VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO i2c_master_top
  CLASS BLOCK ;
  FOREIGN i2c_master_top ;
  ORIGIN 3.500 2.300 ;
  SIZE 559.000 BY 388.600 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.400 380.400 551.600 381.600 ;
        RECT 1.200 377.800 2.000 380.400 ;
        RECT 7.600 375.800 8.400 380.400 ;
        RECT 18.800 377.800 19.600 380.400 ;
        RECT 22.000 377.800 22.800 380.400 ;
        RECT 31.600 375.800 32.400 380.400 ;
        RECT 39.600 375.800 40.400 380.400 ;
        RECT 49.200 377.800 50.000 380.400 ;
        RECT 52.400 377.800 53.200 380.400 ;
        RECT 63.600 375.800 64.400 380.400 ;
        RECT 70.000 377.800 70.800 380.400 ;
        RECT 71.600 377.800 72.400 380.400 ;
        RECT 78.000 375.800 78.800 380.400 ;
        RECT 89.200 377.800 90.000 380.400 ;
        RECT 92.400 377.800 93.200 380.400 ;
        RECT 102.000 375.800 102.800 380.400 ;
        RECT 113.200 377.800 114.000 380.400 ;
        RECT 119.600 375.800 120.400 380.400 ;
        RECT 130.800 377.800 131.600 380.400 ;
        RECT 134.000 377.800 134.800 380.400 ;
        RECT 143.600 375.800 144.400 380.400 ;
        RECT 151.600 375.800 152.400 380.400 ;
        RECT 161.200 377.800 162.000 380.400 ;
        RECT 164.400 377.800 165.200 380.400 ;
        RECT 175.600 375.800 176.400 380.400 ;
        RECT 182.000 377.800 182.800 380.400 ;
        RECT 186.800 375.800 187.600 380.400 ;
        RECT 196.400 377.800 197.200 380.400 ;
        RECT 199.600 377.800 200.400 380.400 ;
        RECT 210.800 375.800 211.600 380.400 ;
        RECT 217.200 377.800 218.000 380.400 ;
        RECT 222.000 375.800 222.800 380.400 ;
        RECT 226.800 376.600 227.600 380.400 ;
        RECT 233.200 376.600 234.000 380.400 ;
        RECT 239.600 375.800 240.400 380.400 ;
        RECT 244.400 376.600 245.200 380.400 ;
        RECT 247.600 375.800 248.400 380.400 ;
        RECT 252.400 377.800 253.200 380.400 ;
        RECT 258.800 375.800 259.600 380.400 ;
        RECT 270.000 377.800 270.800 380.400 ;
        RECT 273.200 377.800 274.000 380.400 ;
        RECT 282.800 375.800 283.600 380.400 ;
        RECT 297.200 376.600 298.000 380.400 ;
        RECT 300.400 375.800 301.200 380.400 ;
        RECT 306.800 375.800 307.600 380.400 ;
        RECT 308.400 373.800 309.200 380.400 ;
        RECT 314.800 377.800 315.600 380.400 ;
        RECT 318.000 377.800 318.800 380.400 ;
        RECT 321.200 376.600 322.000 380.400 ;
        RECT 326.000 373.800 326.800 380.400 ;
        RECT 335.600 375.800 336.400 380.400 ;
        RECT 340.400 375.800 341.200 380.400 ;
        RECT 344.200 376.000 345.000 380.400 ;
        RECT 351.600 375.800 352.400 380.400 ;
        RECT 361.200 377.800 362.000 380.400 ;
        RECT 364.400 377.800 365.200 380.400 ;
        RECT 375.600 375.800 376.400 380.400 ;
        RECT 382.000 377.800 382.800 380.400 ;
        RECT 383.600 377.800 384.400 380.400 ;
        RECT 386.800 377.800 387.600 380.400 ;
        RECT 391.600 376.600 392.400 380.400 ;
        RECT 398.000 375.800 398.800 380.400 ;
        RECT 407.600 377.800 408.400 380.400 ;
        RECT 410.800 377.800 411.600 380.400 ;
        RECT 422.000 375.800 422.800 380.400 ;
        RECT 428.400 377.800 429.200 380.400 ;
        RECT 436.400 377.800 437.200 380.400 ;
        RECT 442.800 375.800 443.600 380.400 ;
        RECT 454.000 377.800 454.800 380.400 ;
        RECT 457.200 377.800 458.000 380.400 ;
        RECT 466.800 375.800 467.600 380.400 ;
        RECT 474.800 375.800 475.600 380.400 ;
        RECT 484.400 377.800 485.200 380.400 ;
        RECT 487.600 377.800 488.400 380.400 ;
        RECT 498.800 375.800 499.600 380.400 ;
        RECT 505.200 377.800 506.000 380.400 ;
        RECT 506.800 375.800 507.600 380.400 ;
        RECT 511.600 377.800 512.400 380.400 ;
        RECT 518.000 375.800 518.800 380.400 ;
        RECT 529.200 377.800 530.000 380.400 ;
        RECT 532.400 377.800 533.200 380.400 ;
        RECT 542.000 375.800 542.800 380.400 ;
        RECT 548.400 377.800 549.200 380.400 ;
        RECT 1.200 341.600 2.000 344.200 ;
        RECT 7.600 341.600 8.400 346.200 ;
        RECT 18.800 341.600 19.600 344.200 ;
        RECT 22.000 341.600 22.800 344.200 ;
        RECT 31.600 341.600 32.400 346.200 ;
        RECT 38.000 341.600 38.800 344.200 ;
        RECT 39.600 341.600 40.400 344.200 ;
        RECT 42.800 341.600 43.600 344.200 ;
        RECT 44.400 341.600 45.200 344.200 ;
        RECT 47.600 341.600 48.400 344.200 ;
        RECT 49.200 341.600 50.000 344.200 ;
        RECT 52.400 341.600 53.200 344.200 ;
        RECT 54.000 341.600 54.800 346.200 ;
        RECT 62.000 341.600 62.800 346.200 ;
        RECT 71.600 341.600 72.400 344.200 ;
        RECT 74.800 341.600 75.600 344.200 ;
        RECT 86.000 341.600 86.800 346.200 ;
        RECT 92.400 341.600 93.200 344.200 ;
        RECT 94.000 341.600 94.800 344.200 ;
        RECT 97.200 341.600 98.000 344.200 ;
        RECT 102.000 341.600 102.800 346.200 ;
        RECT 111.600 341.600 112.400 344.200 ;
        RECT 114.800 341.600 115.600 344.200 ;
        RECT 126.000 341.600 126.800 346.200 ;
        RECT 132.400 341.600 133.200 344.200 ;
        RECT 143.600 341.600 144.400 346.200 ;
        RECT 153.200 341.600 154.000 344.200 ;
        RECT 156.400 341.600 157.200 344.200 ;
        RECT 167.600 341.600 168.400 346.200 ;
        RECT 174.000 341.600 174.800 344.200 ;
        RECT 175.600 341.600 176.400 344.200 ;
        RECT 182.000 341.600 182.800 346.200 ;
        RECT 193.200 341.600 194.000 344.200 ;
        RECT 196.400 341.600 197.200 344.200 ;
        RECT 206.000 341.600 206.800 346.200 ;
        RECT 210.800 341.600 211.600 344.200 ;
        RECT 217.200 341.600 218.000 346.200 ;
        RECT 228.400 341.600 229.200 344.200 ;
        RECT 231.600 341.600 232.400 344.200 ;
        RECT 241.200 341.600 242.000 346.200 ;
        RECT 250.800 341.600 251.600 348.200 ;
        RECT 257.200 341.600 258.000 348.200 ;
        RECT 268.400 341.600 269.200 346.200 ;
        RECT 278.000 341.600 278.800 344.200 ;
        RECT 281.200 341.600 282.000 344.200 ;
        RECT 292.400 341.600 293.200 346.200 ;
        RECT 298.800 341.600 299.600 344.200 ;
        RECT 305.200 341.600 306.000 348.200 ;
        RECT 306.800 341.600 307.600 344.200 ;
        RECT 310.000 341.600 310.800 344.200 ;
        RECT 313.800 341.600 314.600 346.000 ;
        RECT 318.000 341.600 318.800 346.200 ;
        RECT 327.600 341.600 328.400 348.200 ;
        RECT 329.200 341.600 330.000 344.200 ;
        RECT 333.400 341.600 334.200 346.200 ;
        RECT 340.400 341.600 341.200 348.200 ;
        RECT 342.000 341.600 342.800 344.200 ;
        RECT 345.200 341.600 346.000 344.200 ;
        RECT 346.800 341.600 347.600 344.200 ;
        RECT 350.000 341.600 350.800 344.200 ;
        RECT 353.200 341.600 354.000 345.400 ;
        RECT 361.200 341.600 362.000 345.400 ;
        RECT 366.000 341.600 366.800 345.400 ;
        RECT 375.600 341.600 376.400 345.400 ;
        RECT 378.800 341.600 379.600 344.200 ;
        RECT 383.000 341.600 383.800 346.200 ;
        RECT 386.800 341.600 387.600 346.200 ;
        RECT 388.400 341.600 389.200 344.200 ;
        RECT 392.600 341.600 393.400 346.200 ;
        RECT 395.400 341.600 396.200 346.200 ;
        RECT 399.600 341.600 400.400 344.200 ;
        RECT 401.800 341.600 402.600 346.200 ;
        RECT 406.000 341.600 406.800 344.200 ;
        RECT 409.200 341.600 410.000 344.200 ;
        RECT 412.400 341.600 413.200 343.800 ;
        RECT 420.400 341.600 421.200 344.200 ;
        RECT 423.600 341.600 424.400 344.200 ;
        RECT 431.600 341.600 432.400 346.200 ;
        RECT 436.400 341.600 437.200 346.200 ;
        RECT 441.200 341.600 442.000 348.200 ;
        RECT 449.200 341.600 450.000 345.400 ;
        RECT 455.600 341.600 456.400 345.400 ;
        RECT 465.200 341.600 466.000 345.400 ;
        RECT 470.000 341.600 470.800 344.200 ;
        RECT 473.200 341.600 474.000 345.400 ;
        RECT 479.600 341.600 480.400 345.400 ;
        RECT 484.400 341.600 485.200 344.200 ;
        RECT 487.600 341.600 488.400 344.200 ;
        RECT 490.800 341.600 491.600 348.200 ;
        RECT 497.200 341.600 498.000 348.200 ;
        RECT 503.600 341.600 504.400 344.200 ;
        RECT 506.800 341.600 507.600 344.200 ;
        RECT 508.400 341.600 509.200 344.200 ;
        RECT 512.600 341.600 513.400 346.200 ;
        RECT 514.800 341.600 515.600 344.200 ;
        RECT 521.200 341.600 522.000 346.200 ;
        RECT 532.400 341.600 533.200 344.200 ;
        RECT 535.600 341.600 536.400 344.200 ;
        RECT 545.200 341.600 546.000 346.200 ;
        RECT 0.400 340.400 551.600 341.600 ;
        RECT 1.200 337.800 2.000 340.400 ;
        RECT 4.400 337.800 5.200 340.400 ;
        RECT 10.800 335.800 11.600 340.400 ;
        RECT 22.000 337.800 22.800 340.400 ;
        RECT 25.200 337.800 26.000 340.400 ;
        RECT 34.800 335.800 35.600 340.400 ;
        RECT 39.600 335.800 40.400 340.400 ;
        RECT 47.600 336.600 48.400 340.400 ;
        RECT 50.800 333.800 51.600 340.400 ;
        RECT 57.200 333.800 58.000 340.400 ;
        RECT 66.800 336.600 67.600 340.400 ;
        RECT 73.200 335.800 74.000 340.400 ;
        RECT 78.000 335.800 78.800 340.400 ;
        RECT 79.600 337.800 80.400 340.400 ;
        RECT 82.800 337.800 83.600 340.400 ;
        RECT 89.200 333.800 90.000 340.400 ;
        RECT 92.400 337.800 93.200 340.400 ;
        RECT 94.000 337.800 94.800 340.400 ;
        RECT 100.400 335.800 101.200 340.400 ;
        RECT 111.600 337.800 112.400 340.400 ;
        RECT 114.800 337.800 115.600 340.400 ;
        RECT 124.400 335.800 125.200 340.400 ;
        RECT 138.800 335.800 139.600 340.400 ;
        RECT 148.400 337.800 149.200 340.400 ;
        RECT 151.600 337.800 152.400 340.400 ;
        RECT 162.800 335.800 163.600 340.400 ;
        RECT 169.200 337.800 170.000 340.400 ;
        RECT 172.400 335.800 173.200 340.400 ;
        RECT 178.800 336.600 179.600 340.400 ;
        RECT 182.000 337.800 182.800 340.400 ;
        RECT 185.200 333.800 186.000 340.400 ;
        RECT 191.600 337.800 192.400 340.400 ;
        RECT 196.400 336.600 197.200 340.400 ;
        RECT 201.200 335.800 202.000 340.400 ;
        RECT 207.600 335.800 208.400 340.400 ;
        RECT 212.400 337.800 213.200 340.400 ;
        RECT 214.000 337.800 214.800 340.400 ;
        RECT 217.200 337.800 218.000 340.400 ;
        RECT 218.800 337.800 219.600 340.400 ;
        RECT 225.200 335.800 226.000 340.400 ;
        RECT 236.400 337.800 237.200 340.400 ;
        RECT 239.600 337.800 240.400 340.400 ;
        RECT 249.200 335.800 250.000 340.400 ;
        RECT 254.000 335.800 254.800 340.400 ;
        RECT 257.200 335.800 258.000 340.400 ;
        RECT 260.400 335.800 261.200 340.400 ;
        RECT 263.600 335.800 264.400 340.400 ;
        RECT 266.800 335.800 267.600 340.400 ;
        RECT 278.000 335.800 278.800 340.400 ;
        RECT 287.600 337.800 288.400 340.400 ;
        RECT 290.800 337.800 291.600 340.400 ;
        RECT 302.000 335.800 302.800 340.400 ;
        RECT 308.400 337.800 309.200 340.400 ;
        RECT 313.200 335.800 314.000 340.400 ;
        RECT 322.800 337.800 323.600 340.400 ;
        RECT 326.000 337.800 326.800 340.400 ;
        RECT 337.200 335.800 338.000 340.400 ;
        RECT 343.600 337.800 344.400 340.400 ;
        RECT 345.200 335.800 346.000 340.400 ;
        RECT 348.400 335.800 349.200 340.400 ;
        RECT 353.800 335.800 354.600 340.400 ;
        RECT 358.000 337.800 358.800 340.400 ;
        RECT 362.800 336.600 363.600 340.400 ;
        RECT 369.200 336.600 370.000 340.400 ;
        RECT 374.000 337.800 374.800 340.400 ;
        RECT 378.800 335.800 379.600 340.400 ;
        RECT 380.400 335.800 381.200 340.400 ;
        RECT 385.200 335.800 386.000 340.400 ;
        RECT 391.600 336.600 392.400 340.400 ;
        RECT 398.000 335.800 398.800 340.400 ;
        RECT 402.800 335.800 403.600 340.400 ;
        RECT 407.600 336.600 408.400 340.400 ;
        RECT 410.800 337.800 411.600 340.400 ;
        RECT 414.000 337.800 414.800 340.400 ;
        RECT 417.200 337.800 418.000 340.400 ;
        RECT 426.800 337.800 427.600 340.400 ;
        RECT 430.000 338.200 430.800 340.400 ;
        RECT 438.000 333.800 438.800 340.400 ;
        RECT 447.600 336.600 448.400 340.400 ;
        RECT 452.400 335.800 453.200 340.400 ;
        RECT 454.000 337.800 454.800 340.400 ;
        RECT 457.200 337.800 458.000 340.400 ;
        RECT 462.000 335.800 462.800 340.400 ;
        RECT 471.600 337.800 472.400 340.400 ;
        RECT 474.800 337.800 475.600 340.400 ;
        RECT 486.000 335.800 486.800 340.400 ;
        RECT 492.400 337.800 493.200 340.400 ;
        RECT 497.200 335.800 498.000 340.400 ;
        RECT 502.000 336.600 502.800 340.400 ;
        RECT 506.800 337.800 507.600 340.400 ;
        RECT 510.000 336.600 510.800 340.400 ;
        RECT 516.400 336.600 517.200 340.400 ;
        RECT 521.200 337.800 522.000 340.400 ;
        RECT 524.400 337.800 525.200 340.400 ;
        RECT 526.000 337.800 526.800 340.400 ;
        RECT 530.800 336.600 531.600 340.400 ;
        RECT 537.200 336.600 538.000 340.400 ;
        RECT 543.600 337.800 544.400 340.400 ;
        RECT 546.800 335.800 547.600 340.400 ;
        RECT 1.200 301.600 2.000 304.200 ;
        RECT 4.400 301.600 5.200 304.200 ;
        RECT 6.000 301.600 6.800 308.200 ;
        RECT 14.000 301.600 14.800 304.200 ;
        RECT 20.400 301.600 21.200 308.200 ;
        RECT 22.000 301.600 22.800 306.200 ;
        RECT 30.000 301.600 30.800 305.400 ;
        RECT 33.200 301.600 34.000 304.200 ;
        RECT 36.400 301.600 37.200 304.200 ;
        RECT 38.000 301.600 38.800 304.200 ;
        RECT 41.200 301.600 42.000 304.200 ;
        RECT 44.400 301.600 45.200 305.400 ;
        RECT 50.800 301.600 51.600 306.200 ;
        RECT 55.600 301.600 56.400 308.200 ;
        RECT 62.000 301.600 62.800 306.200 ;
        RECT 68.400 301.600 69.200 305.400 ;
        RECT 74.800 301.600 75.600 304.200 ;
        RECT 78.000 301.600 78.800 306.200 ;
        RECT 81.200 301.600 82.000 306.200 ;
        RECT 84.400 301.600 85.200 306.200 ;
        RECT 87.600 301.600 88.400 306.200 ;
        RECT 90.800 301.600 91.600 306.200 ;
        RECT 94.000 301.600 94.800 305.400 ;
        RECT 102.000 301.600 102.800 306.200 ;
        RECT 103.600 301.600 104.400 306.200 ;
        RECT 106.800 301.600 107.600 306.200 ;
        RECT 108.400 301.600 109.200 304.200 ;
        RECT 111.600 301.600 112.400 304.200 ;
        RECT 114.800 301.600 115.600 304.200 ;
        RECT 118.000 301.600 118.800 304.200 ;
        RECT 122.200 301.600 123.000 306.000 ;
        RECT 137.200 301.600 138.000 308.200 ;
        RECT 140.400 301.600 141.200 305.400 ;
        RECT 145.200 301.600 146.000 306.200 ;
        RECT 148.400 301.600 149.200 306.200 ;
        RECT 151.600 301.600 152.400 306.200 ;
        RECT 154.800 301.600 155.600 306.200 ;
        RECT 158.000 301.600 158.800 306.200 ;
        RECT 160.200 301.600 161.000 306.200 ;
        RECT 164.400 301.600 165.200 304.200 ;
        RECT 169.200 301.600 170.000 305.400 ;
        RECT 175.600 301.600 176.400 305.400 ;
        RECT 178.800 301.600 179.600 304.200 ;
        RECT 182.000 301.600 182.800 306.200 ;
        RECT 186.800 301.600 187.600 304.200 ;
        RECT 190.000 301.600 190.800 304.200 ;
        RECT 194.800 301.600 195.600 305.400 ;
        RECT 199.600 301.600 200.400 304.200 ;
        RECT 201.200 301.600 202.000 306.200 ;
        RECT 209.200 301.600 210.000 305.400 ;
        RECT 214.000 301.600 214.800 305.400 ;
        RECT 222.000 301.600 222.800 306.200 ;
        RECT 226.800 301.600 227.600 306.200 ;
        RECT 231.600 301.600 232.400 306.200 ;
        RECT 236.400 301.600 237.200 305.400 ;
        RECT 239.600 301.600 240.400 304.200 ;
        RECT 244.400 301.600 245.200 305.400 ;
        RECT 249.200 301.600 250.000 304.200 ;
        RECT 255.600 301.600 256.400 306.200 ;
        RECT 266.800 301.600 267.600 304.200 ;
        RECT 270.000 301.600 270.800 304.200 ;
        RECT 279.600 301.600 280.400 306.200 ;
        RECT 290.800 301.600 291.600 304.200 ;
        RECT 297.200 301.600 298.000 306.200 ;
        RECT 308.400 301.600 309.200 304.200 ;
        RECT 311.600 301.600 312.400 304.200 ;
        RECT 321.200 301.600 322.000 306.200 ;
        RECT 326.600 301.600 327.400 306.200 ;
        RECT 330.800 301.600 331.600 304.200 ;
        RECT 335.600 301.600 336.400 305.400 ;
        RECT 340.400 301.600 341.200 304.200 ;
        RECT 343.600 301.600 344.400 306.200 ;
        RECT 348.400 301.600 349.200 305.400 ;
        RECT 356.400 301.600 357.200 306.200 ;
        RECT 358.000 301.600 358.800 308.200 ;
        RECT 364.400 301.600 365.200 304.200 ;
        RECT 367.600 301.600 368.400 306.200 ;
        RECT 373.600 301.600 374.400 306.200 ;
        RECT 378.800 301.600 379.600 306.200 ;
        RECT 380.800 301.600 381.600 306.200 ;
        RECT 386.800 301.600 387.600 306.200 ;
        RECT 390.000 301.600 390.800 304.200 ;
        RECT 394.800 301.600 395.600 305.400 ;
        RECT 398.000 301.600 398.800 308.200 ;
        RECT 409.200 301.600 410.000 308.200 ;
        RECT 412.400 301.600 413.200 304.200 ;
        RECT 414.000 301.600 414.800 304.200 ;
        RECT 417.200 301.600 418.000 304.200 ;
        RECT 426.800 301.600 427.600 304.200 ;
        RECT 430.000 301.600 430.800 303.800 ;
        RECT 439.600 301.600 440.400 304.200 ;
        RECT 444.400 301.600 445.200 306.200 ;
        RECT 454.000 301.600 454.800 304.200 ;
        RECT 457.200 301.600 458.000 304.200 ;
        RECT 468.400 301.600 469.200 306.200 ;
        RECT 474.800 301.600 475.600 304.200 ;
        RECT 476.400 301.600 477.200 304.200 ;
        RECT 479.600 301.600 480.400 306.200 ;
        RECT 482.800 301.600 483.600 306.200 ;
        RECT 486.000 301.600 486.800 306.200 ;
        RECT 489.200 301.600 490.000 306.200 ;
        RECT 492.400 301.600 493.200 306.200 ;
        RECT 494.000 301.600 494.800 304.200 ;
        RECT 503.600 301.600 504.400 303.800 ;
        RECT 506.800 301.600 507.600 304.200 ;
        RECT 511.600 301.600 512.400 305.400 ;
        RECT 516.400 301.600 517.200 304.200 ;
        RECT 520.200 301.600 521.000 306.200 ;
        RECT 524.400 301.600 525.200 304.200 ;
        RECT 526.000 301.600 526.800 304.200 ;
        RECT 530.800 301.600 531.600 305.400 ;
        RECT 537.200 301.600 538.000 305.400 ;
        RECT 545.200 301.600 546.000 306.200 ;
        RECT 0.400 300.400 551.600 301.600 ;
        RECT 6.000 293.800 6.800 300.400 ;
        RECT 9.200 297.800 10.000 300.400 ;
        RECT 10.800 297.800 11.600 300.400 ;
        RECT 14.000 297.800 14.800 300.400 ;
        RECT 15.600 297.800 16.400 300.400 ;
        RECT 18.800 297.800 19.600 300.400 ;
        RECT 22.000 293.800 22.800 300.400 ;
        RECT 31.600 295.800 32.400 300.400 ;
        RECT 33.200 297.800 34.000 300.400 ;
        RECT 36.400 297.800 37.200 300.400 ;
        RECT 38.000 297.800 38.800 300.400 ;
        RECT 44.400 295.800 45.200 300.400 ;
        RECT 55.600 297.800 56.400 300.400 ;
        RECT 58.800 297.800 59.600 300.400 ;
        RECT 68.400 295.800 69.200 300.400 ;
        RECT 73.200 297.800 74.000 300.400 ;
        RECT 79.600 295.800 80.400 300.400 ;
        RECT 90.800 297.800 91.600 300.400 ;
        RECT 94.000 297.800 94.800 300.400 ;
        RECT 103.600 295.800 104.400 300.400 ;
        RECT 111.600 295.800 112.400 300.400 ;
        RECT 116.400 296.600 117.200 300.400 ;
        RECT 119.600 297.800 120.400 300.400 ;
        RECT 122.800 297.800 123.600 300.400 ;
        RECT 132.400 296.600 133.200 300.400 ;
        RECT 137.200 297.800 138.000 300.400 ;
        RECT 142.000 296.600 142.800 300.400 ;
        RECT 151.600 293.800 152.400 300.400 ;
        RECT 153.200 297.800 154.000 300.400 ;
        RECT 156.400 297.800 157.200 300.400 ;
        RECT 159.600 296.600 160.400 300.400 ;
        RECT 164.400 295.800 165.200 300.400 ;
        RECT 169.200 297.800 170.000 300.400 ;
        RECT 172.400 297.800 173.200 300.400 ;
        RECT 174.400 295.800 175.200 300.400 ;
        RECT 180.400 295.800 181.200 300.400 ;
        RECT 185.200 295.800 186.000 300.400 ;
        RECT 190.000 296.600 190.800 300.400 ;
        RECT 194.800 296.200 195.600 300.400 ;
        RECT 198.000 297.800 198.800 300.400 ;
        RECT 199.600 295.800 200.400 300.400 ;
        RECT 205.600 295.800 206.400 300.400 ;
        RECT 209.200 296.200 210.000 300.400 ;
        RECT 212.400 297.800 213.200 300.400 ;
        RECT 217.200 295.800 218.000 300.400 ;
        RECT 218.800 295.800 219.600 300.400 ;
        RECT 224.800 295.800 225.600 300.400 ;
        RECT 226.800 295.800 227.600 300.400 ;
        RECT 232.800 295.800 233.600 300.400 ;
        RECT 234.800 295.800 235.600 300.400 ;
        RECT 240.800 295.800 241.600 300.400 ;
        RECT 245.400 296.000 246.200 300.400 ;
        RECT 249.200 297.800 250.000 300.400 ;
        RECT 253.000 295.800 253.800 300.400 ;
        RECT 257.200 297.800 258.000 300.400 ;
        RECT 258.800 297.800 259.600 300.400 ;
        RECT 263.600 296.600 264.400 300.400 ;
        RECT 274.800 297.800 275.600 300.400 ;
        RECT 281.200 295.800 282.000 300.400 ;
        RECT 292.400 297.800 293.200 300.400 ;
        RECT 295.600 297.800 296.400 300.400 ;
        RECT 305.200 295.800 306.000 300.400 ;
        RECT 310.000 295.800 310.800 300.400 ;
        RECT 313.200 295.800 314.000 300.400 ;
        RECT 316.400 295.800 317.200 300.400 ;
        RECT 319.600 295.800 320.400 300.400 ;
        RECT 322.800 295.800 323.600 300.400 ;
        RECT 329.200 293.800 330.000 300.400 ;
        RECT 330.800 297.800 331.600 300.400 ;
        RECT 335.600 296.600 336.400 300.400 ;
        RECT 343.600 296.600 344.400 300.400 ;
        RECT 346.800 297.800 347.600 300.400 ;
        RECT 350.000 297.800 350.800 300.400 ;
        RECT 353.200 297.800 354.000 300.400 ;
        RECT 356.400 298.200 357.200 300.400 ;
        RECT 364.400 297.800 365.200 300.400 ;
        RECT 368.600 295.800 369.400 300.400 ;
        RECT 372.400 295.800 373.200 300.400 ;
        RECT 375.600 297.800 376.400 300.400 ;
        RECT 380.400 296.600 381.200 300.400 ;
        RECT 383.600 297.800 384.400 300.400 ;
        RECT 386.800 297.800 387.600 300.400 ;
        RECT 391.600 295.800 392.400 300.400 ;
        RECT 394.800 296.600 395.600 300.400 ;
        RECT 402.800 295.800 403.600 300.400 ;
        RECT 404.400 295.800 405.200 300.400 ;
        RECT 409.200 297.800 410.000 300.400 ;
        RECT 413.400 295.800 414.200 300.400 ;
        RECT 415.600 297.800 416.400 300.400 ;
        RECT 418.800 297.800 419.600 300.400 ;
        RECT 422.000 297.800 422.800 300.400 ;
        RECT 431.600 295.800 432.400 300.400 ;
        RECT 435.200 295.800 436.000 300.400 ;
        RECT 441.200 295.800 442.000 300.400 ;
        RECT 446.000 295.800 446.800 300.400 ;
        RECT 447.600 297.800 448.400 300.400 ;
        RECT 450.800 297.800 451.600 300.400 ;
        RECT 457.200 295.800 458.000 300.400 ;
        RECT 468.400 297.800 469.200 300.400 ;
        RECT 471.600 297.800 472.400 300.400 ;
        RECT 481.200 295.800 482.000 300.400 ;
        RECT 486.000 297.800 486.800 300.400 ;
        RECT 490.200 295.800 491.000 300.400 ;
        RECT 497.200 296.600 498.000 300.400 ;
        RECT 502.000 295.800 502.800 300.400 ;
        RECT 503.600 297.800 504.400 300.400 ;
        RECT 506.800 297.800 507.600 300.400 ;
        RECT 511.600 295.800 512.400 300.400 ;
        RECT 513.200 297.800 514.000 300.400 ;
        RECT 519.600 295.800 520.400 300.400 ;
        RECT 530.800 297.800 531.600 300.400 ;
        RECT 534.000 297.800 534.800 300.400 ;
        RECT 543.600 295.800 544.400 300.400 ;
        RECT 1.200 261.600 2.000 264.200 ;
        RECT 7.600 261.600 8.400 266.200 ;
        RECT 18.800 261.600 19.600 264.200 ;
        RECT 22.000 261.600 22.800 264.200 ;
        RECT 31.600 261.600 32.400 266.200 ;
        RECT 38.000 261.600 38.800 265.400 ;
        RECT 47.600 261.600 48.400 266.200 ;
        RECT 49.200 261.600 50.000 264.200 ;
        RECT 52.400 261.600 53.200 264.200 ;
        RECT 56.600 261.600 57.400 266.000 ;
        RECT 63.600 261.600 64.400 266.200 ;
        RECT 68.400 261.600 69.200 266.200 ;
        RECT 73.200 261.600 74.000 265.400 ;
        RECT 76.400 261.600 77.200 264.200 ;
        RECT 79.600 261.600 80.400 264.200 ;
        RECT 83.800 261.600 84.600 266.000 ;
        RECT 87.600 261.600 88.400 264.200 ;
        RECT 94.000 261.600 94.800 266.200 ;
        RECT 103.600 261.600 104.400 264.200 ;
        RECT 106.800 261.600 107.600 264.200 ;
        RECT 118.000 261.600 118.800 266.200 ;
        RECT 124.400 261.600 125.200 264.200 ;
        RECT 132.400 261.600 133.200 266.200 ;
        RECT 138.400 261.600 139.200 266.200 ;
        RECT 143.600 261.600 144.400 266.200 ;
        RECT 148.400 261.600 149.200 265.400 ;
        RECT 151.600 261.600 152.400 264.200 ;
        RECT 155.800 261.600 156.600 266.200 ;
        RECT 158.000 261.600 158.800 264.200 ;
        RECT 161.200 261.600 162.000 264.200 ;
        RECT 162.800 261.600 163.600 266.200 ;
        RECT 167.600 261.600 168.400 266.200 ;
        RECT 172.400 261.600 173.200 268.200 ;
        RECT 182.000 261.600 182.800 266.200 ;
        RECT 186.800 261.600 187.600 265.400 ;
        RECT 193.200 261.600 194.000 265.400 ;
        RECT 196.400 261.600 197.200 268.200 ;
        RECT 204.400 261.600 205.200 264.200 ;
        RECT 206.000 261.600 206.800 264.200 ;
        RECT 209.200 261.600 210.000 264.200 ;
        RECT 210.800 261.600 211.600 264.200 ;
        RECT 214.000 261.600 214.800 264.200 ;
        RECT 217.200 261.600 218.000 265.400 ;
        RECT 222.000 261.600 222.800 266.200 ;
        RECT 226.800 261.600 227.600 264.200 ;
        RECT 231.600 261.600 232.400 265.400 ;
        RECT 236.400 261.600 237.200 266.200 ;
        RECT 242.400 261.600 243.200 266.200 ;
        RECT 244.400 261.600 245.200 264.200 ;
        RECT 249.200 261.600 250.000 265.400 ;
        RECT 258.800 261.600 259.600 265.400 ;
        RECT 268.400 261.600 269.200 264.200 ;
        RECT 274.800 261.600 275.600 266.200 ;
        RECT 286.000 261.600 286.800 264.200 ;
        RECT 289.200 261.600 290.000 264.200 ;
        RECT 298.800 261.600 299.600 266.200 ;
        RECT 306.800 261.600 307.600 266.200 ;
        RECT 316.400 261.600 317.200 264.200 ;
        RECT 319.600 261.600 320.400 264.200 ;
        RECT 330.800 261.600 331.600 266.200 ;
        RECT 337.200 261.600 338.000 264.200 ;
        RECT 338.800 261.600 339.600 264.200 ;
        RECT 344.600 261.600 345.400 266.000 ;
        RECT 351.600 261.600 352.400 266.200 ;
        RECT 361.200 261.600 362.000 264.200 ;
        RECT 364.400 261.600 365.200 264.200 ;
        RECT 375.600 261.600 376.400 266.200 ;
        RECT 382.000 261.600 382.800 264.200 ;
        RECT 386.800 261.600 387.600 266.200 ;
        RECT 396.400 261.600 397.200 264.200 ;
        RECT 399.600 261.600 400.400 264.200 ;
        RECT 410.800 261.600 411.600 266.200 ;
        RECT 417.200 261.600 418.000 264.200 ;
        RECT 418.800 261.600 419.600 264.200 ;
        RECT 422.000 261.600 422.800 264.200 ;
        RECT 430.000 261.600 430.800 264.200 ;
        RECT 434.800 261.600 435.600 265.400 ;
        RECT 441.200 261.600 442.000 265.400 ;
        RECT 446.000 261.600 446.800 264.200 ;
        RECT 450.800 261.600 451.600 264.200 ;
        RECT 452.400 261.600 453.200 264.200 ;
        RECT 458.800 261.600 459.600 266.200 ;
        RECT 470.000 261.600 470.800 264.200 ;
        RECT 473.200 261.600 474.000 264.200 ;
        RECT 482.800 261.600 483.600 266.200 ;
        RECT 487.600 261.600 488.400 264.200 ;
        RECT 494.000 261.600 494.800 266.200 ;
        RECT 505.200 261.600 506.000 264.200 ;
        RECT 508.400 261.600 509.200 264.200 ;
        RECT 518.000 261.600 518.800 266.200 ;
        RECT 524.400 261.600 525.200 264.200 ;
        RECT 527.600 261.600 528.400 266.200 ;
        RECT 533.000 261.600 534.000 264.200 ;
        RECT 536.400 261.600 537.200 264.200 ;
        RECT 542.000 261.600 542.800 266.000 ;
        RECT 546.800 261.600 547.600 266.200 ;
        RECT 0.400 260.400 551.600 261.600 ;
        RECT 1.200 257.800 2.000 260.400 ;
        RECT 4.400 257.800 5.200 260.400 ;
        RECT 7.600 257.800 8.400 260.400 ;
        RECT 9.200 255.800 10.000 260.400 ;
        RECT 16.600 256.000 17.400 260.400 ;
        RECT 20.400 257.800 21.200 260.400 ;
        RECT 23.600 257.800 24.400 260.400 ;
        RECT 27.800 256.000 28.600 260.400 ;
        RECT 33.200 256.600 34.000 260.400 ;
        RECT 38.000 257.800 38.800 260.400 ;
        RECT 41.200 257.800 42.000 260.400 ;
        RECT 42.800 255.800 43.600 260.400 ;
        RECT 47.600 253.800 48.400 260.400 ;
        RECT 54.000 255.800 54.800 260.400 ;
        RECT 62.000 255.800 62.800 260.400 ;
        RECT 63.600 257.800 64.400 260.400 ;
        RECT 66.800 257.800 67.600 260.400 ;
        RECT 71.600 256.600 72.400 260.400 ;
        RECT 74.800 257.800 75.600 260.400 ;
        RECT 78.000 257.800 78.800 260.400 ;
        RECT 79.600 257.800 80.400 260.400 ;
        RECT 86.000 255.800 86.800 260.400 ;
        RECT 97.200 257.800 98.000 260.400 ;
        RECT 100.400 257.800 101.200 260.400 ;
        RECT 110.000 255.800 110.800 260.400 ;
        RECT 121.200 258.200 122.000 260.400 ;
        RECT 124.400 257.800 125.200 260.400 ;
        RECT 134.000 255.800 134.800 260.400 ;
        RECT 140.000 255.800 140.800 260.400 ;
        RECT 143.600 257.800 144.400 260.400 ;
        RECT 148.400 255.800 149.200 260.400 ;
        RECT 158.000 257.800 158.800 260.400 ;
        RECT 161.200 257.800 162.000 260.400 ;
        RECT 172.400 255.800 173.200 260.400 ;
        RECT 178.800 257.800 179.600 260.400 ;
        RECT 180.400 255.800 181.200 260.400 ;
        RECT 183.600 255.800 184.400 260.400 ;
        RECT 185.200 255.800 186.000 260.400 ;
        RECT 191.600 257.800 192.400 260.400 ;
        RECT 196.400 256.600 197.200 260.400 ;
        RECT 199.600 257.800 200.400 260.400 ;
        RECT 202.800 256.200 203.600 260.400 ;
        RECT 206.000 257.800 206.800 260.400 ;
        RECT 212.400 255.800 213.200 260.400 ;
        RECT 223.600 257.800 224.400 260.400 ;
        RECT 226.800 257.800 227.600 260.400 ;
        RECT 236.400 255.800 237.200 260.400 ;
        RECT 244.400 255.800 245.200 260.400 ;
        RECT 246.000 257.800 246.800 260.400 ;
        RECT 252.400 255.800 253.200 260.400 ;
        RECT 263.600 257.800 264.400 260.400 ;
        RECT 266.800 257.800 267.600 260.400 ;
        RECT 276.400 255.800 277.200 260.400 ;
        RECT 287.600 257.800 288.400 260.400 ;
        RECT 294.000 255.800 294.800 260.400 ;
        RECT 305.200 257.800 306.000 260.400 ;
        RECT 308.400 257.800 309.200 260.400 ;
        RECT 318.000 255.800 318.800 260.400 ;
        RECT 326.000 256.600 326.800 260.400 ;
        RECT 332.400 256.600 333.200 260.400 ;
        RECT 335.600 255.800 336.400 260.400 ;
        RECT 338.800 255.800 339.600 260.400 ;
        RECT 340.400 257.800 341.200 260.400 ;
        RECT 345.200 256.600 346.000 260.400 ;
        RECT 353.200 255.800 354.000 260.400 ;
        RECT 362.800 257.800 363.600 260.400 ;
        RECT 366.000 257.800 366.800 260.400 ;
        RECT 377.200 255.800 378.000 260.400 ;
        RECT 383.600 257.800 384.400 260.400 ;
        RECT 386.800 257.800 387.600 260.400 ;
        RECT 388.400 257.800 389.200 260.400 ;
        RECT 394.800 255.800 395.600 260.400 ;
        RECT 406.000 257.800 406.800 260.400 ;
        RECT 409.200 257.800 410.000 260.400 ;
        RECT 418.800 255.800 419.600 260.400 ;
        RECT 430.000 257.800 430.800 260.400 ;
        RECT 433.200 257.800 434.000 260.400 ;
        RECT 439.600 255.800 440.400 260.400 ;
        RECT 450.800 257.800 451.600 260.400 ;
        RECT 454.000 257.800 454.800 260.400 ;
        RECT 463.600 255.800 464.400 260.400 ;
        RECT 468.400 257.800 469.200 260.400 ;
        RECT 472.600 255.800 473.400 260.400 ;
        RECT 474.800 257.800 475.600 260.400 ;
        RECT 478.000 257.800 478.800 260.400 ;
        RECT 482.800 255.800 483.600 260.400 ;
        RECT 492.400 257.800 493.200 260.400 ;
        RECT 495.600 257.800 496.400 260.400 ;
        RECT 506.800 255.800 507.600 260.400 ;
        RECT 513.200 257.800 514.000 260.400 ;
        RECT 514.800 255.800 515.600 260.400 ;
        RECT 518.000 255.800 518.800 260.400 ;
        RECT 521.200 255.800 522.000 260.400 ;
        RECT 524.400 255.800 525.200 260.400 ;
        RECT 527.600 255.800 528.400 260.400 ;
        RECT 530.800 256.000 531.600 260.400 ;
        RECT 536.400 257.800 537.200 260.400 ;
        RECT 539.600 257.800 540.600 260.400 ;
        RECT 545.200 255.800 546.000 260.400 ;
        RECT 1.200 221.600 2.000 224.200 ;
        RECT 7.600 221.600 8.400 226.200 ;
        RECT 18.800 221.600 19.600 224.200 ;
        RECT 22.000 221.600 22.800 224.200 ;
        RECT 31.600 221.600 32.400 226.200 ;
        RECT 36.400 221.600 37.200 228.200 ;
        RECT 44.400 221.600 45.200 225.400 ;
        RECT 50.800 221.600 51.600 224.200 ;
        RECT 54.000 221.600 54.800 224.200 ;
        RECT 57.800 221.600 58.600 226.000 ;
        RECT 65.200 221.600 66.000 226.200 ;
        RECT 71.600 221.600 72.400 228.200 ;
        RECT 75.800 221.600 76.600 226.000 ;
        RECT 79.600 221.600 80.400 224.200 ;
        RECT 83.800 221.600 84.600 226.200 ;
        RECT 86.000 221.600 86.800 224.200 ;
        RECT 89.200 221.600 90.000 224.200 ;
        RECT 93.400 221.600 94.200 226.000 ;
        RECT 97.200 221.600 98.000 224.200 ;
        RECT 101.400 221.600 102.200 226.200 ;
        RECT 103.600 221.600 104.400 224.200 ;
        RECT 110.000 221.600 110.800 226.200 ;
        RECT 121.200 221.600 122.000 224.200 ;
        RECT 124.400 221.600 125.200 224.200 ;
        RECT 134.000 221.600 134.800 226.200 ;
        RECT 145.200 221.600 146.000 226.200 ;
        RECT 148.400 221.600 149.200 226.200 ;
        RECT 151.600 221.600 152.400 224.200 ;
        RECT 156.400 221.600 157.200 225.400 ;
        RECT 161.200 221.600 162.000 225.400 ;
        RECT 169.200 221.600 170.000 226.200 ;
        RECT 173.400 221.600 174.200 226.000 ;
        RECT 177.200 221.600 178.000 226.200 ;
        RECT 183.600 221.600 184.400 226.200 ;
        RECT 186.800 221.600 187.600 226.200 ;
        RECT 194.800 221.600 195.600 225.400 ;
        RECT 199.600 221.600 200.400 225.400 ;
        RECT 204.400 221.600 205.200 224.200 ;
        RECT 210.800 221.600 211.600 226.200 ;
        RECT 222.000 221.600 222.800 224.200 ;
        RECT 225.200 221.600 226.000 224.200 ;
        RECT 234.800 221.600 235.600 226.200 ;
        RECT 239.600 221.600 240.400 224.200 ;
        RECT 246.000 221.600 246.800 226.200 ;
        RECT 257.200 221.600 258.000 224.200 ;
        RECT 260.400 221.600 261.200 224.200 ;
        RECT 270.000 221.600 270.800 226.200 ;
        RECT 281.200 221.600 282.000 224.200 ;
        RECT 284.400 221.600 285.200 224.200 ;
        RECT 290.800 221.600 291.600 226.200 ;
        RECT 302.000 221.600 302.800 224.200 ;
        RECT 305.200 221.600 306.000 224.200 ;
        RECT 314.800 221.600 315.600 226.200 ;
        RECT 321.200 221.600 322.000 225.400 ;
        RECT 327.600 221.600 328.400 225.400 ;
        RECT 335.600 221.600 336.400 225.400 ;
        RECT 342.000 221.600 342.800 225.400 ;
        RECT 346.800 221.600 347.600 226.200 ;
        RECT 351.600 221.600 352.400 226.200 ;
        RECT 356.400 221.600 357.200 225.400 ;
        RECT 362.800 221.600 363.600 226.200 ;
        RECT 369.200 221.600 370.000 225.400 ;
        RECT 372.400 221.600 373.200 226.200 ;
        RECT 377.200 221.600 378.000 224.200 ;
        RECT 383.600 221.600 384.400 226.200 ;
        RECT 394.800 221.600 395.600 224.200 ;
        RECT 398.000 221.600 398.800 224.200 ;
        RECT 407.600 221.600 408.400 226.200 ;
        RECT 412.400 221.600 413.200 224.200 ;
        RECT 417.200 221.600 418.000 225.400 ;
        RECT 428.400 221.600 429.200 228.200 ;
        RECT 434.800 221.600 435.600 224.200 ;
        RECT 438.000 221.600 438.800 224.200 ;
        RECT 439.600 221.600 440.400 228.200 ;
        RECT 446.000 221.600 446.800 226.200 ;
        RECT 452.400 221.600 453.200 225.400 ;
        RECT 457.200 221.600 458.000 228.200 ;
        RECT 463.600 221.600 464.400 228.200 ;
        RECT 470.000 221.600 470.800 224.200 ;
        RECT 473.200 221.600 474.000 224.200 ;
        RECT 474.800 221.600 475.600 224.200 ;
        RECT 478.000 221.600 478.800 224.200 ;
        RECT 480.200 221.600 481.000 226.200 ;
        RECT 484.400 221.600 485.200 224.200 ;
        RECT 486.000 221.600 486.800 226.200 ;
        RECT 494.000 221.600 494.800 226.200 ;
        RECT 495.600 221.600 496.400 224.200 ;
        RECT 502.000 221.600 502.800 226.200 ;
        RECT 513.200 221.600 514.000 224.200 ;
        RECT 516.400 221.600 517.200 224.200 ;
        RECT 526.000 221.600 526.800 226.200 ;
        RECT 530.800 221.600 531.600 224.200 ;
        RECT 535.000 221.600 535.800 226.200 ;
        RECT 540.400 221.600 541.200 226.200 ;
        RECT 542.000 221.600 542.800 224.200 ;
        RECT 545.200 221.600 546.000 224.200 ;
        RECT 548.400 221.600 549.200 226.200 ;
        RECT 0.400 220.400 551.600 221.600 ;
        RECT 1.200 215.800 2.000 220.400 ;
        RECT 4.400 215.800 5.200 220.400 ;
        RECT 6.000 217.800 6.800 220.400 ;
        RECT 9.200 217.800 10.000 220.400 ;
        RECT 11.200 215.800 12.000 220.400 ;
        RECT 17.200 215.800 18.000 220.400 ;
        RECT 22.000 215.800 22.800 220.400 ;
        RECT 28.400 213.800 29.200 220.400 ;
        RECT 32.600 216.000 33.400 220.400 ;
        RECT 39.000 216.000 39.800 220.400 ;
        RECT 47.600 213.800 48.400 220.400 ;
        RECT 50.800 217.800 51.600 220.400 ;
        RECT 54.000 218.200 54.800 220.400 ;
        RECT 62.000 213.800 62.800 220.400 ;
        RECT 68.400 213.800 69.200 220.400 ;
        RECT 74.800 213.800 75.600 220.400 ;
        RECT 81.200 217.800 82.000 220.400 ;
        RECT 84.400 216.200 85.200 220.400 ;
        RECT 90.800 215.800 91.600 220.400 ;
        RECT 93.000 215.800 93.800 220.400 ;
        RECT 97.200 217.800 98.000 220.400 ;
        RECT 98.800 215.800 99.600 220.400 ;
        RECT 105.200 216.600 106.000 220.400 ;
        RECT 119.600 215.800 120.400 220.400 ;
        RECT 129.200 217.800 130.000 220.400 ;
        RECT 132.400 217.800 133.200 220.400 ;
        RECT 143.600 215.800 144.400 220.400 ;
        RECT 150.000 217.800 150.800 220.400 ;
        RECT 151.600 217.800 152.400 220.400 ;
        RECT 154.800 217.800 155.600 220.400 ;
        RECT 156.400 215.800 157.200 220.400 ;
        RECT 162.800 216.600 163.600 220.400 ;
        RECT 167.600 215.800 168.400 220.400 ;
        RECT 173.600 215.800 174.400 220.400 ;
        RECT 177.200 217.800 178.000 220.400 ;
        RECT 181.400 216.000 182.200 220.400 ;
        RECT 185.200 217.800 186.000 220.400 ;
        RECT 188.400 217.800 189.200 220.400 ;
        RECT 191.600 216.600 192.400 220.400 ;
        RECT 196.400 215.800 197.200 220.400 ;
        RECT 206.000 213.800 206.800 220.400 ;
        RECT 207.600 215.800 208.400 220.400 ;
        RECT 213.600 215.800 214.400 220.400 ;
        RECT 218.800 215.800 219.600 220.400 ;
        RECT 222.000 216.600 222.800 220.400 ;
        RECT 228.400 216.600 229.200 220.400 ;
        RECT 233.800 215.800 234.600 220.400 ;
        RECT 238.000 217.800 238.800 220.400 ;
        RECT 242.800 216.600 243.600 220.400 ;
        RECT 246.000 217.800 246.800 220.400 ;
        RECT 252.400 215.800 253.200 220.400 ;
        RECT 263.600 217.800 264.400 220.400 ;
        RECT 266.800 217.800 267.600 220.400 ;
        RECT 276.400 215.800 277.200 220.400 ;
        RECT 287.600 217.800 288.400 220.400 ;
        RECT 290.800 217.800 291.600 220.400 ;
        RECT 297.200 215.800 298.000 220.400 ;
        RECT 308.400 217.800 309.200 220.400 ;
        RECT 311.600 217.800 312.400 220.400 ;
        RECT 321.200 215.800 322.000 220.400 ;
        RECT 326.000 217.800 326.800 220.400 ;
        RECT 330.800 216.600 331.600 220.400 ;
        RECT 338.800 216.600 339.600 220.400 ;
        RECT 342.000 217.800 342.800 220.400 ;
        RECT 346.800 216.000 347.600 220.400 ;
        RECT 352.400 217.800 353.200 220.400 ;
        RECT 355.600 217.800 356.600 220.400 ;
        RECT 361.200 215.800 362.000 220.400 ;
        RECT 367.600 216.600 368.400 220.400 ;
        RECT 375.600 216.600 376.400 220.400 ;
        RECT 378.800 217.800 379.600 220.400 ;
        RECT 383.000 215.800 383.800 220.400 ;
        RECT 385.200 215.800 386.000 220.400 ;
        RECT 391.600 216.600 392.400 220.400 ;
        RECT 401.200 216.600 402.000 220.400 ;
        RECT 409.200 216.600 410.000 220.400 ;
        RECT 412.400 217.800 413.200 220.400 ;
        RECT 415.600 217.800 416.400 220.400 ;
        RECT 420.400 216.600 421.200 220.400 ;
        RECT 430.000 215.800 430.800 220.400 ;
        RECT 436.000 215.800 436.800 220.400 ;
        RECT 438.000 217.800 438.800 220.400 ;
        RECT 441.200 217.800 442.000 220.400 ;
        RECT 442.800 217.800 443.600 220.400 ;
        RECT 446.000 217.800 446.800 220.400 ;
        RECT 452.400 216.600 453.200 220.400 ;
        RECT 457.200 216.600 458.000 220.400 ;
        RECT 465.200 215.400 466.000 220.400 ;
        RECT 470.400 215.000 471.200 220.400 ;
        RECT 474.800 216.600 475.600 220.400 ;
        RECT 479.600 217.800 480.400 220.400 ;
        RECT 486.000 215.800 486.800 220.400 ;
        RECT 497.200 217.800 498.000 220.400 ;
        RECT 500.400 217.800 501.200 220.400 ;
        RECT 510.000 215.800 510.800 220.400 ;
        RECT 518.000 215.800 518.800 220.400 ;
        RECT 527.600 217.800 528.400 220.400 ;
        RECT 530.800 217.800 531.600 220.400 ;
        RECT 542.000 215.800 542.800 220.400 ;
        RECT 548.400 217.800 549.200 220.400 ;
        RECT 1.200 181.600 2.000 186.200 ;
        RECT 9.200 181.600 10.000 186.200 ;
        RECT 10.800 181.600 11.600 184.200 ;
        RECT 14.000 181.600 14.800 184.200 ;
        RECT 18.200 181.600 19.000 186.000 ;
        RECT 22.000 181.600 22.800 184.200 ;
        RECT 25.200 181.600 26.000 184.200 ;
        RECT 26.800 181.600 27.600 184.200 ;
        RECT 30.000 181.600 30.800 185.800 ;
        RECT 33.200 181.600 34.000 188.200 ;
        RECT 44.400 181.600 45.200 188.200 ;
        RECT 46.000 181.600 46.800 184.200 ;
        RECT 49.200 181.600 50.000 186.200 ;
        RECT 58.800 181.600 59.600 188.200 ;
        RECT 63.000 181.600 63.800 186.000 ;
        RECT 70.000 181.600 70.800 186.200 ;
        RECT 79.600 181.600 80.400 184.200 ;
        RECT 82.800 181.600 83.600 184.200 ;
        RECT 94.000 181.600 94.800 186.200 ;
        RECT 100.400 181.600 101.200 184.200 ;
        RECT 102.000 181.600 102.800 184.200 ;
        RECT 108.400 181.600 109.200 186.200 ;
        RECT 119.600 181.600 120.400 184.200 ;
        RECT 122.800 181.600 123.600 184.200 ;
        RECT 132.400 181.600 133.200 186.200 ;
        RECT 146.800 181.600 147.600 186.200 ;
        RECT 156.400 181.600 157.200 184.200 ;
        RECT 159.600 181.600 160.400 184.200 ;
        RECT 170.800 181.600 171.600 186.200 ;
        RECT 177.200 181.600 178.000 184.200 ;
        RECT 180.400 181.600 181.200 186.200 ;
        RECT 182.000 181.600 182.800 184.200 ;
        RECT 188.400 181.600 189.200 186.200 ;
        RECT 199.600 181.600 200.400 184.200 ;
        RECT 202.800 181.600 203.600 184.200 ;
        RECT 212.400 181.600 213.200 186.200 ;
        RECT 218.800 181.600 219.600 184.200 ;
        RECT 225.200 181.600 226.000 188.200 ;
        RECT 228.400 181.600 229.200 184.200 ;
        RECT 230.000 181.600 230.800 186.200 ;
        RECT 234.800 181.600 235.600 184.200 ;
        RECT 238.000 181.600 238.800 184.200 ;
        RECT 242.800 181.600 243.600 186.200 ;
        RECT 244.400 181.600 245.200 184.200 ;
        RECT 249.200 181.600 250.000 185.400 ;
        RECT 254.600 181.600 255.400 186.200 ;
        RECT 258.800 181.600 259.600 184.200 ;
        RECT 266.800 181.600 267.600 184.200 ;
        RECT 273.200 181.600 274.000 186.200 ;
        RECT 284.400 181.600 285.200 184.200 ;
        RECT 287.600 181.600 288.400 184.200 ;
        RECT 297.200 181.600 298.000 186.200 ;
        RECT 302.000 181.600 302.800 184.200 ;
        RECT 308.400 181.600 309.200 186.200 ;
        RECT 319.600 181.600 320.400 184.200 ;
        RECT 322.800 181.600 323.600 184.200 ;
        RECT 332.400 181.600 333.200 186.200 ;
        RECT 337.200 181.600 338.000 184.200 ;
        RECT 342.000 181.600 342.800 185.400 ;
        RECT 350.000 181.600 350.800 186.200 ;
        RECT 359.600 181.600 360.400 184.200 ;
        RECT 362.800 181.600 363.600 184.200 ;
        RECT 374.000 181.600 374.800 186.200 ;
        RECT 380.400 181.600 381.200 184.200 ;
        RECT 385.200 181.600 386.000 185.400 ;
        RECT 388.400 181.600 389.200 188.200 ;
        RECT 398.000 181.600 398.800 186.200 ;
        RECT 401.200 181.600 402.000 185.400 ;
        RECT 406.000 181.600 406.800 184.200 ;
        RECT 409.200 181.600 410.000 188.200 ;
        RECT 417.200 181.600 418.000 184.200 ;
        RECT 420.400 181.600 421.200 185.400 ;
        RECT 433.200 181.600 434.000 184.200 ;
        RECT 436.400 181.600 437.200 186.600 ;
        RECT 441.600 181.600 442.400 187.000 ;
        RECT 449.200 181.600 450.000 188.200 ;
        RECT 452.400 181.600 453.200 186.200 ;
        RECT 460.400 181.600 461.200 188.200 ;
        RECT 465.200 181.600 466.000 185.400 ;
        RECT 468.400 181.600 469.200 184.200 ;
        RECT 474.800 181.600 475.600 186.200 ;
        RECT 486.000 181.600 486.800 184.200 ;
        RECT 489.200 181.600 490.000 184.200 ;
        RECT 498.800 181.600 499.600 186.200 ;
        RECT 505.200 181.600 506.000 185.400 ;
        RECT 513.200 181.600 514.000 186.600 ;
        RECT 518.400 181.600 519.200 187.000 ;
        RECT 522.800 181.600 523.600 186.200 ;
        RECT 528.200 181.600 529.200 184.200 ;
        RECT 531.600 181.600 532.400 184.200 ;
        RECT 537.200 181.600 538.000 186.000 ;
        RECT 542.000 181.600 542.800 185.400 ;
        RECT 550.000 181.600 550.800 186.200 ;
        RECT 0.400 180.400 551.600 181.600 ;
        RECT 1.200 177.800 2.000 180.400 ;
        RECT 4.400 177.800 5.200 180.400 ;
        RECT 7.600 177.800 8.400 180.400 ;
        RECT 9.200 177.800 10.000 180.400 ;
        RECT 12.400 177.800 13.200 180.400 ;
        RECT 14.000 177.800 14.800 180.400 ;
        RECT 17.200 177.800 18.000 180.400 ;
        RECT 18.800 177.800 19.600 180.400 ;
        RECT 23.600 177.800 24.400 180.400 ;
        RECT 30.000 173.800 30.800 180.400 ;
        RECT 31.600 173.800 32.400 180.400 ;
        RECT 39.600 176.600 40.400 180.400 ;
        RECT 46.000 175.800 46.800 180.400 ;
        RECT 54.000 175.800 54.800 180.400 ;
        RECT 55.600 177.800 56.400 180.400 ;
        RECT 62.000 175.800 62.800 180.400 ;
        RECT 73.200 177.800 74.000 180.400 ;
        RECT 76.400 177.800 77.200 180.400 ;
        RECT 86.000 175.800 86.800 180.400 ;
        RECT 92.400 176.600 93.200 180.400 ;
        RECT 97.200 177.800 98.000 180.400 ;
        RECT 100.400 177.800 101.200 180.400 ;
        RECT 102.000 175.800 102.800 180.400 ;
        RECT 108.000 175.800 108.800 180.400 ;
        RECT 116.400 177.800 117.200 180.400 ;
        RECT 122.800 175.800 123.600 180.400 ;
        RECT 134.000 177.800 134.800 180.400 ;
        RECT 137.200 177.800 138.000 180.400 ;
        RECT 146.800 175.800 147.600 180.400 ;
        RECT 154.800 175.800 155.600 180.400 ;
        RECT 164.400 177.800 165.200 180.400 ;
        RECT 167.600 177.800 168.400 180.400 ;
        RECT 178.800 175.800 179.600 180.400 ;
        RECT 185.200 177.800 186.000 180.400 ;
        RECT 186.800 175.800 187.600 180.400 ;
        RECT 191.600 177.800 192.400 180.400 ;
        RECT 195.800 175.800 196.600 180.400 ;
        RECT 199.600 177.800 200.400 180.400 ;
        RECT 201.200 177.800 202.000 180.400 ;
        RECT 207.600 175.800 208.400 180.400 ;
        RECT 218.800 177.800 219.600 180.400 ;
        RECT 222.000 177.800 222.800 180.400 ;
        RECT 231.600 175.800 232.400 180.400 ;
        RECT 236.400 177.800 237.200 180.400 ;
        RECT 240.600 175.800 241.400 180.400 ;
        RECT 244.400 177.800 245.200 180.400 ;
        RECT 249.200 176.600 250.000 180.400 ;
        RECT 255.600 175.800 256.400 180.400 ;
        RECT 257.200 177.800 258.000 180.400 ;
        RECT 261.400 175.800 262.200 180.400 ;
        RECT 268.400 173.800 269.200 180.400 ;
        RECT 270.000 177.800 270.800 180.400 ;
        RECT 274.200 175.800 275.000 180.400 ;
        RECT 284.400 176.600 285.200 180.400 ;
        RECT 289.200 177.800 290.000 180.400 ;
        RECT 292.400 177.800 293.200 180.400 ;
        RECT 294.000 177.800 294.800 180.400 ;
        RECT 300.400 175.800 301.200 180.400 ;
        RECT 311.600 177.800 312.400 180.400 ;
        RECT 314.800 177.800 315.600 180.400 ;
        RECT 324.400 175.800 325.200 180.400 ;
        RECT 332.400 175.800 333.200 180.400 ;
        RECT 334.000 177.800 334.800 180.400 ;
        RECT 338.800 176.600 339.600 180.400 ;
        RECT 346.800 176.600 347.600 180.400 ;
        RECT 351.600 175.800 352.400 180.400 ;
        RECT 356.400 177.800 357.200 180.400 ;
        RECT 359.600 176.600 360.400 180.400 ;
        RECT 367.600 175.800 368.400 180.400 ;
        RECT 377.200 177.800 378.000 180.400 ;
        RECT 380.400 177.800 381.200 180.400 ;
        RECT 391.600 175.800 392.400 180.400 ;
        RECT 398.000 177.800 398.800 180.400 ;
        RECT 404.400 173.800 405.200 180.400 ;
        RECT 406.000 177.800 406.800 180.400 ;
        RECT 409.200 177.800 410.000 180.400 ;
        RECT 417.200 177.800 418.000 180.400 ;
        RECT 423.600 175.800 424.400 180.400 ;
        RECT 434.800 177.800 435.600 180.400 ;
        RECT 438.000 177.800 438.800 180.400 ;
        RECT 447.600 175.800 448.400 180.400 ;
        RECT 452.400 177.800 453.200 180.400 ;
        RECT 455.600 177.800 456.400 180.400 ;
        RECT 457.200 175.800 458.000 180.400 ;
        RECT 460.400 175.800 461.200 180.400 ;
        RECT 462.000 177.800 462.800 180.400 ;
        RECT 465.200 177.800 466.000 180.400 ;
        RECT 471.600 173.800 472.400 180.400 ;
        RECT 478.000 173.800 478.800 180.400 ;
        RECT 481.200 175.800 482.000 180.400 ;
        RECT 482.800 173.800 483.600 180.400 ;
        RECT 490.800 177.800 491.600 180.400 ;
        RECT 497.200 173.800 498.000 180.400 ;
        RECT 498.800 175.800 499.600 180.400 ;
        RECT 502.000 177.800 502.800 180.400 ;
        RECT 506.200 175.800 507.000 180.400 ;
        RECT 508.400 175.800 509.200 180.400 ;
        RECT 513.200 177.800 514.000 180.400 ;
        RECT 519.600 175.800 520.400 180.400 ;
        RECT 530.800 177.800 531.600 180.400 ;
        RECT 534.000 177.800 534.800 180.400 ;
        RECT 543.600 175.800 544.400 180.400 ;
        RECT 2.800 141.600 3.600 146.200 ;
        RECT 6.000 141.600 6.800 148.200 ;
        RECT 18.800 141.600 19.600 143.800 ;
        RECT 22.000 141.600 22.800 144.200 ;
        RECT 25.200 141.600 26.000 144.200 ;
        RECT 28.400 141.600 29.200 144.200 ;
        RECT 31.600 141.600 32.400 144.200 ;
        RECT 33.200 141.600 34.000 144.200 ;
        RECT 36.400 141.600 37.200 144.200 ;
        RECT 39.600 141.600 40.400 144.200 ;
        RECT 41.200 141.600 42.000 146.200 ;
        RECT 47.600 141.600 48.400 144.200 ;
        RECT 50.800 141.600 51.600 143.800 ;
        RECT 60.400 141.600 61.200 145.400 ;
        RECT 68.400 141.600 69.200 146.200 ;
        RECT 70.000 141.600 70.800 144.200 ;
        RECT 76.400 141.600 77.200 146.200 ;
        RECT 87.600 141.600 88.400 144.200 ;
        RECT 90.800 141.600 91.600 144.200 ;
        RECT 100.400 141.600 101.200 146.200 ;
        RECT 105.200 141.600 106.000 144.200 ;
        RECT 108.400 141.600 109.200 144.200 ;
        RECT 110.000 141.600 110.800 146.200 ;
        RECT 114.800 141.600 115.600 145.400 ;
        RECT 119.600 141.600 120.400 144.200 ;
        RECT 130.800 141.600 131.600 146.200 ;
        RECT 136.200 141.600 137.200 144.200 ;
        RECT 139.600 141.600 140.400 144.200 ;
        RECT 145.200 141.600 146.000 146.000 ;
        RECT 151.600 141.600 152.400 146.200 ;
        RECT 161.200 141.600 162.000 144.200 ;
        RECT 164.400 141.600 165.200 144.200 ;
        RECT 175.600 141.600 176.400 146.200 ;
        RECT 182.000 141.600 182.800 144.200 ;
        RECT 185.200 141.600 186.000 145.400 ;
        RECT 190.000 141.600 190.800 146.200 ;
        RECT 194.800 141.600 195.600 144.200 ;
        RECT 199.000 141.600 199.800 146.200 ;
        RECT 201.200 141.600 202.000 144.200 ;
        RECT 204.400 141.600 205.200 144.200 ;
        RECT 207.600 141.600 208.400 144.200 ;
        RECT 211.800 141.600 212.600 146.000 ;
        RECT 217.200 141.600 218.000 145.400 ;
        RECT 225.200 141.600 226.000 146.200 ;
        RECT 234.800 141.600 235.600 144.200 ;
        RECT 238.000 141.600 238.800 144.200 ;
        RECT 249.200 141.600 250.000 146.200 ;
        RECT 255.600 141.600 256.400 144.200 ;
        RECT 260.400 141.600 261.200 146.200 ;
        RECT 262.000 141.600 262.800 144.200 ;
        RECT 266.200 141.600 267.000 146.200 ;
        RECT 268.400 141.600 269.200 148.200 ;
        RECT 283.800 141.600 284.600 146.000 ;
        RECT 290.800 141.600 291.600 145.400 ;
        RECT 294.000 141.600 294.800 144.200 ;
        RECT 300.400 141.600 301.200 146.200 ;
        RECT 311.600 141.600 312.400 144.200 ;
        RECT 314.800 141.600 315.600 144.200 ;
        RECT 324.400 141.600 325.200 146.200 ;
        RECT 332.400 141.600 333.200 145.400 ;
        RECT 337.200 141.600 338.000 144.200 ;
        RECT 342.000 141.600 342.800 145.400 ;
        RECT 348.400 141.600 349.200 145.400 ;
        RECT 354.800 141.600 355.600 145.400 ;
        RECT 359.600 141.600 360.400 145.400 ;
        RECT 364.400 141.600 365.200 146.200 ;
        RECT 369.200 141.600 370.000 146.200 ;
        RECT 375.200 141.600 376.000 146.200 ;
        RECT 378.400 141.600 379.200 147.000 ;
        RECT 383.600 141.600 384.400 146.600 ;
        RECT 388.400 141.600 389.200 144.200 ;
        RECT 392.200 141.600 393.000 146.000 ;
        RECT 401.200 141.600 402.000 148.200 ;
        RECT 407.600 141.600 408.400 148.200 ;
        RECT 412.400 141.600 413.200 145.400 ;
        RECT 415.600 141.600 416.400 144.200 ;
        RECT 420.400 141.600 421.200 146.600 ;
        RECT 425.600 141.600 426.400 147.000 ;
        RECT 436.400 141.600 437.200 146.200 ;
        RECT 441.800 141.600 442.800 144.200 ;
        RECT 445.200 141.600 446.000 144.200 ;
        RECT 450.800 141.600 451.600 146.000 ;
        RECT 458.800 141.600 459.600 148.200 ;
        RECT 460.400 141.600 461.200 148.200 ;
        RECT 468.400 141.600 469.200 144.200 ;
        RECT 471.600 141.600 472.400 143.800 ;
        RECT 480.800 141.600 481.600 147.000 ;
        RECT 486.000 141.600 486.800 146.600 ;
        RECT 490.800 141.600 491.600 144.200 ;
        RECT 497.200 141.600 498.000 145.400 ;
        RECT 501.600 141.600 502.400 147.000 ;
        RECT 506.800 141.600 507.600 146.600 ;
        RECT 511.600 141.600 512.400 144.200 ;
        RECT 514.800 141.600 515.600 144.200 ;
        RECT 518.000 141.600 518.800 146.600 ;
        RECT 523.200 141.600 524.000 147.000 ;
        RECT 527.600 141.600 528.400 146.200 ;
        RECT 533.000 141.600 534.000 144.200 ;
        RECT 536.400 141.600 537.200 144.200 ;
        RECT 542.000 141.600 542.800 146.000 ;
        RECT 546.800 141.600 547.600 146.200 ;
        RECT 0.400 140.400 551.600 141.600 ;
        RECT 2.800 135.800 3.600 140.400 ;
        RECT 4.400 137.800 5.200 140.400 ;
        RECT 10.800 135.800 11.600 140.400 ;
        RECT 12.400 137.800 13.200 140.400 ;
        RECT 15.600 137.800 16.400 140.400 ;
        RECT 18.800 136.600 19.600 140.400 ;
        RECT 28.400 133.800 29.200 140.400 ;
        RECT 34.800 133.800 35.600 140.400 ;
        RECT 38.000 136.600 38.800 140.400 ;
        RECT 47.600 133.800 48.400 140.400 ;
        RECT 49.200 137.800 50.000 140.400 ;
        RECT 55.600 135.800 56.400 140.400 ;
        RECT 66.800 137.800 67.600 140.400 ;
        RECT 70.000 137.800 70.800 140.400 ;
        RECT 79.600 135.800 80.400 140.400 ;
        RECT 84.400 137.800 85.200 140.400 ;
        RECT 87.600 137.800 88.400 140.400 ;
        RECT 90.800 135.800 91.600 140.400 ;
        RECT 93.000 135.800 93.800 140.400 ;
        RECT 97.200 137.800 98.000 140.400 ;
        RECT 102.000 135.800 102.800 140.400 ;
        RECT 111.600 137.800 112.400 140.400 ;
        RECT 114.800 137.800 115.600 140.400 ;
        RECT 126.000 135.800 126.800 140.400 ;
        RECT 132.400 137.800 133.200 140.400 ;
        RECT 142.000 137.800 142.800 140.400 ;
        RECT 145.200 136.600 146.000 140.400 ;
        RECT 152.600 136.000 153.400 140.400 ;
        RECT 158.600 136.000 159.400 140.400 ;
        RECT 162.800 137.800 163.600 140.400 ;
        RECT 166.000 137.800 166.800 140.400 ;
        RECT 169.200 136.600 170.000 140.400 ;
        RECT 177.200 135.800 178.000 140.400 ;
        RECT 180.400 137.800 181.200 140.400 ;
        RECT 182.000 137.800 182.800 140.400 ;
        RECT 188.400 135.800 189.200 140.400 ;
        RECT 199.600 137.800 200.400 140.400 ;
        RECT 202.800 137.800 203.600 140.400 ;
        RECT 212.400 135.800 213.200 140.400 ;
        RECT 217.200 137.800 218.000 140.400 ;
        RECT 220.400 137.800 221.200 140.400 ;
        RECT 225.200 136.600 226.000 140.400 ;
        RECT 230.000 136.600 230.800 140.400 ;
        RECT 239.600 133.800 240.400 140.400 ;
        RECT 242.800 137.800 243.600 140.400 ;
        RECT 247.600 135.800 248.400 140.400 ;
        RECT 249.200 137.800 250.000 140.400 ;
        RECT 252.400 137.800 253.200 140.400 ;
        RECT 254.000 137.800 254.800 140.400 ;
        RECT 257.200 137.800 258.000 140.400 ;
        RECT 260.400 136.600 261.200 140.400 ;
        RECT 271.600 137.800 272.400 140.400 ;
        RECT 278.000 135.800 278.800 140.400 ;
        RECT 289.200 137.800 290.000 140.400 ;
        RECT 292.400 137.800 293.200 140.400 ;
        RECT 302.000 135.800 302.800 140.400 ;
        RECT 310.000 136.600 310.800 140.400 ;
        RECT 314.800 137.800 315.600 140.400 ;
        RECT 319.600 136.600 320.400 140.400 ;
        RECT 326.000 135.800 326.800 140.400 ;
        RECT 335.600 137.800 336.400 140.400 ;
        RECT 338.800 137.800 339.600 140.400 ;
        RECT 350.000 135.800 350.800 140.400 ;
        RECT 356.400 137.800 357.200 140.400 ;
        RECT 358.000 137.800 358.800 140.400 ;
        RECT 361.200 137.800 362.000 140.400 ;
        RECT 369.200 136.600 370.000 140.400 ;
        RECT 373.000 135.800 373.800 140.400 ;
        RECT 377.200 137.800 378.000 140.400 ;
        RECT 378.800 137.800 379.600 140.400 ;
        RECT 382.000 137.800 382.800 140.400 ;
        RECT 384.000 135.800 384.800 140.400 ;
        RECT 390.000 135.800 390.800 140.400 ;
        RECT 393.200 137.800 394.000 140.400 ;
        RECT 394.800 137.800 395.600 140.400 ;
        RECT 401.200 135.800 402.000 140.400 ;
        RECT 412.400 137.800 413.200 140.400 ;
        RECT 415.600 137.800 416.400 140.400 ;
        RECT 425.200 135.800 426.000 140.400 ;
        RECT 436.400 137.800 437.200 140.400 ;
        RECT 439.600 137.800 440.400 140.400 ;
        RECT 441.800 135.800 442.600 140.400 ;
        RECT 446.000 137.800 446.800 140.400 ;
        RECT 447.600 133.800 448.400 140.400 ;
        RECT 455.600 136.600 456.400 140.400 ;
        RECT 463.600 137.800 464.400 140.400 ;
        RECT 468.400 135.800 469.200 140.400 ;
        RECT 478.000 137.800 478.800 140.400 ;
        RECT 481.200 137.800 482.000 140.400 ;
        RECT 492.400 135.800 493.200 140.400 ;
        RECT 498.800 137.800 499.600 140.400 ;
        RECT 502.000 135.400 502.800 140.400 ;
        RECT 507.200 135.000 508.000 140.400 ;
        RECT 510.000 135.800 510.800 140.400 ;
        RECT 514.800 137.800 515.600 140.400 ;
        RECT 521.200 135.800 522.000 140.400 ;
        RECT 532.400 137.800 533.200 140.400 ;
        RECT 535.600 137.800 536.400 140.400 ;
        RECT 545.200 135.800 546.000 140.400 ;
        RECT 6.000 101.600 6.800 108.200 ;
        RECT 7.600 101.600 8.400 106.200 ;
        RECT 17.200 101.600 18.000 108.200 ;
        RECT 23.600 101.600 24.400 108.200 ;
        RECT 25.200 101.600 26.000 108.200 ;
        RECT 34.800 101.600 35.600 105.400 ;
        RECT 38.000 101.600 38.800 106.200 ;
        RECT 41.200 101.600 42.000 106.200 ;
        RECT 42.800 101.600 43.600 104.200 ;
        RECT 49.200 101.600 50.000 106.200 ;
        RECT 60.400 101.600 61.200 104.200 ;
        RECT 63.600 101.600 64.400 104.200 ;
        RECT 73.200 101.600 74.000 106.200 ;
        RECT 79.600 101.600 80.400 105.400 ;
        RECT 87.600 101.600 88.400 106.200 ;
        RECT 97.200 101.600 98.000 104.200 ;
        RECT 100.400 101.600 101.200 104.200 ;
        RECT 111.600 101.600 112.400 106.200 ;
        RECT 118.000 101.600 118.800 104.200 ;
        RECT 121.200 101.600 122.000 104.200 ;
        RECT 129.200 101.600 130.000 104.200 ;
        RECT 132.400 101.600 133.200 104.200 ;
        RECT 134.000 101.600 134.800 104.200 ;
        RECT 138.200 101.600 139.000 106.200 ;
        RECT 140.400 101.600 141.200 104.200 ;
        RECT 143.600 101.600 144.400 104.200 ;
        RECT 146.800 101.600 147.600 104.200 ;
        RECT 150.000 101.600 150.800 105.400 ;
        RECT 155.400 101.600 156.200 106.200 ;
        RECT 159.600 101.600 160.400 104.200 ;
        RECT 161.200 101.600 162.000 104.200 ;
        RECT 164.400 101.600 165.200 104.200 ;
        RECT 167.600 101.600 168.400 105.400 ;
        RECT 174.000 101.600 174.800 104.200 ;
        RECT 175.600 101.600 176.400 106.200 ;
        RECT 183.600 101.600 184.400 106.200 ;
        RECT 193.200 101.600 194.000 104.200 ;
        RECT 196.400 101.600 197.200 104.200 ;
        RECT 207.600 101.600 208.400 106.200 ;
        RECT 214.000 101.600 214.800 104.200 ;
        RECT 215.600 101.600 216.400 104.200 ;
        RECT 219.800 101.600 220.600 106.200 ;
        RECT 225.200 101.600 226.000 106.200 ;
        RECT 230.000 101.600 230.800 105.400 ;
        RECT 233.200 101.600 234.000 104.200 ;
        RECT 236.400 101.600 237.200 104.200 ;
        RECT 239.600 101.600 240.400 104.200 ;
        RECT 241.200 101.600 242.000 104.200 ;
        RECT 244.400 101.600 245.200 105.800 ;
        RECT 250.800 101.600 251.600 105.400 ;
        RECT 255.600 101.600 256.400 105.400 ;
        RECT 261.000 101.600 261.800 106.200 ;
        RECT 265.200 101.600 266.000 104.200 ;
        RECT 273.200 101.600 274.000 104.200 ;
        RECT 279.600 101.600 280.400 106.200 ;
        RECT 290.800 101.600 291.600 104.200 ;
        RECT 294.000 101.600 294.800 104.200 ;
        RECT 303.600 101.600 304.400 106.200 ;
        RECT 310.000 101.600 310.800 105.400 ;
        RECT 318.000 101.600 318.800 105.400 ;
        RECT 321.200 101.600 322.000 104.200 ;
        RECT 324.400 101.600 325.200 106.200 ;
        RECT 327.600 101.600 328.400 106.200 ;
        RECT 330.800 101.600 331.600 106.200 ;
        RECT 334.000 101.600 334.800 106.200 ;
        RECT 337.200 101.600 338.000 106.200 ;
        RECT 342.000 101.600 342.800 106.200 ;
        RECT 351.600 101.600 352.400 104.200 ;
        RECT 354.800 101.600 355.600 104.200 ;
        RECT 366.000 101.600 366.800 106.200 ;
        RECT 372.400 101.600 373.200 104.200 ;
        RECT 378.800 101.600 379.600 105.400 ;
        RECT 383.600 101.600 384.400 104.200 ;
        RECT 385.600 101.600 386.400 106.200 ;
        RECT 391.600 101.600 392.400 106.200 ;
        RECT 393.200 101.600 394.000 104.200 ;
        RECT 396.400 101.600 397.200 104.200 ;
        RECT 398.000 101.600 398.800 104.200 ;
        RECT 401.200 101.600 402.000 104.200 ;
        RECT 404.400 101.600 405.200 104.200 ;
        RECT 410.800 101.600 411.600 105.400 ;
        RECT 417.200 101.600 418.000 105.400 ;
        RECT 420.400 101.600 421.200 104.200 ;
        RECT 423.600 101.600 424.400 104.200 ;
        RECT 436.400 101.600 437.200 105.400 ;
        RECT 439.600 101.600 440.400 108.200 ;
        RECT 446.600 101.600 447.400 106.200 ;
        RECT 450.800 101.600 451.600 104.200 ;
        RECT 455.600 101.600 456.400 106.200 ;
        RECT 458.800 101.600 459.600 105.400 ;
        RECT 463.600 101.600 464.400 104.200 ;
        RECT 466.800 101.600 467.600 104.200 ;
        RECT 468.400 101.600 469.200 106.200 ;
        RECT 473.200 101.600 474.000 106.200 ;
        RECT 476.800 101.600 477.600 106.200 ;
        RECT 482.800 101.600 483.600 106.200 ;
        RECT 486.000 101.600 486.800 106.600 ;
        RECT 491.200 101.600 492.000 107.000 ;
        RECT 494.000 101.600 494.800 106.200 ;
        RECT 500.400 101.600 501.200 105.400 ;
        RECT 508.400 101.600 509.200 106.200 ;
        RECT 513.200 101.600 514.000 105.400 ;
        RECT 516.400 101.600 517.200 104.200 ;
        RECT 522.800 101.600 523.600 106.200 ;
        RECT 534.000 101.600 534.800 104.200 ;
        RECT 537.200 101.600 538.000 104.200 ;
        RECT 546.800 101.600 547.600 106.200 ;
        RECT 0.400 100.400 551.600 101.600 ;
        RECT 1.200 95.800 2.000 100.400 ;
        RECT 6.000 97.800 6.800 100.400 ;
        RECT 9.200 97.800 10.000 100.400 ;
        RECT 15.600 93.800 16.400 100.400 ;
        RECT 22.000 93.800 22.800 100.400 ;
        RECT 25.200 96.600 26.000 100.400 ;
        RECT 30.000 95.800 30.800 100.400 ;
        RECT 34.800 95.800 35.600 100.400 ;
        RECT 41.200 96.600 42.000 100.400 ;
        RECT 49.200 95.800 50.000 100.400 ;
        RECT 58.800 97.800 59.600 100.400 ;
        RECT 62.000 97.800 62.800 100.400 ;
        RECT 73.200 95.800 74.000 100.400 ;
        RECT 79.600 97.800 80.400 100.400 ;
        RECT 84.400 96.600 85.200 100.400 ;
        RECT 87.600 97.800 88.400 100.400 ;
        RECT 90.800 97.800 91.600 100.400 ;
        RECT 92.400 97.800 93.200 100.400 ;
        RECT 96.600 95.800 97.400 100.400 ;
        RECT 102.000 95.800 102.800 100.400 ;
        RECT 111.600 97.800 112.400 100.400 ;
        RECT 114.800 97.800 115.600 100.400 ;
        RECT 126.000 95.800 126.800 100.400 ;
        RECT 132.400 97.800 133.200 100.400 ;
        RECT 142.000 97.800 142.800 100.400 ;
        RECT 143.600 97.800 144.400 100.400 ;
        RECT 146.800 96.200 147.600 100.400 ;
        RECT 153.200 96.600 154.000 100.400 ;
        RECT 158.000 95.800 158.800 100.400 ;
        RECT 163.400 97.800 164.400 100.400 ;
        RECT 166.800 97.800 167.600 100.400 ;
        RECT 172.400 96.000 173.200 100.400 ;
        RECT 177.200 95.800 178.000 100.400 ;
        RECT 182.000 95.800 182.800 100.400 ;
        RECT 185.200 97.800 186.000 100.400 ;
        RECT 189.000 95.800 189.800 100.400 ;
        RECT 193.200 97.800 194.000 100.400 ;
        RECT 194.800 95.800 195.600 100.400 ;
        RECT 202.800 95.800 203.600 100.400 ;
        RECT 207.600 96.600 208.400 100.400 ;
        RECT 212.400 97.800 213.200 100.400 ;
        RECT 214.000 95.800 214.800 100.400 ;
        RECT 218.800 97.800 219.600 100.400 ;
        RECT 222.000 97.800 222.800 100.400 ;
        RECT 223.600 95.800 224.400 100.400 ;
        RECT 228.400 97.800 229.200 100.400 ;
        RECT 231.600 97.800 232.400 100.400 ;
        RECT 235.800 95.800 236.600 100.400 ;
        RECT 239.600 96.600 240.400 100.400 ;
        RECT 246.000 97.800 246.800 100.400 ;
        RECT 249.200 98.200 250.000 100.400 ;
        RECT 257.200 97.800 258.000 100.400 ;
        RECT 260.400 97.800 261.200 100.400 ;
        RECT 268.400 97.800 269.200 100.400 ;
        RECT 274.800 95.800 275.600 100.400 ;
        RECT 286.000 97.800 286.800 100.400 ;
        RECT 289.200 97.800 290.000 100.400 ;
        RECT 298.800 95.800 299.600 100.400 ;
        RECT 303.600 97.800 304.400 100.400 ;
        RECT 306.800 97.800 307.600 100.400 ;
        RECT 313.200 95.800 314.000 100.400 ;
        RECT 324.400 97.800 325.200 100.400 ;
        RECT 327.600 97.800 328.400 100.400 ;
        RECT 337.200 95.800 338.000 100.400 ;
        RECT 343.600 96.600 344.400 100.400 ;
        RECT 351.600 96.600 352.400 100.400 ;
        RECT 358.000 95.800 358.800 100.400 ;
        RECT 367.600 97.800 368.400 100.400 ;
        RECT 370.800 97.800 371.600 100.400 ;
        RECT 382.000 95.800 382.800 100.400 ;
        RECT 388.400 97.800 389.200 100.400 ;
        RECT 393.200 95.800 394.000 100.400 ;
        RECT 398.000 95.800 398.800 100.400 ;
        RECT 399.600 95.800 400.400 100.400 ;
        RECT 404.400 95.800 405.200 100.400 ;
        RECT 412.400 96.600 413.200 100.400 ;
        RECT 415.600 97.800 416.400 100.400 ;
        RECT 420.400 95.800 421.200 100.400 ;
        RECT 430.000 97.800 430.800 100.400 ;
        RECT 433.200 97.800 434.000 100.400 ;
        RECT 437.400 95.800 438.200 100.400 ;
        RECT 439.600 93.800 440.400 100.400 ;
        RECT 446.000 95.800 446.800 100.400 ;
        RECT 452.400 95.800 453.200 100.400 ;
        RECT 456.800 95.000 457.600 100.400 ;
        RECT 462.000 95.400 462.800 100.400 ;
        RECT 465.600 95.800 466.400 100.400 ;
        RECT 471.600 95.800 472.400 100.400 ;
        RECT 473.200 95.800 474.000 100.400 ;
        RECT 479.200 95.800 480.000 100.400 ;
        RECT 481.200 97.800 482.000 100.400 ;
        RECT 487.600 95.800 488.400 100.400 ;
        RECT 498.800 97.800 499.600 100.400 ;
        RECT 502.000 97.800 502.800 100.400 ;
        RECT 511.600 95.800 512.400 100.400 ;
        RECT 516.400 97.800 517.200 100.400 ;
        RECT 522.800 95.800 523.600 100.400 ;
        RECT 534.000 97.800 534.800 100.400 ;
        RECT 537.200 97.800 538.000 100.400 ;
        RECT 546.800 95.800 547.600 100.400 ;
        RECT 1.200 61.600 2.000 64.200 ;
        RECT 4.400 61.600 5.200 64.200 ;
        RECT 6.000 61.600 6.800 64.200 ;
        RECT 9.200 61.600 10.000 64.200 ;
        RECT 12.400 61.600 13.200 64.200 ;
        RECT 14.000 61.600 14.800 64.200 ;
        RECT 17.200 61.600 18.000 64.200 ;
        RECT 18.800 61.600 19.600 64.200 ;
        RECT 22.000 61.600 22.800 64.200 ;
        RECT 25.200 61.600 26.000 64.200 ;
        RECT 26.800 61.600 27.600 64.200 ;
        RECT 30.000 61.600 30.800 64.200 ;
        RECT 31.600 61.600 32.400 64.200 ;
        RECT 34.800 61.600 35.600 64.200 ;
        RECT 39.600 61.600 40.400 66.200 ;
        RECT 42.800 61.600 43.600 64.200 ;
        RECT 46.000 61.600 46.800 65.400 ;
        RECT 54.000 61.600 54.800 65.400 ;
        RECT 62.000 61.600 62.800 66.200 ;
        RECT 63.600 61.600 64.400 66.200 ;
        RECT 66.800 61.600 67.600 66.200 ;
        RECT 70.000 61.600 70.800 66.200 ;
        RECT 73.200 61.600 74.000 66.200 ;
        RECT 76.400 61.600 77.200 66.200 ;
        RECT 78.000 61.600 78.800 68.200 ;
        RECT 89.200 61.600 90.000 68.200 ;
        RECT 90.800 61.600 91.600 64.200 ;
        RECT 97.200 61.600 98.000 66.200 ;
        RECT 108.400 61.600 109.200 64.200 ;
        RECT 111.600 61.600 112.400 64.200 ;
        RECT 121.200 61.600 122.000 66.200 ;
        RECT 132.400 61.600 133.200 64.200 ;
        RECT 138.800 61.600 139.600 66.200 ;
        RECT 150.000 61.600 150.800 64.200 ;
        RECT 153.200 61.600 154.000 64.200 ;
        RECT 162.800 61.600 163.600 66.200 ;
        RECT 169.200 61.600 170.000 66.200 ;
        RECT 175.600 61.600 176.400 66.200 ;
        RECT 185.200 61.600 186.000 64.200 ;
        RECT 188.400 61.600 189.200 64.200 ;
        RECT 199.600 61.600 200.400 66.200 ;
        RECT 206.000 61.600 206.800 64.200 ;
        RECT 207.600 61.600 208.400 64.200 ;
        RECT 214.000 61.600 214.800 66.200 ;
        RECT 225.200 61.600 226.000 64.200 ;
        RECT 228.400 61.600 229.200 64.200 ;
        RECT 238.000 61.600 238.800 66.200 ;
        RECT 244.400 61.600 245.200 66.200 ;
        RECT 247.600 61.600 248.400 64.200 ;
        RECT 252.400 61.600 253.200 65.400 ;
        RECT 260.400 61.600 261.200 65.400 ;
        RECT 263.600 61.600 264.400 64.200 ;
        RECT 273.200 61.600 274.000 64.200 ;
        RECT 279.600 61.600 280.400 66.200 ;
        RECT 290.800 61.600 291.600 64.200 ;
        RECT 294.000 61.600 294.800 64.200 ;
        RECT 303.600 61.600 304.400 66.200 ;
        RECT 310.000 61.600 310.800 65.400 ;
        RECT 318.000 61.600 318.800 65.400 ;
        RECT 322.800 61.600 323.600 66.200 ;
        RECT 330.800 61.600 331.600 65.400 ;
        RECT 335.600 61.600 336.400 64.200 ;
        RECT 337.200 61.600 338.000 64.200 ;
        RECT 343.600 61.600 344.400 66.200 ;
        RECT 354.800 61.600 355.600 64.200 ;
        RECT 358.000 61.600 358.800 64.200 ;
        RECT 367.600 61.600 368.400 66.200 ;
        RECT 374.000 61.600 374.800 65.400 ;
        RECT 383.600 61.600 384.400 65.400 ;
        RECT 388.400 61.600 389.200 65.400 ;
        RECT 394.800 61.600 395.600 64.200 ;
        RECT 399.600 61.600 400.400 66.200 ;
        RECT 401.200 61.600 402.000 64.200 ;
        RECT 404.400 61.600 405.200 64.200 ;
        RECT 406.000 61.600 406.800 64.200 ;
        RECT 415.600 61.600 416.400 64.200 ;
        RECT 422.000 61.600 422.800 66.200 ;
        RECT 433.200 61.600 434.000 64.200 ;
        RECT 436.400 61.600 437.200 64.200 ;
        RECT 446.000 61.600 446.800 66.200 ;
        RECT 454.000 61.600 454.800 65.400 ;
        RECT 458.800 61.600 459.600 64.200 ;
        RECT 460.400 61.600 461.200 64.200 ;
        RECT 464.600 61.600 465.400 66.200 ;
        RECT 470.000 61.600 470.800 66.200 ;
        RECT 471.600 61.600 472.400 64.200 ;
        RECT 475.800 61.600 476.600 66.200 ;
        RECT 479.200 61.600 480.000 67.000 ;
        RECT 484.400 61.600 485.200 66.600 ;
        RECT 487.600 61.600 488.400 66.200 ;
        RECT 494.000 61.600 494.800 65.400 ;
        RECT 502.000 61.600 502.800 65.400 ;
        RECT 508.400 61.600 509.200 66.200 ;
        RECT 513.200 61.600 514.000 66.200 ;
        RECT 514.800 61.600 515.600 64.200 ;
        RECT 521.200 61.600 522.000 66.200 ;
        RECT 532.400 61.600 533.200 64.200 ;
        RECT 535.600 61.600 536.400 64.200 ;
        RECT 545.200 61.600 546.000 66.200 ;
        RECT 0.400 60.400 551.600 61.600 ;
        RECT 1.200 57.800 2.000 60.400 ;
        RECT 4.400 55.800 5.200 60.400 ;
        RECT 9.200 57.800 10.000 60.400 ;
        RECT 12.400 55.800 13.200 60.400 ;
        RECT 18.800 56.600 19.600 60.400 ;
        RECT 26.800 56.600 27.600 60.400 ;
        RECT 33.200 55.800 34.000 60.400 ;
        RECT 39.600 57.800 40.400 60.400 ;
        RECT 44.400 55.800 45.200 60.400 ;
        RECT 54.000 57.800 54.800 60.400 ;
        RECT 57.200 57.800 58.000 60.400 ;
        RECT 68.400 55.800 69.200 60.400 ;
        RECT 74.800 57.800 75.600 60.400 ;
        RECT 76.400 55.800 77.200 60.400 ;
        RECT 79.600 55.800 80.400 60.400 ;
        RECT 82.800 55.800 83.600 60.400 ;
        RECT 86.000 55.800 86.800 60.400 ;
        RECT 89.200 55.800 90.000 60.400 ;
        RECT 94.000 55.800 94.800 60.400 ;
        RECT 103.600 57.800 104.400 60.400 ;
        RECT 106.800 57.800 107.600 60.400 ;
        RECT 118.000 55.800 118.800 60.400 ;
        RECT 124.400 57.800 125.200 60.400 ;
        RECT 132.400 57.800 133.200 60.400 ;
        RECT 135.600 57.800 136.400 60.400 ;
        RECT 138.800 57.800 139.600 60.400 ;
        RECT 140.400 57.800 141.200 60.400 ;
        RECT 143.600 57.800 144.400 60.400 ;
        RECT 148.400 55.800 149.200 60.400 ;
        RECT 150.000 55.800 150.800 60.400 ;
        RECT 154.800 57.800 155.600 60.400 ;
        RECT 158.000 57.800 158.800 60.400 ;
        RECT 162.800 55.800 163.600 60.400 ;
        RECT 166.000 57.800 166.800 60.400 ;
        RECT 167.600 57.800 168.400 60.400 ;
        RECT 170.800 57.800 171.600 60.400 ;
        RECT 172.400 55.800 173.200 60.400 ;
        RECT 175.600 55.800 176.400 60.400 ;
        RECT 180.400 55.800 181.200 60.400 ;
        RECT 190.000 57.800 190.800 60.400 ;
        RECT 193.200 57.800 194.000 60.400 ;
        RECT 204.400 55.800 205.200 60.400 ;
        RECT 210.800 57.800 211.600 60.400 ;
        RECT 214.000 56.600 214.800 60.400 ;
        RECT 222.000 56.600 222.800 60.400 ;
        RECT 226.800 57.800 227.600 60.400 ;
        RECT 230.000 56.600 230.800 60.400 ;
        RECT 234.800 57.800 235.600 60.400 ;
        RECT 241.200 55.800 242.000 60.400 ;
        RECT 252.400 57.800 253.200 60.400 ;
        RECT 255.600 57.800 256.400 60.400 ;
        RECT 265.200 55.800 266.000 60.400 ;
        RECT 271.600 55.800 272.400 60.400 ;
        RECT 284.400 55.800 285.200 60.400 ;
        RECT 294.000 57.800 294.800 60.400 ;
        RECT 297.200 57.800 298.000 60.400 ;
        RECT 308.400 55.800 309.200 60.400 ;
        RECT 314.800 57.800 315.600 60.400 ;
        RECT 316.400 57.800 317.200 60.400 ;
        RECT 322.800 55.800 323.600 60.400 ;
        RECT 332.400 57.800 333.200 60.400 ;
        RECT 335.600 57.800 336.400 60.400 ;
        RECT 346.800 55.800 347.600 60.400 ;
        RECT 353.200 57.800 354.000 60.400 ;
        RECT 354.800 57.800 355.600 60.400 ;
        RECT 358.000 57.800 358.800 60.400 ;
        RECT 359.600 57.800 360.400 60.400 ;
        RECT 364.400 56.600 365.200 60.400 ;
        RECT 372.400 55.800 373.200 60.400 ;
        RECT 377.200 55.800 378.000 60.400 ;
        RECT 386.800 57.800 387.600 60.400 ;
        RECT 390.000 57.800 390.800 60.400 ;
        RECT 401.200 55.800 402.000 60.400 ;
        RECT 407.600 57.800 408.400 60.400 ;
        RECT 410.400 55.000 411.200 60.400 ;
        RECT 415.600 55.400 416.400 60.400 ;
        RECT 420.400 57.800 421.200 60.400 ;
        RECT 429.600 55.000 430.400 60.400 ;
        RECT 434.800 55.400 435.600 60.400 ;
        RECT 439.600 57.800 440.400 60.400 ;
        RECT 441.200 57.800 442.000 60.400 ;
        RECT 447.600 55.800 448.400 60.400 ;
        RECT 458.800 57.800 459.600 60.400 ;
        RECT 462.000 57.800 462.800 60.400 ;
        RECT 471.600 55.800 472.400 60.400 ;
        RECT 476.400 55.800 477.200 60.400 ;
        RECT 482.400 55.000 483.200 60.400 ;
        RECT 487.600 55.400 488.400 60.400 ;
        RECT 492.400 55.400 493.200 60.400 ;
        RECT 497.600 55.000 498.400 60.400 ;
        RECT 502.000 56.600 502.800 60.400 ;
        RECT 508.400 56.600 509.200 60.400 ;
        RECT 513.200 57.800 514.000 60.400 ;
        RECT 519.600 55.800 520.400 60.400 ;
        RECT 530.800 57.800 531.600 60.400 ;
        RECT 534.000 57.800 534.800 60.400 ;
        RECT 543.600 55.800 544.400 60.400 ;
        RECT 1.200 21.600 2.000 24.200 ;
        RECT 7.600 21.600 8.400 26.200 ;
        RECT 18.800 21.600 19.600 24.200 ;
        RECT 22.000 21.600 22.800 24.200 ;
        RECT 31.600 21.600 32.400 26.200 ;
        RECT 36.400 21.600 37.200 24.200 ;
        RECT 42.800 21.600 43.600 26.200 ;
        RECT 54.000 21.600 54.800 24.200 ;
        RECT 57.200 21.600 58.000 24.200 ;
        RECT 66.800 21.600 67.600 26.200 ;
        RECT 73.200 21.600 74.000 26.200 ;
        RECT 76.400 21.600 77.200 26.200 ;
        RECT 79.600 21.600 80.400 26.200 ;
        RECT 82.800 21.600 83.600 26.200 ;
        RECT 86.000 21.600 86.800 26.200 ;
        RECT 89.200 21.600 90.000 26.200 ;
        RECT 94.000 21.600 94.800 26.200 ;
        RECT 103.600 21.600 104.400 24.200 ;
        RECT 106.800 21.600 107.600 24.200 ;
        RECT 118.000 21.600 118.800 26.200 ;
        RECT 124.400 21.600 125.200 24.200 ;
        RECT 132.400 21.600 133.200 24.200 ;
        RECT 138.800 21.600 139.600 26.200 ;
        RECT 150.000 21.600 150.800 24.200 ;
        RECT 153.200 21.600 154.000 24.200 ;
        RECT 162.800 21.600 163.600 26.200 ;
        RECT 174.000 24.300 174.800 26.200 ;
        RECT 175.600 24.300 176.400 24.400 ;
        RECT 167.600 21.600 168.400 24.200 ;
        RECT 174.000 23.700 176.400 24.300 ;
        RECT 174.000 21.600 174.800 23.700 ;
        RECT 175.600 23.600 176.400 23.700 ;
        RECT 185.200 21.600 186.000 24.200 ;
        RECT 188.400 21.600 189.200 24.200 ;
        RECT 198.000 21.600 198.800 26.200 ;
        RECT 202.800 21.600 203.600 26.200 ;
        RECT 210.800 21.600 211.600 25.400 ;
        RECT 214.000 21.600 214.800 24.200 ;
        RECT 218.800 21.600 219.600 25.400 ;
        RECT 225.200 21.600 226.000 25.400 ;
        RECT 230.000 21.600 230.800 24.200 ;
        RECT 236.400 21.600 237.200 26.200 ;
        RECT 247.600 21.600 248.400 24.200 ;
        RECT 250.800 21.600 251.600 24.200 ;
        RECT 260.400 21.600 261.200 26.200 ;
        RECT 265.200 21.600 266.000 24.200 ;
        RECT 270.000 21.600 270.800 25.400 ;
        RECT 284.400 21.600 285.200 25.400 ;
        RECT 287.600 21.600 288.400 24.200 ;
        RECT 294.000 21.600 294.800 26.200 ;
        RECT 305.200 21.600 306.000 24.200 ;
        RECT 308.400 21.600 309.200 24.200 ;
        RECT 318.000 21.600 318.800 26.200 ;
        RECT 322.800 21.600 323.600 24.200 ;
        RECT 329.200 21.600 330.000 26.200 ;
        RECT 340.400 21.600 341.200 24.200 ;
        RECT 343.600 21.600 344.400 24.200 ;
        RECT 353.200 21.600 354.000 26.200 ;
        RECT 358.000 21.600 358.800 26.200 ;
        RECT 361.200 21.600 362.000 26.200 ;
        RECT 364.400 21.600 365.200 26.200 ;
        RECT 367.600 21.600 368.400 26.200 ;
        RECT 370.800 21.600 371.600 26.200 ;
        RECT 375.600 21.600 376.400 26.200 ;
        RECT 385.200 21.600 386.000 24.200 ;
        RECT 388.400 21.600 389.200 24.200 ;
        RECT 399.600 21.600 400.400 26.200 ;
        RECT 406.000 21.600 406.800 24.200 ;
        RECT 407.600 21.600 408.400 24.200 ;
        RECT 420.400 21.600 421.200 26.200 ;
        RECT 430.000 21.600 430.800 24.200 ;
        RECT 433.200 21.600 434.000 24.200 ;
        RECT 444.400 21.600 445.200 26.200 ;
        RECT 450.800 21.600 451.600 24.200 ;
        RECT 454.000 21.600 454.800 26.000 ;
        RECT 459.600 21.600 460.400 24.200 ;
        RECT 462.800 21.600 463.800 24.200 ;
        RECT 468.400 21.600 469.200 26.200 ;
        RECT 471.600 21.600 472.400 24.200 ;
        RECT 476.400 21.600 477.200 25.400 ;
        RECT 481.200 21.600 482.000 24.200 ;
        RECT 487.600 21.600 488.400 26.200 ;
        RECT 498.800 21.600 499.600 24.200 ;
        RECT 502.000 21.600 502.800 24.200 ;
        RECT 511.600 21.600 512.400 26.200 ;
        RECT 517.600 21.600 518.400 27.000 ;
        RECT 522.800 21.600 523.600 26.600 ;
        RECT 527.600 21.600 528.400 26.600 ;
        RECT 532.800 21.600 533.600 27.000 ;
        RECT 535.600 21.600 536.400 26.200 ;
        RECT 538.800 21.600 539.600 26.200 ;
        RECT 542.000 21.600 542.800 26.200 ;
        RECT 545.200 21.600 546.000 26.200 ;
        RECT 548.400 21.600 549.200 26.200 ;
        RECT 0.400 20.400 551.600 21.600 ;
        RECT 1.200 17.800 2.000 20.400 ;
        RECT 7.600 15.800 8.400 20.400 ;
        RECT 18.800 17.800 19.600 20.400 ;
        RECT 22.000 17.800 22.800 20.400 ;
        RECT 31.600 15.800 32.400 20.400 ;
        RECT 39.600 15.800 40.400 20.400 ;
        RECT 49.200 17.800 50.000 20.400 ;
        RECT 52.400 17.800 53.200 20.400 ;
        RECT 63.600 15.800 64.400 20.400 ;
        RECT 70.000 17.800 70.800 20.400 ;
        RECT 73.800 16.000 74.600 20.400 ;
        RECT 80.600 16.000 81.400 20.400 ;
        RECT 87.600 15.800 88.400 20.400 ;
        RECT 97.200 17.800 98.000 20.400 ;
        RECT 100.400 17.800 101.200 20.400 ;
        RECT 111.600 15.800 112.400 20.400 ;
        RECT 118.000 17.800 118.800 20.400 ;
        RECT 119.600 17.800 120.400 20.400 ;
        RECT 122.800 17.800 123.600 20.400 ;
        RECT 134.000 16.600 134.800 20.400 ;
        RECT 137.200 17.800 138.000 20.400 ;
        RECT 143.600 15.800 144.400 20.400 ;
        RECT 154.800 17.800 155.600 20.400 ;
        RECT 158.000 17.800 158.800 20.400 ;
        RECT 167.600 15.800 168.400 20.400 ;
        RECT 174.000 15.800 174.800 20.400 ;
        RECT 178.800 15.800 179.600 20.400 ;
        RECT 185.200 15.800 186.000 20.400 ;
        RECT 194.800 17.800 195.600 20.400 ;
        RECT 198.000 17.800 198.800 20.400 ;
        RECT 209.200 15.800 210.000 20.400 ;
        RECT 215.600 17.800 216.400 20.400 ;
        RECT 217.200 17.800 218.000 20.400 ;
        RECT 222.000 16.600 222.800 20.400 ;
        RECT 228.400 16.600 229.200 20.400 ;
        RECT 233.200 15.800 234.000 20.400 ;
        RECT 239.600 16.600 240.400 20.400 ;
        RECT 246.000 16.600 246.800 20.400 ;
        RECT 254.000 16.600 254.800 20.400 ;
        RECT 260.400 16.600 261.200 20.400 ;
        RECT 265.200 17.800 266.000 20.400 ;
        RECT 266.800 17.800 267.600 20.400 ;
        RECT 271.600 16.600 272.400 20.400 ;
        RECT 284.400 16.600 285.200 20.400 ;
        RECT 289.200 17.800 290.000 20.400 ;
        RECT 295.600 15.800 296.400 20.400 ;
        RECT 306.800 17.800 307.600 20.400 ;
        RECT 310.000 17.800 310.800 20.400 ;
        RECT 319.600 15.800 320.400 20.400 ;
        RECT 327.000 16.000 327.800 20.400 ;
        RECT 333.400 16.000 334.200 20.400 ;
        RECT 337.200 17.800 338.000 20.400 ;
        RECT 343.600 15.800 344.400 20.400 ;
        RECT 354.800 17.800 355.600 20.400 ;
        RECT 358.000 17.800 358.800 20.400 ;
        RECT 367.600 15.800 368.400 20.400 ;
        RECT 374.000 15.800 374.800 20.400 ;
        RECT 378.800 16.000 379.600 20.400 ;
        RECT 384.400 17.800 385.200 20.400 ;
        RECT 387.600 17.800 388.600 20.400 ;
        RECT 393.200 15.800 394.000 20.400 ;
        RECT 399.600 15.800 400.400 20.400 ;
        RECT 409.200 17.800 410.000 20.400 ;
        RECT 412.400 17.800 413.200 20.400 ;
        RECT 423.600 15.800 424.400 20.400 ;
        RECT 430.000 17.800 430.800 20.400 ;
        RECT 439.600 15.800 440.400 20.400 ;
        RECT 445.000 17.800 446.000 20.400 ;
        RECT 448.400 17.800 449.200 20.400 ;
        RECT 454.000 16.000 454.800 20.400 ;
        RECT 458.800 15.800 459.600 20.400 ;
        RECT 463.600 15.800 464.400 20.400 ;
        RECT 470.000 15.800 470.800 20.400 ;
        RECT 479.600 17.800 480.400 20.400 ;
        RECT 482.800 17.800 483.600 20.400 ;
        RECT 494.000 15.800 494.800 20.400 ;
        RECT 500.400 17.800 501.200 20.400 ;
        RECT 502.000 17.800 502.800 20.400 ;
        RECT 508.400 15.800 509.200 20.400 ;
        RECT 518.000 17.800 518.800 20.400 ;
        RECT 521.200 17.800 522.000 20.400 ;
        RECT 532.400 15.800 533.200 20.400 ;
        RECT 538.800 17.800 539.600 20.400 ;
        RECT 542.000 15.800 542.800 20.400 ;
        RECT 546.800 15.800 547.600 20.400 ;
        RECT 175.600 12.300 176.400 13.200 ;
        RECT 177.200 12.300 178.000 13.200 ;
        RECT 175.600 11.700 178.000 12.300 ;
        RECT 175.600 11.600 176.400 11.700 ;
        RECT 177.200 11.600 178.000 11.700 ;
      LAYER via1 ;
        RECT 272.300 380.600 273.100 381.400 ;
        RECT 273.300 380.600 274.100 381.400 ;
        RECT 274.300 380.600 275.100 381.400 ;
        RECT 275.300 380.600 276.100 381.400 ;
        RECT 276.300 380.600 277.100 381.400 ;
        RECT 277.300 380.600 278.100 381.400 ;
        RECT 272.300 340.600 273.100 341.400 ;
        RECT 273.300 340.600 274.100 341.400 ;
        RECT 274.300 340.600 275.100 341.400 ;
        RECT 275.300 340.600 276.100 341.400 ;
        RECT 276.300 340.600 277.100 341.400 ;
        RECT 277.300 340.600 278.100 341.400 ;
        RECT 272.300 300.600 273.100 301.400 ;
        RECT 273.300 300.600 274.100 301.400 ;
        RECT 274.300 300.600 275.100 301.400 ;
        RECT 275.300 300.600 276.100 301.400 ;
        RECT 276.300 300.600 277.100 301.400 ;
        RECT 277.300 300.600 278.100 301.400 ;
        RECT 272.300 260.600 273.100 261.400 ;
        RECT 273.300 260.600 274.100 261.400 ;
        RECT 274.300 260.600 275.100 261.400 ;
        RECT 275.300 260.600 276.100 261.400 ;
        RECT 276.300 260.600 277.100 261.400 ;
        RECT 277.300 260.600 278.100 261.400 ;
        RECT 272.300 220.600 273.100 221.400 ;
        RECT 273.300 220.600 274.100 221.400 ;
        RECT 274.300 220.600 275.100 221.400 ;
        RECT 275.300 220.600 276.100 221.400 ;
        RECT 276.300 220.600 277.100 221.400 ;
        RECT 277.300 220.600 278.100 221.400 ;
        RECT 272.300 180.600 273.100 181.400 ;
        RECT 273.300 180.600 274.100 181.400 ;
        RECT 274.300 180.600 275.100 181.400 ;
        RECT 275.300 180.600 276.100 181.400 ;
        RECT 276.300 180.600 277.100 181.400 ;
        RECT 277.300 180.600 278.100 181.400 ;
        RECT 272.300 140.600 273.100 141.400 ;
        RECT 273.300 140.600 274.100 141.400 ;
        RECT 274.300 140.600 275.100 141.400 ;
        RECT 275.300 140.600 276.100 141.400 ;
        RECT 276.300 140.600 277.100 141.400 ;
        RECT 277.300 140.600 278.100 141.400 ;
        RECT 272.300 100.600 273.100 101.400 ;
        RECT 273.300 100.600 274.100 101.400 ;
        RECT 274.300 100.600 275.100 101.400 ;
        RECT 275.300 100.600 276.100 101.400 ;
        RECT 276.300 100.600 277.100 101.400 ;
        RECT 277.300 100.600 278.100 101.400 ;
        RECT 272.300 60.600 273.100 61.400 ;
        RECT 273.300 60.600 274.100 61.400 ;
        RECT 274.300 60.600 275.100 61.400 ;
        RECT 275.300 60.600 276.100 61.400 ;
        RECT 276.300 60.600 277.100 61.400 ;
        RECT 277.300 60.600 278.100 61.400 ;
        RECT 272.300 20.600 273.100 21.400 ;
        RECT 273.300 20.600 274.100 21.400 ;
        RECT 274.300 20.600 275.100 21.400 ;
        RECT 275.300 20.600 276.100 21.400 ;
        RECT 276.300 20.600 277.100 21.400 ;
        RECT 277.300 20.600 278.100 21.400 ;
      LAYER metal2 ;
        RECT 274.600 381.400 275.800 381.600 ;
        RECT 272.300 380.600 278.100 381.400 ;
        RECT 274.600 380.400 275.800 380.600 ;
        RECT 274.600 341.400 275.800 341.600 ;
        RECT 272.300 340.600 278.100 341.400 ;
        RECT 274.600 340.400 275.800 340.600 ;
        RECT 274.600 301.400 275.800 301.600 ;
        RECT 272.300 300.600 278.100 301.400 ;
        RECT 274.600 300.400 275.800 300.600 ;
        RECT 274.600 261.400 275.800 261.600 ;
        RECT 272.300 260.600 278.100 261.400 ;
        RECT 274.600 260.400 275.800 260.600 ;
        RECT 274.600 221.400 275.800 221.600 ;
        RECT 272.300 220.600 278.100 221.400 ;
        RECT 274.600 220.400 275.800 220.600 ;
        RECT 274.600 181.400 275.800 181.600 ;
        RECT 272.300 180.600 278.100 181.400 ;
        RECT 274.600 180.400 275.800 180.600 ;
        RECT 274.600 141.400 275.800 141.600 ;
        RECT 272.300 140.600 278.100 141.400 ;
        RECT 274.600 140.400 275.800 140.600 ;
        RECT 274.600 101.400 275.800 101.600 ;
        RECT 272.300 100.600 278.100 101.400 ;
        RECT 274.600 100.400 275.800 100.600 ;
        RECT 274.600 61.400 275.800 61.600 ;
        RECT 272.300 60.600 278.100 61.400 ;
        RECT 274.600 60.400 275.800 60.600 ;
        RECT 175.600 23.600 176.400 24.400 ;
        RECT 175.700 12.400 176.300 23.600 ;
        RECT 274.600 21.400 275.800 21.600 ;
        RECT 272.300 20.600 278.100 21.400 ;
        RECT 274.600 20.400 275.800 20.600 ;
        RECT 175.600 11.600 176.400 12.400 ;
      LAYER via2 ;
        RECT 273.300 380.600 274.100 381.400 ;
        RECT 274.300 380.600 275.100 381.400 ;
        RECT 275.300 380.600 276.100 381.400 ;
        RECT 276.300 380.600 277.100 381.400 ;
        RECT 277.300 380.600 278.100 381.400 ;
        RECT 273.300 340.600 274.100 341.400 ;
        RECT 274.300 340.600 275.100 341.400 ;
        RECT 275.300 340.600 276.100 341.400 ;
        RECT 276.300 340.600 277.100 341.400 ;
        RECT 277.300 340.600 278.100 341.400 ;
        RECT 273.300 300.600 274.100 301.400 ;
        RECT 274.300 300.600 275.100 301.400 ;
        RECT 275.300 300.600 276.100 301.400 ;
        RECT 276.300 300.600 277.100 301.400 ;
        RECT 277.300 300.600 278.100 301.400 ;
        RECT 273.300 260.600 274.100 261.400 ;
        RECT 274.300 260.600 275.100 261.400 ;
        RECT 275.300 260.600 276.100 261.400 ;
        RECT 276.300 260.600 277.100 261.400 ;
        RECT 277.300 260.600 278.100 261.400 ;
        RECT 273.300 220.600 274.100 221.400 ;
        RECT 274.300 220.600 275.100 221.400 ;
        RECT 275.300 220.600 276.100 221.400 ;
        RECT 276.300 220.600 277.100 221.400 ;
        RECT 277.300 220.600 278.100 221.400 ;
        RECT 273.300 180.600 274.100 181.400 ;
        RECT 274.300 180.600 275.100 181.400 ;
        RECT 275.300 180.600 276.100 181.400 ;
        RECT 276.300 180.600 277.100 181.400 ;
        RECT 277.300 180.600 278.100 181.400 ;
        RECT 273.300 140.600 274.100 141.400 ;
        RECT 274.300 140.600 275.100 141.400 ;
        RECT 275.300 140.600 276.100 141.400 ;
        RECT 276.300 140.600 277.100 141.400 ;
        RECT 277.300 140.600 278.100 141.400 ;
        RECT 273.300 100.600 274.100 101.400 ;
        RECT 274.300 100.600 275.100 101.400 ;
        RECT 275.300 100.600 276.100 101.400 ;
        RECT 276.300 100.600 277.100 101.400 ;
        RECT 277.300 100.600 278.100 101.400 ;
        RECT 273.300 60.600 274.100 61.400 ;
        RECT 274.300 60.600 275.100 61.400 ;
        RECT 275.300 60.600 276.100 61.400 ;
        RECT 276.300 60.600 277.100 61.400 ;
        RECT 277.300 60.600 278.100 61.400 ;
        RECT 273.300 20.600 274.100 21.400 ;
        RECT 274.300 20.600 275.100 21.400 ;
        RECT 275.300 20.600 276.100 21.400 ;
        RECT 276.300 20.600 277.100 21.400 ;
        RECT 277.300 20.600 278.100 21.400 ;
      LAYER metal3 ;
        RECT 272.200 380.400 278.200 381.600 ;
        RECT 272.200 340.400 278.200 341.600 ;
        RECT 272.200 300.400 278.200 301.600 ;
        RECT 272.200 260.400 278.200 261.600 ;
        RECT 272.200 220.400 278.200 221.600 ;
        RECT 272.200 180.400 278.200 181.600 ;
        RECT 272.200 140.400 278.200 141.600 ;
        RECT 272.200 100.400 278.200 101.600 ;
        RECT 272.200 60.400 278.200 61.600 ;
        RECT 272.200 20.400 278.200 21.600 ;
      LAYER via3 ;
        RECT 272.400 380.600 273.200 381.400 ;
        RECT 273.600 380.600 274.400 381.400 ;
        RECT 274.800 380.600 275.600 381.400 ;
        RECT 276.000 380.600 276.800 381.400 ;
        RECT 277.200 380.600 278.000 381.400 ;
        RECT 272.400 340.600 273.200 341.400 ;
        RECT 273.600 340.600 274.400 341.400 ;
        RECT 274.800 340.600 275.600 341.400 ;
        RECT 276.000 340.600 276.800 341.400 ;
        RECT 277.200 340.600 278.000 341.400 ;
        RECT 272.400 300.600 273.200 301.400 ;
        RECT 273.600 300.600 274.400 301.400 ;
        RECT 274.800 300.600 275.600 301.400 ;
        RECT 276.000 300.600 276.800 301.400 ;
        RECT 277.200 300.600 278.000 301.400 ;
        RECT 272.400 260.600 273.200 261.400 ;
        RECT 273.600 260.600 274.400 261.400 ;
        RECT 274.800 260.600 275.600 261.400 ;
        RECT 276.000 260.600 276.800 261.400 ;
        RECT 277.200 260.600 278.000 261.400 ;
        RECT 272.400 220.600 273.200 221.400 ;
        RECT 273.600 220.600 274.400 221.400 ;
        RECT 274.800 220.600 275.600 221.400 ;
        RECT 276.000 220.600 276.800 221.400 ;
        RECT 277.200 220.600 278.000 221.400 ;
        RECT 272.400 180.600 273.200 181.400 ;
        RECT 273.600 180.600 274.400 181.400 ;
        RECT 274.800 180.600 275.600 181.400 ;
        RECT 276.000 180.600 276.800 181.400 ;
        RECT 277.200 180.600 278.000 181.400 ;
        RECT 272.400 140.600 273.200 141.400 ;
        RECT 273.600 140.600 274.400 141.400 ;
        RECT 274.800 140.600 275.600 141.400 ;
        RECT 276.000 140.600 276.800 141.400 ;
        RECT 277.200 140.600 278.000 141.400 ;
        RECT 272.400 100.600 273.200 101.400 ;
        RECT 273.600 100.600 274.400 101.400 ;
        RECT 274.800 100.600 275.600 101.400 ;
        RECT 276.000 100.600 276.800 101.400 ;
        RECT 277.200 100.600 278.000 101.400 ;
        RECT 272.400 60.600 273.200 61.400 ;
        RECT 273.600 60.600 274.400 61.400 ;
        RECT 274.800 60.600 275.600 61.400 ;
        RECT 276.000 60.600 276.800 61.400 ;
        RECT 277.200 60.600 278.000 61.400 ;
        RECT 272.400 20.600 273.200 21.400 ;
        RECT 273.600 20.600 274.400 21.400 ;
        RECT 274.800 20.600 275.600 21.400 ;
        RECT 276.000 20.600 276.800 21.400 ;
        RECT 277.200 20.600 278.000 21.400 ;
      LAYER metal4 ;
        RECT 272.000 -1.000 278.400 381.600 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 349.800 372.000 350.600 372.200 ;
        RECT 354.800 372.000 355.600 372.400 ;
        RECT 372.400 372.000 373.200 372.600 ;
        RECT 349.800 371.400 373.200 372.000 ;
        RECT 5.400 370.800 6.200 371.000 ;
        RECT 65.800 370.800 66.600 371.000 ;
        RECT 5.400 370.200 32.400 370.800 ;
        RECT 28.200 370.000 29.000 370.200 ;
        RECT 31.600 369.600 32.400 370.200 ;
        RECT 39.600 370.200 66.600 370.800 ;
        RECT 75.800 370.800 76.600 371.000 ;
        RECT 117.400 370.800 118.200 371.000 ;
        RECT 177.800 370.800 178.600 371.000 ;
        RECT 213.000 370.800 213.800 371.000 ;
        RECT 75.800 370.200 102.800 370.800 ;
        RECT 117.400 370.200 144.400 370.800 ;
        RECT 39.600 369.600 40.400 370.200 ;
        RECT 42.800 370.000 43.800 370.200 ;
        RECT 98.600 370.000 99.600 370.200 ;
        RECT 102.000 369.600 102.800 370.200 ;
        RECT 140.200 370.000 141.000 370.200 ;
        RECT 143.600 369.600 144.400 370.200 ;
        RECT 151.600 370.200 178.600 370.800 ;
        RECT 186.800 370.200 213.800 370.800 ;
        RECT 256.600 370.800 257.400 371.000 ;
        RECT 424.200 370.800 425.000 371.000 ;
        RECT 256.600 370.200 283.600 370.800 ;
        RECT 398.000 370.200 425.000 370.800 ;
        RECT 440.600 370.800 441.400 371.000 ;
        RECT 501.000 370.800 501.800 371.000 ;
        RECT 440.600 370.200 467.600 370.800 ;
        RECT 151.600 369.600 152.400 370.200 ;
        RECT 154.800 370.000 155.800 370.200 ;
        RECT 186.800 369.600 187.600 370.200 ;
        RECT 190.000 370.000 191.000 370.200 ;
        RECT 1.200 361.600 2.000 366.200 ;
        RECT 4.400 361.600 5.200 366.200 ;
        RECT 7.600 361.600 8.400 366.200 ;
        RECT 10.800 361.600 11.600 366.200 ;
        RECT 18.800 361.600 19.600 366.200 ;
        RECT 22.000 361.600 22.800 366.200 ;
        RECT 28.400 361.600 29.200 366.200 ;
        RECT 31.600 361.600 32.400 366.200 ;
        RECT 34.800 361.600 35.600 366.200 ;
        RECT 36.400 361.600 37.200 366.200 ;
        RECT 39.600 361.600 40.400 366.200 ;
        RECT 42.800 361.600 43.600 366.200 ;
        RECT 49.200 361.600 50.000 366.200 ;
        RECT 52.400 361.600 53.200 366.200 ;
        RECT 60.400 361.600 61.200 366.200 ;
        RECT 63.600 361.600 64.400 366.200 ;
        RECT 66.800 361.600 67.600 366.200 ;
        RECT 70.000 361.600 70.800 366.200 ;
        RECT 71.600 361.600 72.400 366.200 ;
        RECT 74.800 361.600 75.600 366.200 ;
        RECT 78.000 361.600 78.800 366.200 ;
        RECT 81.200 361.600 82.000 366.200 ;
        RECT 89.200 361.600 90.000 366.200 ;
        RECT 92.400 361.600 93.200 366.200 ;
        RECT 98.800 361.600 99.600 366.200 ;
        RECT 102.000 361.600 102.800 366.200 ;
        RECT 105.200 361.600 106.000 366.200 ;
        RECT 113.200 361.600 114.000 366.200 ;
        RECT 116.400 361.600 117.200 366.200 ;
        RECT 119.600 361.600 120.400 366.200 ;
        RECT 122.800 361.600 123.600 366.200 ;
        RECT 130.800 361.600 131.600 366.200 ;
        RECT 134.000 361.600 134.800 366.200 ;
        RECT 140.400 361.600 141.200 366.200 ;
        RECT 143.600 361.600 144.400 366.200 ;
        RECT 146.800 361.600 147.600 366.200 ;
        RECT 148.400 361.600 149.200 366.200 ;
        RECT 151.600 361.600 152.400 366.200 ;
        RECT 154.800 361.600 155.600 366.200 ;
        RECT 161.200 361.600 162.000 366.200 ;
        RECT 164.400 361.600 165.200 366.200 ;
        RECT 172.400 361.600 173.200 366.200 ;
        RECT 175.600 361.600 176.400 366.200 ;
        RECT 178.800 361.600 179.600 366.200 ;
        RECT 182.000 361.600 182.800 366.200 ;
        RECT 183.600 361.600 184.400 366.200 ;
        RECT 186.800 361.600 187.600 366.200 ;
        RECT 190.000 361.600 190.800 366.200 ;
        RECT 196.400 361.600 197.200 366.200 ;
        RECT 199.600 361.600 200.400 366.200 ;
        RECT 207.600 361.600 208.400 366.200 ;
        RECT 210.800 361.600 211.600 366.200 ;
        RECT 214.000 361.600 214.800 366.200 ;
        RECT 217.200 361.600 218.000 366.200 ;
        RECT 218.800 361.600 219.600 366.200 ;
        RECT 222.000 361.600 222.800 366.200 ;
        RECT 224.200 361.600 225.000 366.200 ;
        RECT 228.400 361.600 229.200 370.200 ;
        RECT 230.600 361.600 231.400 366.200 ;
        RECT 234.800 361.600 235.600 370.200 ;
        RECT 236.400 361.600 237.200 366.200 ;
        RECT 239.600 361.600 240.400 366.200 ;
        RECT 241.800 361.600 242.600 366.200 ;
        RECT 246.000 361.600 246.800 370.200 ;
        RECT 279.400 370.000 280.200 370.200 ;
        RECT 282.800 369.600 283.600 370.200 ;
        RECT 247.600 361.600 248.400 366.200 ;
        RECT 250.800 361.600 251.600 366.200 ;
        RECT 252.400 361.600 253.200 366.200 ;
        RECT 255.600 361.600 256.400 366.200 ;
        RECT 258.800 361.600 259.600 366.200 ;
        RECT 262.000 361.600 262.800 366.200 ;
        RECT 270.000 361.600 270.800 366.200 ;
        RECT 273.200 361.600 274.000 366.200 ;
        RECT 279.600 361.600 280.400 366.200 ;
        RECT 282.800 361.600 283.600 366.200 ;
        RECT 286.000 361.600 286.800 366.200 ;
        RECT 294.600 361.600 295.400 366.200 ;
        RECT 298.800 361.600 299.600 370.200 ;
        RECT 300.400 361.600 301.200 366.200 ;
        RECT 303.600 361.600 304.400 366.200 ;
        RECT 306.800 361.600 307.600 370.200 ;
        RECT 308.400 361.600 309.200 366.200 ;
        RECT 311.600 361.600 312.400 365.800 ;
        RECT 314.800 361.600 315.600 370.200 ;
        RECT 319.600 361.600 320.400 370.200 ;
        RECT 323.800 361.600 324.600 366.200 ;
        RECT 326.000 361.600 326.800 366.200 ;
        RECT 329.200 361.600 330.000 365.800 ;
        RECT 332.400 361.600 333.200 366.200 ;
        RECT 335.600 361.600 336.400 366.200 ;
        RECT 337.200 361.600 338.000 366.200 ;
        RECT 340.400 361.600 341.200 366.200 ;
        RECT 343.600 361.600 344.400 369.800 ;
        RECT 346.800 361.600 347.600 366.200 ;
        RECT 348.400 361.600 349.200 366.200 ;
        RECT 351.600 361.600 352.400 366.200 ;
        RECT 354.800 361.600 355.600 366.200 ;
        RECT 361.200 361.600 362.000 366.200 ;
        RECT 364.400 361.600 365.200 366.200 ;
        RECT 372.400 361.600 373.200 366.200 ;
        RECT 375.600 361.600 376.400 366.200 ;
        RECT 378.800 361.600 379.600 366.200 ;
        RECT 382.000 361.600 382.800 366.200 ;
        RECT 383.600 361.600 384.400 370.200 ;
        RECT 389.000 361.600 389.800 366.200 ;
        RECT 393.200 361.600 394.000 370.200 ;
        RECT 398.000 369.600 398.800 370.200 ;
        RECT 401.400 370.000 402.200 370.200 ;
        RECT 463.400 370.000 464.200 370.200 ;
        RECT 466.800 369.600 467.600 370.200 ;
        RECT 474.800 370.200 501.800 370.800 ;
        RECT 515.800 370.800 516.600 371.000 ;
        RECT 515.800 370.200 542.800 370.800 ;
        RECT 474.800 369.600 475.600 370.200 ;
        RECT 478.000 370.000 479.000 370.200 ;
        RECT 538.600 370.000 539.600 370.200 ;
        RECT 542.000 369.600 542.800 370.200 ;
        RECT 394.800 361.600 395.600 366.200 ;
        RECT 398.000 361.600 398.800 366.200 ;
        RECT 401.200 361.600 402.000 366.200 ;
        RECT 407.600 361.600 408.400 366.200 ;
        RECT 410.800 361.600 411.600 366.200 ;
        RECT 418.800 361.600 419.600 366.200 ;
        RECT 422.000 361.600 422.800 366.200 ;
        RECT 425.200 361.600 426.000 366.200 ;
        RECT 428.400 361.600 429.200 366.200 ;
        RECT 436.400 361.600 437.200 366.200 ;
        RECT 439.600 361.600 440.400 366.200 ;
        RECT 442.800 361.600 443.600 366.200 ;
        RECT 446.000 361.600 446.800 366.200 ;
        RECT 454.000 361.600 454.800 366.200 ;
        RECT 457.200 361.600 458.000 366.200 ;
        RECT 463.600 361.600 464.400 366.200 ;
        RECT 466.800 361.600 467.600 366.200 ;
        RECT 470.000 361.600 470.800 366.200 ;
        RECT 471.600 361.600 472.400 366.200 ;
        RECT 474.800 361.600 475.600 366.200 ;
        RECT 478.000 361.600 478.800 366.200 ;
        RECT 484.400 361.600 485.200 366.200 ;
        RECT 487.600 361.600 488.400 366.200 ;
        RECT 495.600 361.600 496.400 366.200 ;
        RECT 498.800 361.600 499.600 366.200 ;
        RECT 502.000 361.600 502.800 366.200 ;
        RECT 505.200 361.600 506.000 366.200 ;
        RECT 506.800 361.600 507.600 366.200 ;
        RECT 510.000 361.600 510.800 366.200 ;
        RECT 511.600 361.600 512.400 366.200 ;
        RECT 514.800 361.600 515.600 366.200 ;
        RECT 518.000 361.600 518.800 366.200 ;
        RECT 521.200 361.600 522.000 366.200 ;
        RECT 529.200 361.600 530.000 366.200 ;
        RECT 532.400 361.600 533.200 366.200 ;
        RECT 538.800 361.600 539.600 366.200 ;
        RECT 542.000 361.600 542.800 366.200 ;
        RECT 545.200 361.600 546.000 366.200 ;
        RECT 548.400 361.600 549.200 366.200 ;
        RECT 0.400 360.400 551.600 361.600 ;
        RECT 1.200 355.800 2.000 360.400 ;
        RECT 4.400 355.800 5.200 360.400 ;
        RECT 7.600 355.800 8.400 360.400 ;
        RECT 10.800 355.800 11.600 360.400 ;
        RECT 18.800 355.800 19.600 360.400 ;
        RECT 22.000 355.800 22.800 360.400 ;
        RECT 28.400 355.800 29.200 360.400 ;
        RECT 31.600 355.800 32.400 360.400 ;
        RECT 34.800 355.800 35.600 360.400 ;
        RECT 38.000 355.800 38.800 360.400 ;
        RECT 28.200 351.800 29.000 352.000 ;
        RECT 31.600 351.800 32.400 352.400 ;
        RECT 42.800 351.800 43.600 360.400 ;
        RECT 47.600 351.800 48.400 360.400 ;
        RECT 49.200 351.800 50.000 360.400 ;
        RECT 54.000 355.800 54.800 360.400 ;
        RECT 57.200 355.800 58.000 360.400 ;
        RECT 58.800 355.800 59.600 360.400 ;
        RECT 62.000 355.800 62.800 360.400 ;
        RECT 65.200 355.800 66.000 360.400 ;
        RECT 71.600 355.800 72.400 360.400 ;
        RECT 74.800 355.800 75.600 360.400 ;
        RECT 82.800 355.800 83.600 360.400 ;
        RECT 86.000 355.800 86.800 360.400 ;
        RECT 89.200 355.800 90.000 360.400 ;
        RECT 92.400 355.800 93.200 360.400 ;
        RECT 62.000 351.800 62.800 352.400 ;
        RECT 65.200 351.800 66.200 352.000 ;
        RECT 97.200 351.800 98.000 360.400 ;
        RECT 98.800 355.800 99.600 360.400 ;
        RECT 102.000 355.800 102.800 360.400 ;
        RECT 105.200 355.800 106.000 360.400 ;
        RECT 111.600 355.800 112.400 360.400 ;
        RECT 114.800 355.800 115.600 360.400 ;
        RECT 122.800 355.800 123.600 360.400 ;
        RECT 126.000 355.800 126.800 360.400 ;
        RECT 129.200 355.800 130.000 360.400 ;
        RECT 132.400 355.800 133.200 360.400 ;
        RECT 140.400 355.800 141.200 360.400 ;
        RECT 143.600 355.800 144.400 360.400 ;
        RECT 146.800 355.800 147.600 360.400 ;
        RECT 153.200 355.800 154.000 360.400 ;
        RECT 156.400 355.800 157.200 360.400 ;
        RECT 164.400 355.800 165.200 360.400 ;
        RECT 167.600 355.800 168.400 360.400 ;
        RECT 170.800 355.800 171.600 360.400 ;
        RECT 174.000 355.800 174.800 360.400 ;
        RECT 175.600 355.800 176.400 360.400 ;
        RECT 178.800 355.800 179.600 360.400 ;
        RECT 182.000 355.800 182.800 360.400 ;
        RECT 185.200 355.800 186.000 360.400 ;
        RECT 193.200 355.800 194.000 360.400 ;
        RECT 196.400 355.800 197.200 360.400 ;
        RECT 202.800 355.800 203.600 360.400 ;
        RECT 206.000 355.800 206.800 360.400 ;
        RECT 209.200 355.800 210.000 360.400 ;
        RECT 210.800 355.800 211.600 360.400 ;
        RECT 214.000 355.800 214.800 360.400 ;
        RECT 217.200 355.800 218.000 360.400 ;
        RECT 220.400 355.800 221.200 360.400 ;
        RECT 228.400 355.800 229.200 360.400 ;
        RECT 231.600 355.800 232.400 360.400 ;
        RECT 238.000 355.800 238.800 360.400 ;
        RECT 241.200 355.800 242.000 360.400 ;
        RECT 244.400 355.800 245.200 360.400 ;
        RECT 247.600 356.200 248.400 360.400 ;
        RECT 250.800 355.800 251.600 360.400 ;
        RECT 254.000 356.200 254.800 360.400 ;
        RECT 257.200 355.800 258.000 360.400 ;
        RECT 265.200 355.800 266.000 360.400 ;
        RECT 268.400 355.800 269.200 360.400 ;
        RECT 271.600 355.800 272.400 360.400 ;
        RECT 278.000 355.800 278.800 360.400 ;
        RECT 281.200 355.800 282.000 360.400 ;
        RECT 289.200 355.800 290.000 360.400 ;
        RECT 292.400 355.800 293.200 360.400 ;
        RECT 295.600 355.800 296.400 360.400 ;
        RECT 298.800 355.800 299.600 360.400 ;
        RECT 302.000 356.200 302.800 360.400 ;
        RECT 305.200 355.800 306.000 360.400 ;
        RECT 102.000 351.800 102.800 352.400 ;
        RECT 105.200 351.800 106.200 352.000 ;
        RECT 143.600 351.800 144.400 352.400 ;
        RECT 147.000 351.800 147.800 352.000 ;
        RECT 202.600 351.800 203.600 352.000 ;
        RECT 206.000 351.800 206.800 352.400 ;
        RECT 237.800 351.800 238.800 352.000 ;
        RECT 241.200 351.800 242.000 352.400 ;
        RECT 5.400 351.200 32.400 351.800 ;
        RECT 62.000 351.200 89.000 351.800 ;
        RECT 102.000 351.200 129.000 351.800 ;
        RECT 143.600 351.200 170.600 351.800 ;
        RECT 5.400 351.000 6.200 351.200 ;
        RECT 88.200 351.000 89.000 351.200 ;
        RECT 128.200 351.000 129.000 351.200 ;
        RECT 169.800 351.000 170.600 351.200 ;
        RECT 179.800 351.200 206.800 351.800 ;
        RECT 215.000 351.200 242.000 351.800 ;
        RECT 268.400 351.800 269.200 352.400 ;
        RECT 271.800 351.800 272.600 352.000 ;
        RECT 310.000 351.800 310.800 360.400 ;
        RECT 313.200 352.200 314.000 360.400 ;
        RECT 316.400 355.800 317.200 360.400 ;
        RECT 318.000 355.800 318.800 360.400 ;
        RECT 321.200 355.800 322.000 360.400 ;
        RECT 324.400 356.200 325.200 360.400 ;
        RECT 327.600 355.800 328.400 360.400 ;
        RECT 332.400 353.000 333.200 360.400 ;
        RECT 337.200 356.200 338.000 360.400 ;
        RECT 340.400 355.800 341.200 360.400 ;
        RECT 345.200 351.800 346.000 360.400 ;
        RECT 350.000 351.800 350.800 360.400 ;
        RECT 351.600 351.800 352.400 360.400 ;
        RECT 355.800 355.800 356.600 360.400 ;
        RECT 358.600 355.800 359.400 360.400 ;
        RECT 362.800 351.800 363.600 360.400 ;
        RECT 364.400 351.800 365.200 360.400 ;
        RECT 370.800 351.800 371.600 360.400 ;
        RECT 373.000 355.800 373.800 360.400 ;
        RECT 377.200 351.800 378.000 360.400 ;
        RECT 382.000 353.000 382.800 360.400 ;
        RECT 386.800 351.800 387.600 360.400 ;
        RECT 391.600 353.000 392.400 360.400 ;
        RECT 396.400 353.000 397.200 360.400 ;
        RECT 402.800 353.000 403.600 360.400 ;
        RECT 409.200 353.800 410.000 360.400 ;
        RECT 423.600 351.800 424.400 360.400 ;
        RECT 431.600 355.800 432.400 360.400 ;
        RECT 434.800 355.800 435.600 360.400 ;
        RECT 436.400 355.800 437.200 360.400 ;
        RECT 439.600 355.800 440.400 360.400 ;
        RECT 441.200 355.800 442.000 360.400 ;
        RECT 444.400 356.200 445.200 360.400 ;
        RECT 447.600 351.800 448.400 360.400 ;
        RECT 451.800 355.800 452.600 360.400 ;
        RECT 454.000 351.800 454.800 360.400 ;
        RECT 460.400 351.800 461.200 360.400 ;
        RECT 462.600 355.800 463.400 360.400 ;
        RECT 466.800 351.800 467.600 360.400 ;
        RECT 470.000 355.800 470.800 360.400 ;
        RECT 471.600 351.800 472.400 360.400 ;
        RECT 475.800 355.800 476.600 360.400 ;
        RECT 478.000 351.800 478.800 360.400 ;
        RECT 482.200 355.800 483.000 360.400 ;
        RECT 484.400 355.800 485.200 360.400 ;
        RECT 487.600 355.800 488.400 360.400 ;
        RECT 490.800 355.800 491.600 360.400 ;
        RECT 494.000 356.200 494.800 360.400 ;
        RECT 497.200 355.800 498.000 360.400 ;
        RECT 500.400 356.200 501.200 360.400 ;
        RECT 506.800 351.800 507.600 360.400 ;
        RECT 511.600 353.000 512.400 360.400 ;
        RECT 514.800 355.800 515.600 360.400 ;
        RECT 518.000 355.800 518.800 360.400 ;
        RECT 521.200 355.800 522.000 360.400 ;
        RECT 524.400 355.800 525.200 360.400 ;
        RECT 532.400 355.800 533.200 360.400 ;
        RECT 535.600 355.800 536.400 360.400 ;
        RECT 542.000 355.800 542.800 360.400 ;
        RECT 545.200 355.800 546.000 360.400 ;
        RECT 548.400 355.800 549.200 360.400 ;
        RECT 541.800 351.800 542.600 352.000 ;
        RECT 545.200 351.800 546.000 352.400 ;
        RECT 268.400 351.200 295.400 351.800 ;
        RECT 179.800 351.000 180.600 351.200 ;
        RECT 215.000 351.000 215.800 351.200 ;
        RECT 294.600 351.000 295.400 351.200 ;
        RECT 519.000 351.200 546.000 351.800 ;
        RECT 519.000 351.000 519.800 351.200 ;
        RECT 8.600 330.800 9.400 331.000 ;
        RECT 98.200 330.800 99.000 331.000 ;
        RECT 165.000 330.800 165.800 331.000 ;
        RECT 8.600 330.200 35.600 330.800 ;
        RECT 98.200 330.200 125.200 330.800 ;
        RECT 31.400 330.000 32.200 330.200 ;
        RECT 34.800 329.600 35.600 330.200 ;
        RECT 1.200 321.600 2.000 326.200 ;
        RECT 4.400 321.600 5.200 326.200 ;
        RECT 7.600 321.600 8.400 326.200 ;
        RECT 10.800 321.600 11.600 326.200 ;
        RECT 14.000 321.600 14.800 326.200 ;
        RECT 22.000 321.600 22.800 326.200 ;
        RECT 25.200 321.600 26.000 326.200 ;
        RECT 31.600 321.600 32.400 326.200 ;
        RECT 34.800 321.600 35.600 326.200 ;
        RECT 38.000 321.600 38.800 326.200 ;
        RECT 39.600 321.600 40.400 326.200 ;
        RECT 42.800 321.600 43.600 326.200 ;
        RECT 45.000 321.600 45.800 326.200 ;
        RECT 49.200 321.600 50.000 330.200 ;
        RECT 50.800 321.600 51.600 326.200 ;
        RECT 54.000 321.600 54.800 325.800 ;
        RECT 57.200 321.600 58.000 326.200 ;
        RECT 60.400 321.600 61.200 325.800 ;
        RECT 64.200 321.600 65.000 326.200 ;
        RECT 68.400 321.600 69.200 330.200 ;
        RECT 70.000 321.600 70.800 326.200 ;
        RECT 73.200 321.600 74.000 326.200 ;
        RECT 74.800 321.600 75.600 326.200 ;
        RECT 78.000 321.600 78.800 326.200 ;
        RECT 79.600 321.600 80.400 330.200 ;
        RECT 121.000 330.000 122.000 330.200 ;
        RECT 124.400 329.600 125.200 330.200 ;
        RECT 138.800 330.200 165.800 330.800 ;
        RECT 223.000 330.800 223.800 331.000 ;
        RECT 304.200 330.800 305.000 331.000 ;
        RECT 339.400 330.800 340.200 331.000 ;
        RECT 488.200 330.800 489.000 331.000 ;
        RECT 223.000 330.200 250.000 330.800 ;
        RECT 278.000 330.200 305.000 330.800 ;
        RECT 313.200 330.200 340.200 330.800 ;
        RECT 462.000 330.200 489.000 330.800 ;
        RECT 138.800 329.600 139.600 330.200 ;
        RECT 142.000 330.000 143.000 330.200 ;
        RECT 86.000 321.600 86.800 325.800 ;
        RECT 89.200 321.600 90.000 326.200 ;
        RECT 92.400 321.600 93.200 326.200 ;
        RECT 94.000 321.600 94.800 326.200 ;
        RECT 97.200 321.600 98.000 326.200 ;
        RECT 100.400 321.600 101.200 326.200 ;
        RECT 103.600 321.600 104.400 326.200 ;
        RECT 111.600 321.600 112.400 326.200 ;
        RECT 114.800 321.600 115.600 326.200 ;
        RECT 121.200 321.600 122.000 326.200 ;
        RECT 124.400 321.600 125.200 326.200 ;
        RECT 127.600 321.600 128.400 326.200 ;
        RECT 135.600 321.600 136.400 326.200 ;
        RECT 138.800 321.600 139.600 326.200 ;
        RECT 142.000 321.600 142.800 326.200 ;
        RECT 148.400 321.600 149.200 326.200 ;
        RECT 151.600 321.600 152.400 326.200 ;
        RECT 159.600 321.600 160.400 326.200 ;
        RECT 162.800 321.600 163.600 326.200 ;
        RECT 166.000 321.600 166.800 326.200 ;
        RECT 169.200 321.600 170.000 326.200 ;
        RECT 172.400 321.600 173.200 329.000 ;
        RECT 176.200 321.600 177.000 326.200 ;
        RECT 180.400 321.600 181.200 330.200 ;
        RECT 182.000 321.600 182.800 326.200 ;
        RECT 185.200 321.600 186.000 326.200 ;
        RECT 188.400 321.600 189.200 325.800 ;
        RECT 191.600 321.600 192.400 326.200 ;
        RECT 194.800 321.600 195.600 330.200 ;
        RECT 199.000 321.600 199.800 326.200 ;
        RECT 201.200 321.600 202.000 326.200 ;
        RECT 204.400 321.600 205.200 326.200 ;
        RECT 207.600 321.600 208.400 329.000 ;
        RECT 212.400 321.600 213.200 326.200 ;
        RECT 214.000 321.600 214.800 330.200 ;
        RECT 245.800 330.000 246.800 330.200 ;
        RECT 249.200 329.600 250.000 330.200 ;
        RECT 218.800 321.600 219.600 326.200 ;
        RECT 222.000 321.600 222.800 326.200 ;
        RECT 225.200 321.600 226.000 326.200 ;
        RECT 228.400 321.600 229.200 326.200 ;
        RECT 236.400 321.600 237.200 326.200 ;
        RECT 239.600 321.600 240.400 326.200 ;
        RECT 246.000 321.600 246.800 326.200 ;
        RECT 249.200 321.600 250.000 326.200 ;
        RECT 252.400 321.600 253.200 326.200 ;
        RECT 254.000 321.600 254.800 330.200 ;
        RECT 257.200 321.600 258.000 330.200 ;
        RECT 260.400 321.600 261.200 330.200 ;
        RECT 263.600 321.600 264.400 330.200 ;
        RECT 266.800 321.600 267.600 330.200 ;
        RECT 278.000 329.600 278.800 330.200 ;
        RECT 281.400 330.000 282.200 330.200 ;
        RECT 313.200 329.600 314.000 330.200 ;
        RECT 316.400 330.000 317.400 330.200 ;
        RECT 274.800 321.600 275.600 326.200 ;
        RECT 278.000 321.600 278.800 326.200 ;
        RECT 281.200 321.600 282.000 326.200 ;
        RECT 287.600 321.600 288.400 326.200 ;
        RECT 290.800 321.600 291.600 326.200 ;
        RECT 298.800 321.600 299.600 326.200 ;
        RECT 302.000 321.600 302.800 326.200 ;
        RECT 305.200 321.600 306.000 326.200 ;
        RECT 308.400 321.600 309.200 326.200 ;
        RECT 310.000 321.600 310.800 326.200 ;
        RECT 313.200 321.600 314.000 326.200 ;
        RECT 316.400 321.600 317.200 326.200 ;
        RECT 322.800 321.600 323.600 326.200 ;
        RECT 326.000 321.600 326.800 326.200 ;
        RECT 334.000 321.600 334.800 326.200 ;
        RECT 337.200 321.600 338.000 326.200 ;
        RECT 340.400 321.600 341.200 326.200 ;
        RECT 343.600 321.600 344.400 326.200 ;
        RECT 345.200 321.600 346.000 330.200 ;
        RECT 348.400 321.600 349.200 326.200 ;
        RECT 351.600 321.600 352.400 326.200 ;
        RECT 354.800 321.600 355.600 329.000 ;
        RECT 360.200 321.600 361.000 326.200 ;
        RECT 364.400 321.600 365.200 330.200 ;
        RECT 366.600 321.600 367.400 326.200 ;
        RECT 370.800 321.600 371.600 330.200 ;
        RECT 374.000 321.600 374.800 326.200 ;
        RECT 375.600 321.600 376.400 326.200 ;
        RECT 378.800 321.600 379.600 326.200 ;
        RECT 380.400 321.600 381.200 326.200 ;
        RECT 383.600 321.600 384.400 326.200 ;
        RECT 385.200 321.600 386.000 330.200 ;
        RECT 389.000 321.600 389.800 326.200 ;
        RECT 393.200 321.600 394.000 330.200 ;
        RECT 394.800 321.600 395.600 326.200 ;
        RECT 398.000 321.600 398.800 326.200 ;
        RECT 399.600 321.600 400.400 326.200 ;
        RECT 402.800 321.600 403.600 326.200 ;
        RECT 405.000 321.600 405.800 326.200 ;
        RECT 409.200 321.600 410.000 330.200 ;
        RECT 414.000 321.600 414.800 330.200 ;
        RECT 417.200 321.600 418.000 326.200 ;
        RECT 426.800 321.600 427.600 328.200 ;
        RECT 438.000 321.600 438.800 326.200 ;
        RECT 441.200 321.600 442.000 325.800 ;
        RECT 445.000 321.600 445.800 326.200 ;
        RECT 449.200 321.600 450.000 330.200 ;
        RECT 452.400 321.600 453.200 330.200 ;
        RECT 457.200 321.600 458.000 330.200 ;
        RECT 462.000 329.600 462.800 330.200 ;
        RECT 465.400 330.000 466.200 330.200 ;
        RECT 458.800 321.600 459.600 326.200 ;
        RECT 462.000 321.600 462.800 326.200 ;
        RECT 465.200 321.600 466.000 326.200 ;
        RECT 471.600 321.600 472.400 326.200 ;
        RECT 474.800 321.600 475.600 326.200 ;
        RECT 482.800 321.600 483.600 326.200 ;
        RECT 486.000 321.600 486.800 326.200 ;
        RECT 489.200 321.600 490.000 326.200 ;
        RECT 492.400 321.600 493.200 326.200 ;
        RECT 494.000 321.600 494.800 326.200 ;
        RECT 497.200 321.600 498.000 326.200 ;
        RECT 499.400 321.600 500.200 326.200 ;
        RECT 503.600 321.600 504.400 330.200 ;
        RECT 506.800 321.600 507.600 326.200 ;
        RECT 508.400 321.600 509.200 330.200 ;
        RECT 512.600 321.600 513.400 326.200 ;
        RECT 514.800 321.600 515.600 330.200 ;
        RECT 519.000 321.600 519.800 326.200 ;
        RECT 524.400 321.600 525.200 330.200 ;
        RECT 526.000 321.600 526.800 326.200 ;
        RECT 529.200 321.600 530.000 330.200 ;
        RECT 533.400 321.600 534.200 326.200 ;
        RECT 535.600 321.600 536.400 330.200 ;
        RECT 539.800 321.600 540.600 326.200 ;
        RECT 543.600 321.600 544.400 326.200 ;
        RECT 546.800 321.600 547.600 329.000 ;
        RECT 0.400 320.400 551.600 321.600 ;
        RECT 4.400 311.800 5.200 320.400 ;
        RECT 6.000 315.800 6.800 320.400 ;
        RECT 9.200 316.200 10.000 320.400 ;
        RECT 14.000 315.800 14.800 320.400 ;
        RECT 17.200 316.200 18.000 320.400 ;
        RECT 20.400 315.800 21.200 320.400 ;
        RECT 22.000 315.800 22.800 320.400 ;
        RECT 25.200 315.800 26.000 320.400 ;
        RECT 27.400 315.800 28.200 320.400 ;
        RECT 31.600 311.800 32.400 320.400 ;
        RECT 33.200 311.800 34.000 320.400 ;
        RECT 38.000 311.800 38.800 320.400 ;
        RECT 42.800 311.800 43.600 320.400 ;
        RECT 49.200 311.800 50.000 320.400 ;
        RECT 50.800 315.800 51.600 320.400 ;
        RECT 54.000 315.800 54.800 320.400 ;
        RECT 55.600 315.800 56.400 320.400 ;
        RECT 58.800 316.200 59.600 320.400 ;
        RECT 62.000 315.800 62.800 320.400 ;
        RECT 65.200 315.800 66.000 320.400 ;
        RECT 66.800 311.800 67.600 320.400 ;
        RECT 73.200 311.800 74.000 320.400 ;
        RECT 74.800 315.800 75.600 320.400 ;
        RECT 78.000 311.800 78.800 320.400 ;
        RECT 81.200 311.800 82.000 320.400 ;
        RECT 84.400 311.800 85.200 320.400 ;
        RECT 87.600 311.800 88.400 320.400 ;
        RECT 90.800 311.800 91.600 320.400 ;
        RECT 92.400 311.800 93.200 320.400 ;
        RECT 96.600 315.800 97.400 320.400 ;
        RECT 98.800 315.800 99.600 320.400 ;
        RECT 102.000 315.800 102.800 320.400 ;
        RECT 103.600 311.800 104.400 320.400 ;
        RECT 106.800 311.800 107.600 320.400 ;
        RECT 108.400 315.800 109.200 320.400 ;
        RECT 111.600 315.800 112.400 320.400 ;
        RECT 114.800 311.800 115.600 320.400 ;
        RECT 119.600 315.800 120.400 320.400 ;
        RECT 122.800 312.200 123.600 320.400 ;
        RECT 134.000 316.200 134.800 320.400 ;
        RECT 137.200 315.800 138.000 320.400 ;
        RECT 138.800 311.800 139.600 320.400 ;
        RECT 143.000 315.800 143.800 320.400 ;
        RECT 145.200 311.800 146.000 320.400 ;
        RECT 148.400 311.800 149.200 320.400 ;
        RECT 151.600 311.800 152.400 320.400 ;
        RECT 154.800 311.800 155.600 320.400 ;
        RECT 158.000 311.800 158.800 320.400 ;
        RECT 161.200 313.000 162.000 320.400 ;
        RECT 166.600 315.800 167.400 320.400 ;
        RECT 170.800 311.800 171.600 320.400 ;
        RECT 173.000 315.800 173.800 320.400 ;
        RECT 177.200 311.800 178.000 320.400 ;
        RECT 178.800 315.800 179.600 320.400 ;
        RECT 182.000 315.800 182.800 320.400 ;
        RECT 185.200 315.800 186.000 320.400 ;
        RECT 186.800 311.800 187.600 320.400 ;
        RECT 192.200 315.800 193.000 320.400 ;
        RECT 196.400 311.800 197.200 320.400 ;
        RECT 199.600 315.800 200.400 320.400 ;
        RECT 201.200 315.800 202.000 320.400 ;
        RECT 204.400 315.800 205.200 320.400 ;
        RECT 206.600 315.800 207.400 320.400 ;
        RECT 210.800 311.800 211.600 320.400 ;
        RECT 212.400 311.800 213.200 320.400 ;
        RECT 216.600 315.800 217.400 320.400 ;
        RECT 218.800 315.800 219.600 320.400 ;
        RECT 222.000 315.800 222.800 320.400 ;
        RECT 223.600 315.800 224.400 320.400 ;
        RECT 226.800 315.800 227.600 320.400 ;
        RECT 228.400 315.800 229.200 320.400 ;
        RECT 231.600 315.800 232.400 320.400 ;
        RECT 233.800 315.800 234.600 320.400 ;
        RECT 238.000 311.800 238.800 320.400 ;
        RECT 239.600 315.800 240.400 320.400 ;
        RECT 242.800 311.800 243.600 320.400 ;
        RECT 247.000 315.800 247.800 320.400 ;
        RECT 249.200 315.800 250.000 320.400 ;
        RECT 252.400 315.800 253.200 320.400 ;
        RECT 255.600 315.800 256.400 320.400 ;
        RECT 258.800 315.800 259.600 320.400 ;
        RECT 266.800 315.800 267.600 320.400 ;
        RECT 270.000 315.800 270.800 320.400 ;
        RECT 276.400 315.800 277.200 320.400 ;
        RECT 279.600 315.800 280.400 320.400 ;
        RECT 282.800 315.800 283.600 320.400 ;
        RECT 290.800 315.800 291.600 320.400 ;
        RECT 294.000 315.800 294.800 320.400 ;
        RECT 297.200 315.800 298.000 320.400 ;
        RECT 300.400 315.800 301.200 320.400 ;
        RECT 308.400 315.800 309.200 320.400 ;
        RECT 311.600 315.600 312.400 320.400 ;
        RECT 318.000 315.800 318.800 320.400 ;
        RECT 321.200 315.800 322.000 320.400 ;
        RECT 324.400 315.800 325.200 320.400 ;
        RECT 327.600 313.000 328.400 320.400 ;
        RECT 333.000 315.800 333.800 320.400 ;
        RECT 276.200 311.800 277.000 312.000 ;
        RECT 279.600 311.800 280.400 312.400 ;
        RECT 337.200 311.800 338.000 320.400 ;
        RECT 340.400 315.800 341.200 320.400 ;
        RECT 343.600 313.000 344.400 320.400 ;
        RECT 346.800 311.800 347.600 320.400 ;
        RECT 351.000 315.800 351.800 320.400 ;
        RECT 353.200 315.800 354.000 320.400 ;
        RECT 356.400 315.800 357.200 320.400 ;
        RECT 358.000 315.800 358.800 320.400 ;
        RECT 361.200 316.200 362.000 320.400 ;
        RECT 364.400 315.800 365.200 320.400 ;
        RECT 372.400 313.000 373.200 320.400 ;
        RECT 375.600 315.800 376.400 320.400 ;
        RECT 378.800 315.800 379.600 320.400 ;
        RECT 382.000 313.000 382.800 320.400 ;
        RECT 390.000 315.800 390.800 320.400 ;
        RECT 392.200 315.800 393.000 320.400 ;
        RECT 396.400 311.800 397.200 320.400 ;
        RECT 398.000 315.800 398.800 320.400 ;
        RECT 401.200 316.200 402.000 320.400 ;
        RECT 406.000 316.200 406.800 320.400 ;
        RECT 409.200 315.800 410.000 320.400 ;
        RECT 412.400 315.800 413.200 320.400 ;
        RECT 417.200 311.800 418.000 320.400 ;
        RECT 426.800 313.800 427.600 320.400 ;
        RECT 439.600 315.800 440.400 320.400 ;
        RECT 441.200 315.800 442.000 320.400 ;
        RECT 444.400 315.800 445.200 320.400 ;
        RECT 447.600 315.800 448.400 320.400 ;
        RECT 454.000 315.800 454.800 320.400 ;
        RECT 457.200 315.800 458.000 320.400 ;
        RECT 465.200 315.800 466.000 320.400 ;
        RECT 468.400 315.800 469.200 320.400 ;
        RECT 471.600 315.800 472.400 320.400 ;
        RECT 474.800 315.800 475.600 320.400 ;
        RECT 476.400 315.800 477.200 320.400 ;
        RECT 444.400 311.800 445.200 312.400 ;
        RECT 447.800 311.800 448.600 312.000 ;
        RECT 479.600 311.800 480.400 320.400 ;
        RECT 482.800 311.800 483.600 320.400 ;
        RECT 486.000 311.800 486.800 320.400 ;
        RECT 489.200 311.800 490.000 320.400 ;
        RECT 492.400 311.800 493.200 320.400 ;
        RECT 494.000 315.800 494.800 320.400 ;
        RECT 506.800 313.800 507.600 320.400 ;
        RECT 510.000 311.800 510.800 320.400 ;
        RECT 514.200 315.800 515.000 320.400 ;
        RECT 516.400 315.800 517.200 320.400 ;
        RECT 521.200 313.000 522.000 320.400 ;
        RECT 526.000 315.800 526.800 320.400 ;
        RECT 529.200 311.800 530.000 320.400 ;
        RECT 533.400 315.800 534.200 320.400 ;
        RECT 535.600 311.800 536.400 320.400 ;
        RECT 539.800 315.800 540.600 320.400 ;
        RECT 542.000 315.800 542.800 320.400 ;
        RECT 545.200 315.800 546.000 320.400 ;
        RECT 253.400 311.200 280.400 311.800 ;
        RECT 444.400 311.200 471.400 311.800 ;
        RECT 253.400 311.000 254.200 311.200 ;
        RECT 470.600 311.000 471.400 311.200 ;
        RECT 300.400 310.000 323.800 310.600 ;
        RECT 300.400 309.400 301.200 310.000 ;
        RECT 311.600 309.600 312.400 310.000 ;
        RECT 318.000 309.600 318.800 310.000 ;
        RECT 323.000 309.800 323.800 310.000 ;
        RECT 42.200 290.800 43.000 291.000 ;
        RECT 77.400 290.800 78.200 291.000 ;
        RECT 279.000 290.800 279.800 291.000 ;
        RECT 455.000 290.800 455.800 291.000 ;
        RECT 517.400 290.800 518.200 291.000 ;
        RECT 42.200 290.200 69.200 290.800 ;
        RECT 77.400 290.200 104.400 290.800 ;
        RECT 279.000 290.200 306.000 290.800 ;
        RECT 455.000 290.200 482.000 290.800 ;
        RECT 517.400 290.200 544.400 290.800 ;
        RECT 2.800 281.600 3.600 285.800 ;
        RECT 6.000 281.600 6.800 286.200 ;
        RECT 9.200 281.600 10.000 286.200 ;
        RECT 10.800 281.600 11.600 290.200 ;
        RECT 15.600 281.600 16.400 286.200 ;
        RECT 18.800 281.600 19.600 286.200 ;
        RECT 22.000 281.600 22.800 286.200 ;
        RECT 25.200 281.600 26.000 285.800 ;
        RECT 28.400 281.600 29.200 286.200 ;
        RECT 31.600 281.600 32.400 286.200 ;
        RECT 33.200 281.600 34.000 290.200 ;
        RECT 65.000 290.000 66.000 290.200 ;
        RECT 68.400 289.600 69.200 290.200 ;
        RECT 100.200 290.000 101.200 290.200 ;
        RECT 103.600 289.600 104.400 290.200 ;
        RECT 38.000 281.600 38.800 286.200 ;
        RECT 41.200 281.600 42.000 286.200 ;
        RECT 44.400 281.600 45.200 286.200 ;
        RECT 47.600 281.600 48.400 286.200 ;
        RECT 55.600 281.600 56.400 286.200 ;
        RECT 58.800 281.600 59.600 286.200 ;
        RECT 65.200 281.600 66.000 286.200 ;
        RECT 68.400 281.600 69.200 286.200 ;
        RECT 71.600 281.600 72.400 286.200 ;
        RECT 73.200 281.600 74.000 286.200 ;
        RECT 76.400 281.600 77.200 286.200 ;
        RECT 79.600 281.600 80.400 286.200 ;
        RECT 82.800 281.600 83.600 286.200 ;
        RECT 90.800 281.600 91.600 286.200 ;
        RECT 94.000 281.600 94.800 286.200 ;
        RECT 100.400 281.600 101.200 286.200 ;
        RECT 103.600 281.600 104.400 286.200 ;
        RECT 106.800 281.600 107.600 286.200 ;
        RECT 108.400 281.600 109.200 286.200 ;
        RECT 111.600 281.600 112.400 286.200 ;
        RECT 113.800 281.600 114.600 286.200 ;
        RECT 118.000 281.600 118.800 290.200 ;
        RECT 119.600 281.600 120.400 290.200 ;
        RECT 130.800 281.600 131.600 290.200 ;
        RECT 135.000 281.600 135.800 286.200 ;
        RECT 137.200 281.600 138.000 286.200 ;
        RECT 140.400 281.600 141.200 290.200 ;
        RECT 144.600 281.600 145.400 286.200 ;
        RECT 148.400 281.600 149.200 285.800 ;
        RECT 151.600 281.600 152.400 286.200 ;
        RECT 156.400 281.600 157.200 290.200 ;
        RECT 158.000 281.600 158.800 290.200 ;
        RECT 162.200 281.600 163.000 286.200 ;
        RECT 164.400 281.600 165.200 286.200 ;
        RECT 167.600 281.600 168.400 286.200 ;
        RECT 169.200 281.600 170.000 290.200 ;
        RECT 175.600 281.600 176.400 289.000 ;
        RECT 182.000 281.600 182.800 286.200 ;
        RECT 185.200 281.600 186.000 286.200 ;
        RECT 187.400 281.600 188.200 286.200 ;
        RECT 191.600 281.600 192.400 290.200 ;
        RECT 195.400 281.600 196.200 290.200 ;
        RECT 204.400 281.600 205.200 289.000 ;
        RECT 209.800 281.600 210.600 290.200 ;
        RECT 214.000 281.600 214.800 286.200 ;
        RECT 217.200 281.600 218.000 286.200 ;
        RECT 223.600 281.600 224.400 289.000 ;
        RECT 231.600 281.600 232.400 289.000 ;
        RECT 239.600 281.600 240.400 289.000 ;
        RECT 242.800 281.600 243.600 286.200 ;
        RECT 246.000 281.600 246.800 289.800 ;
        RECT 249.200 281.600 250.000 286.200 ;
        RECT 254.000 281.600 254.800 289.000 ;
        RECT 258.800 281.600 259.600 286.200 ;
        RECT 262.000 281.600 262.800 290.200 ;
        RECT 301.800 290.000 302.800 290.200 ;
        RECT 305.200 289.600 306.000 290.200 ;
        RECT 266.200 281.600 267.000 286.200 ;
        RECT 274.800 281.600 275.600 286.200 ;
        RECT 278.000 281.600 278.800 286.200 ;
        RECT 281.200 281.600 282.000 286.200 ;
        RECT 284.400 281.600 285.200 286.200 ;
        RECT 292.400 281.600 293.200 286.200 ;
        RECT 295.600 281.600 296.400 286.200 ;
        RECT 302.000 281.600 302.800 286.200 ;
        RECT 305.200 281.600 306.000 286.200 ;
        RECT 308.400 281.600 309.200 286.200 ;
        RECT 310.000 281.600 310.800 290.200 ;
        RECT 313.200 281.600 314.000 290.200 ;
        RECT 316.400 281.600 317.200 290.200 ;
        RECT 319.600 281.600 320.400 290.200 ;
        RECT 322.800 281.600 323.600 290.200 ;
        RECT 326.000 281.600 326.800 285.800 ;
        RECT 329.200 281.600 330.000 286.200 ;
        RECT 330.800 281.600 331.600 286.200 ;
        RECT 334.000 281.600 334.800 290.200 ;
        RECT 338.200 281.600 339.000 286.200 ;
        RECT 341.000 281.600 341.800 286.200 ;
        RECT 345.200 281.600 346.000 290.200 ;
        RECT 350.000 281.600 350.800 290.200 ;
        RECT 353.200 281.600 354.000 288.200 ;
        RECT 367.600 281.600 368.400 289.000 ;
        RECT 372.400 281.600 373.200 290.200 ;
        RECT 375.600 281.600 376.400 286.200 ;
        RECT 377.800 281.600 378.600 286.200 ;
        RECT 382.000 281.600 382.800 290.200 ;
        RECT 383.600 281.600 384.400 290.200 ;
        RECT 388.400 281.600 389.200 286.200 ;
        RECT 391.600 281.600 392.400 286.200 ;
        RECT 393.200 281.600 394.000 290.200 ;
        RECT 397.400 281.600 398.200 286.200 ;
        RECT 399.600 281.600 400.400 286.200 ;
        RECT 402.800 281.600 403.600 286.200 ;
        RECT 404.400 281.600 405.200 286.200 ;
        RECT 407.600 281.600 408.400 286.200 ;
        RECT 412.400 281.600 413.200 289.000 ;
        RECT 415.600 281.600 416.400 286.200 ;
        RECT 418.800 281.600 419.600 290.200 ;
        RECT 477.800 290.000 478.800 290.200 ;
        RECT 481.200 289.600 482.000 290.200 ;
        RECT 431.600 281.600 432.400 289.000 ;
        RECT 436.400 281.600 437.200 289.000 ;
        RECT 442.800 281.600 443.600 286.200 ;
        RECT 446.000 281.600 446.800 286.200 ;
        RECT 447.600 281.600 448.400 286.200 ;
        RECT 450.800 281.600 451.600 286.200 ;
        RECT 454.000 281.600 454.800 286.200 ;
        RECT 457.200 281.600 458.000 286.200 ;
        RECT 460.400 281.600 461.200 286.200 ;
        RECT 468.400 281.600 469.200 286.200 ;
        RECT 471.600 281.600 472.400 286.200 ;
        RECT 478.000 281.600 478.800 286.200 ;
        RECT 481.200 281.600 482.000 286.200 ;
        RECT 484.400 281.600 485.200 286.200 ;
        RECT 489.200 281.600 490.000 289.000 ;
        RECT 492.400 281.600 493.200 290.200 ;
        RECT 498.800 281.600 499.600 290.200 ;
        RECT 502.000 281.600 502.800 290.200 ;
        RECT 503.600 281.600 504.400 290.200 ;
        RECT 540.200 290.000 541.200 290.200 ;
        RECT 543.600 289.600 544.400 290.200 ;
        RECT 508.400 281.600 509.200 286.200 ;
        RECT 511.600 281.600 512.400 286.200 ;
        RECT 513.200 281.600 514.000 286.200 ;
        RECT 516.400 281.600 517.200 286.200 ;
        RECT 519.600 281.600 520.400 286.200 ;
        RECT 522.800 281.600 523.600 286.200 ;
        RECT 530.800 281.600 531.600 286.200 ;
        RECT 534.000 281.600 534.800 286.200 ;
        RECT 540.400 281.600 541.200 286.200 ;
        RECT 543.600 281.600 544.400 286.200 ;
        RECT 546.800 281.600 547.600 286.200 ;
        RECT 0.400 280.400 551.600 281.600 ;
        RECT 1.200 275.800 2.000 280.400 ;
        RECT 4.400 275.800 5.200 280.400 ;
        RECT 7.600 275.800 8.400 280.400 ;
        RECT 10.800 275.800 11.600 280.400 ;
        RECT 18.800 275.800 19.600 280.400 ;
        RECT 22.000 275.800 22.800 280.400 ;
        RECT 28.400 275.800 29.200 280.400 ;
        RECT 31.600 275.800 32.400 280.400 ;
        RECT 34.800 275.800 35.600 280.400 ;
        RECT 28.200 271.800 29.000 272.000 ;
        RECT 31.600 271.800 32.400 272.400 ;
        RECT 36.400 271.800 37.200 280.400 ;
        RECT 42.800 271.800 43.600 280.400 ;
        RECT 44.400 275.800 45.200 280.400 ;
        RECT 47.600 275.800 48.400 280.400 ;
        RECT 52.400 271.800 53.200 280.400 ;
        RECT 54.000 275.800 54.800 280.400 ;
        RECT 57.200 272.200 58.000 280.400 ;
        RECT 60.400 275.800 61.200 280.400 ;
        RECT 63.600 275.800 64.400 280.400 ;
        RECT 65.200 275.800 66.000 280.400 ;
        RECT 68.400 275.800 69.200 280.400 ;
        RECT 70.600 275.800 71.400 280.400 ;
        RECT 74.800 271.800 75.600 280.400 ;
        RECT 76.400 271.800 77.200 280.400 ;
        RECT 81.200 275.800 82.000 280.400 ;
        RECT 84.400 272.200 85.200 280.400 ;
        RECT 87.600 275.800 88.400 280.400 ;
        RECT 90.800 275.800 91.600 280.400 ;
        RECT 94.000 275.800 94.800 280.400 ;
        RECT 97.200 275.800 98.000 280.400 ;
        RECT 103.600 275.800 104.400 280.400 ;
        RECT 106.800 275.800 107.600 280.400 ;
        RECT 114.800 275.800 115.600 280.400 ;
        RECT 118.000 275.800 118.800 280.400 ;
        RECT 121.200 275.800 122.000 280.400 ;
        RECT 124.400 275.800 125.200 280.400 ;
        RECT 137.200 273.000 138.000 280.400 ;
        RECT 140.400 275.800 141.200 280.400 ;
        RECT 143.600 275.800 144.400 280.400 ;
        RECT 145.800 275.800 146.600 280.400 ;
        RECT 94.000 271.800 94.800 272.400 ;
        RECT 97.200 271.800 98.200 272.000 ;
        RECT 150.000 271.800 150.800 280.400 ;
        RECT 154.800 273.000 155.600 280.400 ;
        RECT 158.000 271.800 158.800 280.400 ;
        RECT 162.800 275.800 163.600 280.400 ;
        RECT 166.000 275.800 166.800 280.400 ;
        RECT 167.600 275.800 168.400 280.400 ;
        RECT 170.800 275.800 171.600 280.400 ;
        RECT 172.400 275.800 173.200 280.400 ;
        RECT 175.600 276.200 176.400 280.400 ;
        RECT 178.800 275.800 179.600 280.400 ;
        RECT 182.000 275.800 182.800 280.400 ;
        RECT 184.200 275.800 185.000 280.400 ;
        RECT 188.400 271.800 189.200 280.400 ;
        RECT 190.600 275.800 191.400 280.400 ;
        RECT 194.800 271.800 195.600 280.400 ;
        RECT 196.400 275.800 197.200 280.400 ;
        RECT 199.600 276.200 200.400 280.400 ;
        RECT 204.400 275.800 205.200 280.400 ;
        RECT 206.000 271.800 206.800 280.400 ;
        RECT 214.000 271.800 214.800 280.400 ;
        RECT 215.600 271.800 216.400 280.400 ;
        RECT 219.800 275.800 220.600 280.400 ;
        RECT 222.000 275.800 222.800 280.400 ;
        RECT 225.200 275.800 226.000 280.400 ;
        RECT 226.800 275.800 227.600 280.400 ;
        RECT 230.000 271.800 230.800 280.400 ;
        RECT 234.200 275.800 235.000 280.400 ;
        RECT 241.200 273.000 242.000 280.400 ;
        RECT 244.400 275.800 245.200 280.400 ;
        RECT 247.600 271.800 248.400 280.400 ;
        RECT 251.800 275.800 252.600 280.400 ;
        RECT 254.000 271.800 254.800 280.400 ;
        RECT 260.400 271.800 261.200 280.400 ;
        RECT 268.400 275.800 269.200 280.400 ;
        RECT 271.600 275.800 272.400 280.400 ;
        RECT 274.800 275.800 275.600 280.400 ;
        RECT 278.000 275.800 278.800 280.400 ;
        RECT 286.000 275.800 286.800 280.400 ;
        RECT 289.200 275.600 290.000 280.400 ;
        RECT 295.600 275.800 296.400 280.400 ;
        RECT 298.800 275.800 299.600 280.400 ;
        RECT 302.000 275.800 302.800 280.400 ;
        RECT 303.600 275.800 304.400 280.400 ;
        RECT 306.800 275.800 307.600 280.400 ;
        RECT 310.000 275.800 310.800 280.400 ;
        RECT 316.400 275.600 317.200 280.400 ;
        RECT 319.600 275.800 320.400 280.400 ;
        RECT 327.600 275.800 328.400 280.400 ;
        RECT 330.800 275.800 331.600 280.400 ;
        RECT 334.000 275.800 334.800 280.400 ;
        RECT 337.200 275.800 338.000 280.400 ;
        RECT 338.800 275.800 339.600 280.400 ;
        RECT 342.000 275.800 342.800 280.400 ;
        RECT 345.200 272.200 346.000 280.400 ;
        RECT 348.400 275.800 349.200 280.400 ;
        RECT 351.600 275.800 352.400 280.400 ;
        RECT 354.800 275.800 355.600 280.400 ;
        RECT 361.200 275.600 362.000 280.400 ;
        RECT 364.400 275.800 365.200 280.400 ;
        RECT 372.400 275.800 373.200 280.400 ;
        RECT 375.600 275.800 376.400 280.400 ;
        RECT 378.800 275.800 379.600 280.400 ;
        RECT 382.000 275.800 382.800 280.400 ;
        RECT 383.600 275.800 384.400 280.400 ;
        RECT 386.800 275.800 387.600 280.400 ;
        RECT 390.000 275.800 390.800 280.400 ;
        RECT 396.400 275.800 397.200 280.400 ;
        RECT 399.600 275.800 400.400 280.400 ;
        RECT 407.600 275.800 408.400 280.400 ;
        RECT 410.800 275.800 411.600 280.400 ;
        RECT 414.000 275.800 414.800 280.400 ;
        RECT 417.200 275.800 418.000 280.400 ;
        RECT 386.800 271.800 387.600 272.400 ;
        RECT 390.000 271.800 391.000 272.000 ;
        RECT 422.000 271.800 422.800 280.400 ;
        RECT 430.000 275.800 430.800 280.400 ;
        RECT 433.200 271.800 434.000 280.400 ;
        RECT 437.400 275.800 438.200 280.400 ;
        RECT 439.600 271.800 440.400 280.400 ;
        RECT 443.800 275.800 444.600 280.400 ;
        RECT 446.000 275.800 446.800 280.400 ;
        RECT 450.800 275.800 451.600 280.400 ;
        RECT 452.400 275.800 453.200 280.400 ;
        RECT 455.600 275.800 456.400 280.400 ;
        RECT 458.800 275.800 459.600 280.400 ;
        RECT 462.000 275.800 462.800 280.400 ;
        RECT 470.000 275.800 470.800 280.400 ;
        RECT 473.200 275.800 474.000 280.400 ;
        RECT 479.600 275.800 480.400 280.400 ;
        RECT 482.800 275.800 483.600 280.400 ;
        RECT 486.000 275.800 486.800 280.400 ;
        RECT 487.600 275.800 488.400 280.400 ;
        RECT 490.800 275.800 491.600 280.400 ;
        RECT 494.000 275.800 494.800 280.400 ;
        RECT 497.200 275.800 498.000 280.400 ;
        RECT 505.200 275.800 506.000 280.400 ;
        RECT 508.400 275.800 509.200 280.400 ;
        RECT 514.800 275.800 515.600 280.400 ;
        RECT 518.000 275.800 518.800 280.400 ;
        RECT 521.200 275.800 522.000 280.400 ;
        RECT 524.400 275.800 525.200 280.400 ;
        RECT 479.400 271.800 480.200 272.000 ;
        RECT 482.800 271.800 483.600 272.400 ;
        RECT 514.600 271.800 515.400 272.000 ;
        RECT 518.000 271.800 518.800 272.400 ;
        RECT 527.600 272.000 528.400 280.400 ;
        RECT 533.200 275.800 534.000 280.400 ;
        RECT 536.400 275.800 537.200 280.400 ;
        RECT 542.000 271.800 542.800 280.400 ;
        RECT 546.800 273.000 547.600 280.400 ;
        RECT 5.400 271.200 32.400 271.800 ;
        RECT 94.000 271.200 121.000 271.800 ;
        RECT 386.800 271.200 413.800 271.800 ;
        RECT 5.400 271.000 6.200 271.200 ;
        RECT 120.200 271.000 121.000 271.200 ;
        RECT 413.000 271.000 413.800 271.200 ;
        RECT 456.600 271.200 483.600 271.800 ;
        RECT 491.800 271.200 518.800 271.800 ;
        RECT 456.600 271.000 457.400 271.200 ;
        RECT 491.800 271.000 492.600 271.200 ;
        RECT 278.000 270.000 301.400 270.600 ;
        RECT 278.000 269.400 278.800 270.000 ;
        RECT 289.200 269.600 290.000 270.000 ;
        RECT 295.600 269.600 296.400 270.000 ;
        RECT 300.600 269.800 301.400 270.000 ;
        RECT 305.000 270.000 328.400 270.600 ;
        RECT 305.000 269.800 305.800 270.000 ;
        RECT 310.000 269.600 310.800 270.000 ;
        RECT 316.400 269.600 317.200 270.000 ;
        RECT 327.600 269.400 328.400 270.000 ;
        RECT 349.800 270.000 373.200 270.600 ;
        RECT 349.800 269.800 350.600 270.000 ;
        RECT 354.800 269.600 355.600 270.000 ;
        RECT 361.200 269.600 362.000 270.000 ;
        RECT 372.400 269.400 373.200 270.000 ;
        RECT 255.600 252.000 256.400 252.600 ;
        RECT 273.200 252.000 274.000 252.400 ;
        RECT 278.200 252.000 279.000 252.200 ;
        RECT 255.600 251.400 279.000 252.000 ;
        RECT 297.200 252.000 298.000 252.600 ;
        RECT 314.800 252.000 315.600 252.400 ;
        RECT 319.800 252.000 320.600 252.200 ;
        RECT 297.200 251.400 320.600 252.000 ;
        RECT 83.800 250.800 84.600 251.000 ;
        RECT 174.600 250.800 175.400 251.000 ;
        RECT 83.800 250.200 110.800 250.800 ;
        RECT 1.200 241.600 2.000 246.200 ;
        RECT 4.400 241.600 5.200 250.200 ;
        RECT 9.200 241.600 10.000 246.200 ;
        RECT 12.400 241.600 13.200 246.200 ;
        RECT 14.000 241.600 14.800 246.200 ;
        RECT 17.200 241.600 18.000 249.800 ;
        RECT 23.600 241.600 24.400 250.200 ;
        RECT 25.200 241.600 26.000 246.200 ;
        RECT 28.400 241.600 29.200 249.800 ;
        RECT 31.600 241.600 32.400 250.200 ;
        RECT 35.800 241.600 36.600 246.200 ;
        RECT 41.200 241.600 42.000 250.200 ;
        RECT 42.800 241.600 43.600 246.200 ;
        RECT 46.000 241.600 46.800 246.200 ;
        RECT 47.600 241.600 48.400 246.200 ;
        RECT 50.800 241.600 51.600 245.800 ;
        RECT 54.000 241.600 54.800 246.200 ;
        RECT 57.200 241.600 58.000 246.200 ;
        RECT 58.800 241.600 59.600 246.200 ;
        RECT 62.000 241.600 62.800 246.200 ;
        RECT 63.600 241.600 64.400 250.200 ;
        RECT 69.000 241.600 69.800 246.200 ;
        RECT 73.200 241.600 74.000 250.200 ;
        RECT 74.800 241.600 75.600 250.200 ;
        RECT 106.600 250.000 107.600 250.200 ;
        RECT 110.000 249.600 110.800 250.200 ;
        RECT 148.400 250.200 175.400 250.800 ;
        RECT 210.200 250.800 211.000 251.000 ;
        RECT 379.400 250.800 380.200 251.000 ;
        RECT 210.200 250.200 237.200 250.800 ;
        RECT 353.200 250.200 380.200 250.800 ;
        RECT 392.600 250.800 393.400 251.000 ;
        RECT 437.400 250.800 438.200 251.000 ;
        RECT 509.000 250.800 509.800 251.000 ;
        RECT 392.600 250.200 419.600 250.800 ;
        RECT 437.400 250.200 464.400 250.800 ;
        RECT 482.800 250.200 509.800 250.800 ;
        RECT 148.400 249.600 149.200 250.200 ;
        RECT 151.600 250.000 152.600 250.200 ;
        RECT 79.600 241.600 80.400 246.200 ;
        RECT 82.800 241.600 83.600 246.200 ;
        RECT 86.000 241.600 86.800 246.200 ;
        RECT 89.200 241.600 90.000 246.200 ;
        RECT 97.200 241.600 98.000 246.200 ;
        RECT 100.400 241.600 101.200 246.200 ;
        RECT 106.800 241.600 107.600 246.200 ;
        RECT 110.000 241.600 110.800 246.200 ;
        RECT 113.200 241.600 114.000 246.200 ;
        RECT 124.400 241.600 125.200 248.200 ;
        RECT 138.800 241.600 139.600 249.000 ;
        RECT 143.600 241.600 144.400 246.200 ;
        RECT 145.200 241.600 146.000 246.200 ;
        RECT 148.400 241.600 149.200 246.200 ;
        RECT 151.600 241.600 152.400 246.200 ;
        RECT 158.000 241.600 158.800 246.200 ;
        RECT 161.200 241.600 162.000 246.200 ;
        RECT 169.200 241.600 170.000 246.200 ;
        RECT 172.400 241.600 173.200 246.200 ;
        RECT 175.600 241.600 176.400 246.200 ;
        RECT 178.800 241.600 179.600 246.200 ;
        RECT 180.400 241.600 181.200 250.200 ;
        RECT 183.600 241.600 184.400 250.200 ;
        RECT 185.200 241.600 186.000 246.200 ;
        RECT 188.400 241.600 189.200 246.200 ;
        RECT 191.600 241.600 192.400 246.200 ;
        RECT 193.800 241.600 194.600 246.200 ;
        RECT 198.000 241.600 198.800 250.200 ;
        RECT 202.200 241.600 203.000 250.200 ;
        RECT 233.000 250.000 233.800 250.200 ;
        RECT 236.400 249.600 237.200 250.200 ;
        RECT 206.000 241.600 206.800 246.200 ;
        RECT 209.200 241.600 210.000 246.200 ;
        RECT 212.400 241.600 213.200 246.200 ;
        RECT 215.600 241.600 216.400 246.200 ;
        RECT 223.600 241.600 224.400 246.200 ;
        RECT 226.800 241.600 227.600 246.200 ;
        RECT 233.200 241.600 234.000 246.200 ;
        RECT 236.400 241.600 237.200 246.200 ;
        RECT 239.600 241.600 240.400 246.200 ;
        RECT 241.200 241.600 242.000 246.200 ;
        RECT 244.400 241.600 245.200 246.200 ;
        RECT 246.000 241.600 246.800 246.200 ;
        RECT 249.200 241.600 250.000 246.200 ;
        RECT 252.400 241.600 253.200 246.200 ;
        RECT 255.600 241.600 256.400 246.200 ;
        RECT 263.600 241.600 264.400 246.200 ;
        RECT 266.800 241.600 267.600 246.200 ;
        RECT 273.200 241.600 274.000 246.200 ;
        RECT 276.400 241.600 277.200 246.200 ;
        RECT 279.600 241.600 280.400 246.200 ;
        RECT 287.600 241.600 288.400 246.200 ;
        RECT 290.800 241.600 291.600 246.200 ;
        RECT 294.000 241.600 294.800 246.200 ;
        RECT 297.200 241.600 298.000 246.200 ;
        RECT 305.200 241.600 306.000 246.200 ;
        RECT 308.400 241.600 309.200 246.200 ;
        RECT 314.800 241.600 315.600 246.200 ;
        RECT 318.000 241.600 318.800 246.200 ;
        RECT 321.200 241.600 322.000 246.200 ;
        RECT 323.400 241.600 324.200 246.200 ;
        RECT 327.600 241.600 328.400 250.200 ;
        RECT 329.800 241.600 330.600 246.200 ;
        RECT 334.000 241.600 334.800 250.200 ;
        RECT 335.600 241.600 336.400 250.200 ;
        RECT 338.800 241.600 339.600 250.200 ;
        RECT 340.400 241.600 341.200 246.200 ;
        RECT 343.600 241.600 344.400 250.200 ;
        RECT 353.200 249.600 354.000 250.200 ;
        RECT 356.400 250.000 357.400 250.200 ;
        RECT 415.400 250.000 416.400 250.200 ;
        RECT 418.800 249.600 419.600 250.200 ;
        RECT 460.200 250.000 461.200 250.200 ;
        RECT 463.600 249.600 464.400 250.200 ;
        RECT 347.800 241.600 348.600 246.200 ;
        RECT 350.000 241.600 350.800 246.200 ;
        RECT 353.200 241.600 354.000 246.200 ;
        RECT 356.400 241.600 357.200 246.200 ;
        RECT 362.800 241.600 363.600 246.200 ;
        RECT 366.000 241.600 366.800 246.200 ;
        RECT 374.000 241.600 374.800 246.200 ;
        RECT 377.200 241.600 378.000 246.200 ;
        RECT 380.400 241.600 381.200 246.200 ;
        RECT 383.600 241.600 384.400 246.200 ;
        RECT 386.800 241.600 387.600 246.200 ;
        RECT 388.400 241.600 389.200 246.200 ;
        RECT 391.600 241.600 392.400 246.200 ;
        RECT 394.800 241.600 395.600 246.200 ;
        RECT 398.000 241.600 398.800 246.200 ;
        RECT 406.000 241.600 406.800 246.200 ;
        RECT 409.200 241.600 410.000 246.200 ;
        RECT 415.600 241.600 416.400 246.200 ;
        RECT 418.800 241.600 419.600 246.200 ;
        RECT 422.000 241.600 422.800 246.200 ;
        RECT 430.000 241.600 430.800 246.200 ;
        RECT 433.200 241.600 434.000 246.200 ;
        RECT 436.400 241.600 437.200 246.200 ;
        RECT 439.600 241.600 440.400 246.200 ;
        RECT 442.800 241.600 443.600 246.200 ;
        RECT 450.800 241.600 451.600 246.200 ;
        RECT 454.000 241.600 454.800 246.200 ;
        RECT 460.400 241.600 461.200 246.200 ;
        RECT 463.600 241.600 464.400 246.200 ;
        RECT 466.800 241.600 467.600 246.200 ;
        RECT 471.600 241.600 472.400 249.000 ;
        RECT 478.000 241.600 478.800 250.200 ;
        RECT 482.800 249.600 483.600 250.200 ;
        RECT 486.000 250.000 487.000 250.200 ;
        RECT 479.600 241.600 480.400 246.200 ;
        RECT 482.800 241.600 483.600 246.200 ;
        RECT 486.000 241.600 486.800 246.200 ;
        RECT 492.400 241.600 493.200 246.200 ;
        RECT 495.600 241.600 496.400 246.200 ;
        RECT 503.600 241.600 504.400 246.200 ;
        RECT 506.800 241.600 507.600 246.200 ;
        RECT 510.000 241.600 510.800 246.200 ;
        RECT 513.200 241.600 514.000 246.200 ;
        RECT 514.800 241.600 515.600 250.200 ;
        RECT 518.000 241.600 518.800 250.200 ;
        RECT 521.200 241.600 522.000 250.200 ;
        RECT 524.400 241.600 525.200 250.200 ;
        RECT 527.600 241.600 528.400 250.200 ;
        RECT 530.800 241.600 531.600 250.200 ;
        RECT 536.400 241.600 537.200 246.200 ;
        RECT 539.600 241.600 540.400 246.200 ;
        RECT 545.200 241.600 546.000 250.000 ;
        RECT 0.400 240.400 551.600 241.600 ;
        RECT 1.200 235.800 2.000 240.400 ;
        RECT 4.400 235.800 5.200 240.400 ;
        RECT 7.600 235.800 8.400 240.400 ;
        RECT 10.800 235.800 11.600 240.400 ;
        RECT 18.800 235.800 19.600 240.400 ;
        RECT 22.000 235.800 22.800 240.400 ;
        RECT 28.400 235.800 29.200 240.400 ;
        RECT 31.600 235.800 32.400 240.400 ;
        RECT 34.800 235.800 35.600 240.400 ;
        RECT 36.400 235.800 37.200 240.400 ;
        RECT 39.600 236.200 40.400 240.400 ;
        RECT 28.200 231.800 29.000 232.000 ;
        RECT 31.600 231.800 32.400 232.400 ;
        RECT 42.800 231.800 43.600 240.400 ;
        RECT 49.200 231.800 50.000 240.400 ;
        RECT 54.000 231.800 54.800 240.400 ;
        RECT 57.200 232.200 58.000 240.400 ;
        RECT 60.400 235.800 61.200 240.400 ;
        RECT 62.000 235.800 62.800 240.400 ;
        RECT 65.200 235.800 66.000 240.400 ;
        RECT 68.400 236.200 69.200 240.400 ;
        RECT 71.600 235.800 72.400 240.400 ;
        RECT 73.200 235.800 74.000 240.400 ;
        RECT 76.400 232.200 77.200 240.400 ;
        RECT 82.800 233.000 83.600 240.400 ;
        RECT 86.000 231.800 86.800 240.400 ;
        RECT 90.800 235.800 91.600 240.400 ;
        RECT 94.000 232.200 94.800 240.400 ;
        RECT 100.400 233.000 101.200 240.400 ;
        RECT 103.600 235.800 104.400 240.400 ;
        RECT 106.800 235.800 107.600 240.400 ;
        RECT 110.000 235.800 110.800 240.400 ;
        RECT 113.200 235.800 114.000 240.400 ;
        RECT 121.200 235.800 122.000 240.400 ;
        RECT 124.400 235.800 125.200 240.400 ;
        RECT 130.800 235.800 131.600 240.400 ;
        RECT 134.000 235.800 134.800 240.400 ;
        RECT 137.200 235.800 138.000 240.400 ;
        RECT 130.600 231.800 131.600 232.000 ;
        RECT 134.000 231.800 134.800 232.400 ;
        RECT 145.200 231.800 146.000 240.400 ;
        RECT 148.400 231.800 149.200 240.400 ;
        RECT 151.600 235.800 152.400 240.400 ;
        RECT 153.800 235.800 154.600 240.400 ;
        RECT 158.000 231.800 158.800 240.400 ;
        RECT 159.600 231.800 160.400 240.400 ;
        RECT 163.800 235.800 164.600 240.400 ;
        RECT 166.000 235.800 166.800 240.400 ;
        RECT 169.200 235.800 170.000 240.400 ;
        RECT 170.800 235.800 171.600 240.400 ;
        RECT 174.000 232.200 174.800 240.400 ;
        RECT 177.200 235.800 178.000 240.400 ;
        RECT 180.400 235.800 181.200 240.400 ;
        RECT 183.600 233.000 184.400 240.400 ;
        RECT 186.800 235.800 187.600 240.400 ;
        RECT 190.000 235.800 190.800 240.400 ;
        RECT 192.200 235.800 193.000 240.400 ;
        RECT 196.400 231.800 197.200 240.400 ;
        RECT 198.000 231.800 198.800 240.400 ;
        RECT 202.200 235.800 203.000 240.400 ;
        RECT 204.400 235.800 205.200 240.400 ;
        RECT 207.600 235.800 208.400 240.400 ;
        RECT 210.800 235.800 211.600 240.400 ;
        RECT 214.000 235.800 214.800 240.400 ;
        RECT 222.000 235.800 222.800 240.400 ;
        RECT 225.200 235.800 226.000 240.400 ;
        RECT 231.600 235.800 232.400 240.400 ;
        RECT 234.800 235.800 235.600 240.400 ;
        RECT 238.000 235.800 238.800 240.400 ;
        RECT 239.600 235.800 240.400 240.400 ;
        RECT 242.800 235.800 243.600 240.400 ;
        RECT 246.000 235.800 246.800 240.400 ;
        RECT 249.200 235.800 250.000 240.400 ;
        RECT 257.200 235.800 258.000 240.400 ;
        RECT 260.400 235.800 261.200 240.400 ;
        RECT 266.800 235.800 267.600 240.400 ;
        RECT 270.000 235.800 270.800 240.400 ;
        RECT 273.200 235.800 274.000 240.400 ;
        RECT 281.200 235.800 282.000 240.400 ;
        RECT 284.400 235.800 285.200 240.400 ;
        RECT 287.600 235.800 288.400 240.400 ;
        RECT 290.800 235.800 291.600 240.400 ;
        RECT 294.000 235.800 294.800 240.400 ;
        RECT 302.000 235.800 302.800 240.400 ;
        RECT 305.200 235.600 306.000 240.400 ;
        RECT 311.600 235.800 312.400 240.400 ;
        RECT 314.800 235.800 315.600 240.400 ;
        RECT 318.000 235.800 318.800 240.400 ;
        RECT 231.400 231.800 232.200 232.000 ;
        RECT 234.800 231.800 235.600 232.400 ;
        RECT 266.600 231.800 267.600 232.000 ;
        RECT 270.000 231.800 270.800 232.400 ;
        RECT 319.600 231.800 320.400 240.400 ;
        RECT 323.800 235.800 324.600 240.400 ;
        RECT 326.000 231.800 326.800 240.400 ;
        RECT 330.200 235.800 331.000 240.400 ;
        RECT 333.000 235.800 333.800 240.400 ;
        RECT 337.200 231.800 338.000 240.400 ;
        RECT 339.400 235.800 340.200 240.400 ;
        RECT 343.600 231.800 344.400 240.400 ;
        RECT 346.800 233.000 347.600 240.400 ;
        RECT 351.600 233.000 352.400 240.400 ;
        RECT 354.800 231.800 355.600 240.400 ;
        RECT 359.000 235.800 359.800 240.400 ;
        RECT 362.800 233.000 363.600 240.400 ;
        RECT 366.600 235.800 367.400 240.400 ;
        RECT 370.800 231.800 371.600 240.400 ;
        RECT 372.400 235.800 373.200 240.400 ;
        RECT 375.600 235.800 376.400 240.400 ;
        RECT 377.200 235.800 378.000 240.400 ;
        RECT 380.400 235.800 381.200 240.400 ;
        RECT 383.600 235.800 384.400 240.400 ;
        RECT 386.800 235.800 387.600 240.400 ;
        RECT 394.800 235.800 395.600 240.400 ;
        RECT 398.000 235.800 398.800 240.400 ;
        RECT 404.400 235.800 405.200 240.400 ;
        RECT 407.600 235.800 408.400 240.400 ;
        RECT 410.800 235.800 411.600 240.400 ;
        RECT 412.400 235.800 413.200 240.400 ;
        RECT 404.200 231.800 405.200 232.000 ;
        RECT 407.600 231.800 408.400 232.400 ;
        RECT 415.600 231.800 416.400 240.400 ;
        RECT 419.800 235.800 420.600 240.400 ;
        RECT 428.400 235.800 429.200 240.400 ;
        RECT 431.600 236.200 432.400 240.400 ;
        RECT 438.000 231.800 438.800 240.400 ;
        RECT 439.600 235.800 440.400 240.400 ;
        RECT 442.800 236.200 443.600 240.400 ;
        RECT 446.000 235.800 446.800 240.400 ;
        RECT 449.200 235.800 450.000 240.400 ;
        RECT 450.800 231.800 451.600 240.400 ;
        RECT 455.000 235.800 455.800 240.400 ;
        RECT 457.200 235.800 458.000 240.400 ;
        RECT 460.400 236.200 461.200 240.400 ;
        RECT 463.600 235.800 464.400 240.400 ;
        RECT 466.800 236.200 467.600 240.400 ;
        RECT 470.000 231.800 470.800 240.400 ;
        RECT 474.800 231.800 475.600 240.400 ;
        RECT 481.200 233.000 482.000 240.400 ;
        RECT 486.000 235.800 486.800 240.400 ;
        RECT 489.200 235.800 490.000 240.400 ;
        RECT 490.800 235.800 491.600 240.400 ;
        RECT 494.000 235.800 494.800 240.400 ;
        RECT 495.600 235.800 496.400 240.400 ;
        RECT 498.800 235.800 499.600 240.400 ;
        RECT 502.000 235.800 502.800 240.400 ;
        RECT 505.200 235.800 506.000 240.400 ;
        RECT 513.200 235.800 514.000 240.400 ;
        RECT 516.400 235.800 517.200 240.400 ;
        RECT 522.800 235.800 523.600 240.400 ;
        RECT 526.000 235.800 526.800 240.400 ;
        RECT 529.200 235.800 530.000 240.400 ;
        RECT 534.000 233.000 534.800 240.400 ;
        RECT 537.200 235.800 538.000 240.400 ;
        RECT 540.400 235.800 541.200 240.400 ;
        RECT 522.600 231.800 523.400 232.000 ;
        RECT 526.000 231.800 526.800 232.400 ;
        RECT 542.000 231.800 542.800 240.400 ;
        RECT 548.400 233.000 549.200 240.400 ;
        RECT 5.400 231.200 32.400 231.800 ;
        RECT 107.800 231.200 134.800 231.800 ;
        RECT 208.600 231.200 235.600 231.800 ;
        RECT 243.800 231.200 270.800 231.800 ;
        RECT 381.400 231.200 408.400 231.800 ;
        RECT 499.800 231.200 526.800 231.800 ;
        RECT 5.400 231.000 6.200 231.200 ;
        RECT 107.800 231.000 108.600 231.200 ;
        RECT 208.600 231.000 209.400 231.200 ;
        RECT 243.800 231.000 244.600 231.200 ;
        RECT 381.400 231.000 382.200 231.200 ;
        RECT 499.800 231.000 500.600 231.200 ;
        RECT 294.000 230.000 317.400 230.600 ;
        RECT 294.000 229.400 294.800 230.000 ;
        RECT 305.200 229.600 306.000 230.000 ;
        RECT 311.600 229.600 312.400 230.000 ;
        RECT 316.600 229.800 317.400 230.000 ;
        RECT 300.400 212.000 301.200 212.600 ;
        RECT 318.000 212.000 318.800 212.400 ;
        RECT 323.000 212.000 323.800 212.200 ;
        RECT 300.400 211.400 323.800 212.000 ;
        RECT 145.800 210.800 146.600 211.000 ;
        RECT 119.600 210.200 146.600 210.800 ;
        RECT 250.200 210.800 251.000 211.000 ;
        RECT 483.800 210.800 484.600 211.000 ;
        RECT 544.200 210.800 545.000 211.000 ;
        RECT 250.200 210.200 277.200 210.800 ;
        RECT 483.800 210.200 510.800 210.800 ;
        RECT 1.200 201.600 2.000 210.200 ;
        RECT 4.400 201.600 5.200 210.200 ;
        RECT 6.000 201.600 6.800 210.200 ;
        RECT 12.400 201.600 13.200 209.000 ;
        RECT 18.800 201.600 19.600 206.200 ;
        RECT 22.000 201.600 22.800 206.200 ;
        RECT 25.200 201.600 26.000 205.800 ;
        RECT 28.400 201.600 29.200 206.200 ;
        RECT 30.000 201.600 30.800 206.200 ;
        RECT 33.200 201.600 34.000 209.800 ;
        RECT 36.400 201.600 37.200 206.200 ;
        RECT 39.600 201.600 40.400 209.800 ;
        RECT 44.400 201.600 45.200 205.800 ;
        RECT 47.600 201.600 48.400 206.200 ;
        RECT 50.800 201.600 51.600 208.200 ;
        RECT 62.000 201.600 62.800 206.200 ;
        RECT 65.200 201.600 66.000 205.800 ;
        RECT 68.400 201.600 69.200 206.200 ;
        RECT 71.600 201.600 72.400 205.800 ;
        RECT 74.800 201.600 75.600 206.200 ;
        RECT 78.000 201.600 78.800 205.800 ;
        RECT 83.800 201.600 84.600 210.200 ;
        RECT 87.600 201.600 88.400 206.200 ;
        RECT 90.800 201.600 91.600 206.200 ;
        RECT 94.000 201.600 94.800 209.000 ;
        RECT 98.800 201.600 99.600 206.200 ;
        RECT 102.000 201.600 102.800 206.200 ;
        RECT 103.600 201.600 104.400 210.200 ;
        RECT 119.600 209.600 120.400 210.200 ;
        RECT 123.000 210.000 123.800 210.200 ;
        RECT 107.800 201.600 108.600 206.200 ;
        RECT 116.400 201.600 117.200 206.200 ;
        RECT 119.600 201.600 120.400 206.200 ;
        RECT 122.800 201.600 123.600 206.200 ;
        RECT 129.200 201.600 130.000 206.200 ;
        RECT 132.400 201.600 133.200 206.200 ;
        RECT 140.400 201.600 141.200 206.200 ;
        RECT 143.600 201.600 144.400 206.200 ;
        RECT 146.800 201.600 147.600 206.200 ;
        RECT 150.000 201.600 150.800 206.200 ;
        RECT 154.800 201.600 155.600 210.200 ;
        RECT 156.400 201.600 157.200 206.200 ;
        RECT 159.600 201.600 160.400 206.200 ;
        RECT 161.200 201.600 162.000 210.200 ;
        RECT 165.400 201.600 166.200 206.200 ;
        RECT 172.400 201.600 173.200 209.000 ;
        RECT 177.200 201.600 178.000 206.200 ;
        RECT 178.800 201.600 179.600 206.200 ;
        RECT 182.000 201.600 182.800 209.800 ;
        RECT 188.400 201.600 189.200 210.200 ;
        RECT 190.000 201.600 190.800 210.200 ;
        RECT 194.200 201.600 195.000 206.200 ;
        RECT 196.400 201.600 197.200 206.200 ;
        RECT 199.600 201.600 200.400 206.200 ;
        RECT 202.800 201.600 203.600 205.800 ;
        RECT 206.000 201.600 206.800 206.200 ;
        RECT 212.400 201.600 213.200 209.000 ;
        RECT 215.600 201.600 216.400 206.200 ;
        RECT 218.800 201.600 219.600 206.200 ;
        RECT 220.400 201.600 221.200 210.200 ;
        RECT 224.600 201.600 225.400 206.200 ;
        RECT 226.800 201.600 227.600 210.200 ;
        RECT 231.000 201.600 231.800 206.200 ;
        RECT 234.800 201.600 235.600 209.000 ;
        RECT 240.200 201.600 241.000 206.200 ;
        RECT 244.400 201.600 245.200 210.200 ;
        RECT 273.000 210.000 274.000 210.200 ;
        RECT 276.400 209.600 277.200 210.200 ;
        RECT 246.000 201.600 246.800 206.200 ;
        RECT 249.200 201.600 250.000 206.200 ;
        RECT 252.400 201.600 253.200 206.200 ;
        RECT 255.600 201.600 256.400 206.200 ;
        RECT 263.600 201.600 264.400 206.200 ;
        RECT 266.800 201.600 267.600 206.200 ;
        RECT 273.200 201.600 274.000 206.200 ;
        RECT 276.400 201.600 277.200 206.200 ;
        RECT 279.600 201.600 280.400 206.200 ;
        RECT 287.600 201.600 288.400 206.200 ;
        RECT 290.800 201.600 291.600 206.200 ;
        RECT 294.000 201.600 294.800 206.200 ;
        RECT 297.200 201.600 298.000 206.200 ;
        RECT 300.400 201.600 301.200 206.200 ;
        RECT 308.400 201.600 309.200 206.200 ;
        RECT 311.600 201.600 312.400 206.200 ;
        RECT 318.000 201.600 318.800 206.200 ;
        RECT 321.200 201.600 322.000 206.200 ;
        RECT 324.400 201.600 325.200 206.200 ;
        RECT 326.000 201.600 326.800 206.200 ;
        RECT 329.200 201.600 330.000 210.200 ;
        RECT 333.400 201.600 334.200 206.200 ;
        RECT 336.200 201.600 337.000 206.200 ;
        RECT 340.400 201.600 341.200 210.200 ;
        RECT 342.000 201.600 342.800 206.200 ;
        RECT 346.800 201.600 347.600 210.200 ;
        RECT 352.400 201.600 353.200 206.200 ;
        RECT 355.600 201.600 356.400 206.200 ;
        RECT 361.200 201.600 362.000 210.000 ;
        RECT 365.000 201.600 365.800 206.200 ;
        RECT 369.200 201.600 370.000 210.200 ;
        RECT 370.800 201.600 371.600 210.200 ;
        RECT 377.200 201.600 378.000 210.200 ;
        RECT 382.000 201.600 382.800 209.000 ;
        RECT 385.200 201.600 386.000 206.200 ;
        RECT 388.400 201.600 389.200 206.200 ;
        RECT 390.000 201.600 390.800 210.200 ;
        RECT 394.200 201.600 395.000 206.200 ;
        RECT 396.400 201.600 397.200 210.200 ;
        RECT 402.800 201.600 403.600 210.200 ;
        RECT 404.400 201.600 405.200 210.200 ;
        RECT 410.800 201.600 411.600 210.200 ;
        RECT 415.600 201.600 416.400 210.200 ;
        RECT 417.800 201.600 418.600 206.200 ;
        RECT 422.000 201.600 422.800 210.200 ;
        RECT 434.800 201.600 435.600 209.000 ;
        RECT 438.000 201.600 438.800 210.200 ;
        RECT 446.000 201.600 446.800 210.200 ;
        RECT 447.600 201.600 448.400 210.200 ;
        RECT 454.000 201.600 454.800 210.200 ;
        RECT 455.600 201.600 456.400 210.200 ;
        RECT 462.000 201.600 462.800 210.200 ;
        RECT 465.200 201.600 466.000 209.800 ;
        RECT 470.400 201.600 471.200 210.200 ;
        RECT 473.200 201.600 474.000 210.200 ;
        RECT 506.600 210.000 507.400 210.200 ;
        RECT 510.000 209.600 510.800 210.200 ;
        RECT 518.000 210.200 545.000 210.800 ;
        RECT 518.000 209.600 518.800 210.200 ;
        RECT 521.200 210.000 522.200 210.200 ;
        RECT 477.400 201.600 478.200 206.200 ;
        RECT 479.600 201.600 480.400 206.200 ;
        RECT 482.800 201.600 483.600 206.200 ;
        RECT 486.000 201.600 486.800 206.200 ;
        RECT 489.200 201.600 490.000 206.200 ;
        RECT 497.200 201.600 498.000 206.200 ;
        RECT 500.400 201.600 501.200 206.200 ;
        RECT 506.800 201.600 507.600 206.200 ;
        RECT 510.000 201.600 510.800 206.200 ;
        RECT 513.200 201.600 514.000 206.200 ;
        RECT 514.800 201.600 515.600 206.200 ;
        RECT 518.000 201.600 518.800 206.200 ;
        RECT 521.200 201.600 522.000 206.200 ;
        RECT 527.600 201.600 528.400 206.200 ;
        RECT 530.800 201.600 531.600 206.200 ;
        RECT 538.800 201.600 539.600 206.200 ;
        RECT 542.000 201.600 542.800 206.200 ;
        RECT 545.200 201.600 546.000 206.200 ;
        RECT 548.400 201.600 549.200 206.200 ;
        RECT 0.400 200.400 551.600 201.600 ;
        RECT 1.200 195.800 2.000 200.400 ;
        RECT 4.400 195.800 5.200 200.400 ;
        RECT 6.000 195.800 6.800 200.400 ;
        RECT 9.200 195.800 10.000 200.400 ;
        RECT 14.000 191.800 14.800 200.400 ;
        RECT 15.600 195.800 16.400 200.400 ;
        RECT 18.800 192.200 19.600 200.400 ;
        RECT 22.000 191.800 22.800 200.400 ;
        RECT 29.400 191.800 30.200 200.400 ;
        RECT 33.200 195.800 34.000 200.400 ;
        RECT 36.400 196.200 37.200 200.400 ;
        RECT 41.200 196.200 42.000 200.400 ;
        RECT 44.400 195.800 45.200 200.400 ;
        RECT 46.000 195.800 46.800 200.400 ;
        RECT 49.200 195.800 50.000 200.400 ;
        RECT 52.400 195.800 53.200 200.400 ;
        RECT 55.600 196.200 56.400 200.400 ;
        RECT 58.800 195.800 59.600 200.400 ;
        RECT 60.400 195.800 61.200 200.400 ;
        RECT 63.600 192.200 64.400 200.400 ;
        RECT 66.800 195.800 67.600 200.400 ;
        RECT 70.000 195.800 70.800 200.400 ;
        RECT 73.200 195.800 74.000 200.400 ;
        RECT 79.600 195.800 80.400 200.400 ;
        RECT 82.800 195.800 83.600 200.400 ;
        RECT 90.800 195.800 91.600 200.400 ;
        RECT 94.000 195.800 94.800 200.400 ;
        RECT 97.200 195.800 98.000 200.400 ;
        RECT 100.400 195.800 101.200 200.400 ;
        RECT 102.000 195.800 102.800 200.400 ;
        RECT 105.200 195.800 106.000 200.400 ;
        RECT 108.400 195.800 109.200 200.400 ;
        RECT 111.600 195.800 112.400 200.400 ;
        RECT 119.600 195.800 120.400 200.400 ;
        RECT 122.800 195.600 123.600 200.400 ;
        RECT 129.200 195.800 130.000 200.400 ;
        RECT 132.400 195.800 133.200 200.400 ;
        RECT 135.600 195.800 136.400 200.400 ;
        RECT 143.600 195.800 144.400 200.400 ;
        RECT 146.800 195.800 147.600 200.400 ;
        RECT 150.000 195.800 150.800 200.400 ;
        RECT 156.400 195.800 157.200 200.400 ;
        RECT 159.600 195.800 160.400 200.400 ;
        RECT 167.600 195.800 168.400 200.400 ;
        RECT 170.800 195.800 171.600 200.400 ;
        RECT 174.000 195.800 174.800 200.400 ;
        RECT 177.200 195.800 178.000 200.400 ;
        RECT 70.000 191.800 70.800 192.400 ;
        RECT 73.200 191.800 74.200 192.000 ;
        RECT 146.800 191.800 147.600 192.400 ;
        RECT 150.200 191.800 151.000 192.000 ;
        RECT 180.400 191.800 181.200 200.400 ;
        RECT 182.000 195.800 182.800 200.400 ;
        RECT 185.200 195.800 186.000 200.400 ;
        RECT 188.400 195.800 189.200 200.400 ;
        RECT 191.600 195.800 192.400 200.400 ;
        RECT 199.600 195.800 200.400 200.400 ;
        RECT 202.800 195.800 203.600 200.400 ;
        RECT 209.200 195.800 210.000 200.400 ;
        RECT 212.400 195.800 213.200 200.400 ;
        RECT 215.600 195.800 216.400 200.400 ;
        RECT 218.800 195.800 219.600 200.400 ;
        RECT 222.000 196.200 222.800 200.400 ;
        RECT 225.200 195.800 226.000 200.400 ;
        RECT 228.400 195.800 229.200 200.400 ;
        RECT 230.000 195.800 230.800 200.400 ;
        RECT 233.200 195.800 234.000 200.400 ;
        RECT 209.000 191.800 209.800 192.000 ;
        RECT 212.400 191.800 213.200 192.400 ;
        RECT 238.000 191.800 238.800 200.400 ;
        RECT 239.600 195.800 240.400 200.400 ;
        RECT 242.800 195.800 243.600 200.400 ;
        RECT 244.400 195.800 245.200 200.400 ;
        RECT 247.600 191.800 248.400 200.400 ;
        RECT 251.800 195.800 252.600 200.400 ;
        RECT 255.600 193.000 256.400 200.400 ;
        RECT 266.800 195.800 267.600 200.400 ;
        RECT 270.000 195.800 270.800 200.400 ;
        RECT 273.200 195.800 274.000 200.400 ;
        RECT 276.400 195.800 277.200 200.400 ;
        RECT 284.400 195.800 285.200 200.400 ;
        RECT 287.600 195.800 288.400 200.400 ;
        RECT 294.000 195.800 294.800 200.400 ;
        RECT 297.200 195.800 298.000 200.400 ;
        RECT 300.400 195.800 301.200 200.400 ;
        RECT 302.000 195.800 302.800 200.400 ;
        RECT 305.200 195.800 306.000 200.400 ;
        RECT 308.400 195.800 309.200 200.400 ;
        RECT 311.600 195.800 312.400 200.400 ;
        RECT 319.600 195.800 320.400 200.400 ;
        RECT 322.800 195.600 323.600 200.400 ;
        RECT 329.200 195.800 330.000 200.400 ;
        RECT 332.400 195.800 333.200 200.400 ;
        RECT 335.600 195.800 336.400 200.400 ;
        RECT 337.200 195.800 338.000 200.400 ;
        RECT 293.800 191.800 294.800 192.000 ;
        RECT 297.200 191.800 298.000 192.400 ;
        RECT 340.400 191.800 341.200 200.400 ;
        RECT 344.600 195.800 345.400 200.400 ;
        RECT 346.800 195.800 347.600 200.400 ;
        RECT 350.000 195.800 350.800 200.400 ;
        RECT 353.200 195.800 354.000 200.400 ;
        RECT 359.600 195.600 360.400 200.400 ;
        RECT 362.800 195.800 363.600 200.400 ;
        RECT 370.800 195.800 371.600 200.400 ;
        RECT 374.000 195.800 374.800 200.400 ;
        RECT 377.200 195.800 378.000 200.400 ;
        RECT 380.400 195.800 381.200 200.400 ;
        RECT 382.600 195.800 383.400 200.400 ;
        RECT 386.800 191.800 387.600 200.400 ;
        RECT 388.400 195.800 389.200 200.400 ;
        RECT 391.600 196.200 392.400 200.400 ;
        RECT 394.800 195.800 395.600 200.400 ;
        RECT 398.000 195.800 398.800 200.400 ;
        RECT 399.600 191.800 400.400 200.400 ;
        RECT 403.800 195.800 404.600 200.400 ;
        RECT 406.000 195.800 406.800 200.400 ;
        RECT 409.200 195.800 410.000 200.400 ;
        RECT 412.400 196.200 413.200 200.400 ;
        RECT 417.200 195.800 418.000 200.400 ;
        RECT 418.800 191.800 419.600 200.400 ;
        RECT 423.000 195.800 423.800 200.400 ;
        RECT 433.200 195.800 434.000 200.400 ;
        RECT 436.400 192.200 437.200 200.400 ;
        RECT 441.600 191.800 442.400 200.400 ;
        RECT 446.000 196.200 446.800 200.400 ;
        RECT 449.200 195.800 450.000 200.400 ;
        RECT 452.400 193.000 453.200 200.400 ;
        RECT 457.200 196.200 458.000 200.400 ;
        RECT 460.400 195.800 461.200 200.400 ;
        RECT 462.600 195.800 463.400 200.400 ;
        RECT 466.800 191.800 467.600 200.400 ;
        RECT 468.400 195.800 469.200 200.400 ;
        RECT 471.600 195.800 472.400 200.400 ;
        RECT 474.800 195.800 475.600 200.400 ;
        RECT 478.000 195.800 478.800 200.400 ;
        RECT 486.000 195.800 486.800 200.400 ;
        RECT 489.200 195.800 490.000 200.400 ;
        RECT 495.600 195.800 496.400 200.400 ;
        RECT 498.800 195.800 499.600 200.400 ;
        RECT 502.000 195.800 502.800 200.400 ;
        RECT 495.400 191.800 496.200 192.000 ;
        RECT 498.800 191.800 499.600 192.400 ;
        RECT 503.600 191.800 504.400 200.400 ;
        RECT 510.000 191.800 510.800 200.400 ;
        RECT 513.200 192.200 514.000 200.400 ;
        RECT 518.400 191.800 519.200 200.400 ;
        RECT 522.800 192.000 523.600 200.400 ;
        RECT 528.400 195.800 529.200 200.400 ;
        RECT 531.600 195.800 532.400 200.400 ;
        RECT 537.200 191.800 538.000 200.400 ;
        RECT 540.400 191.800 541.200 200.400 ;
        RECT 544.600 195.800 545.400 200.400 ;
        RECT 546.800 195.800 547.600 200.400 ;
        RECT 550.000 195.800 550.800 200.400 ;
        RECT 70.000 191.200 97.000 191.800 ;
        RECT 146.800 191.200 173.800 191.800 ;
        RECT 96.200 191.000 97.000 191.200 ;
        RECT 173.000 191.000 173.800 191.200 ;
        RECT 186.200 191.200 213.200 191.800 ;
        RECT 271.000 191.200 298.000 191.800 ;
        RECT 472.600 191.200 499.600 191.800 ;
        RECT 186.200 191.000 187.000 191.200 ;
        RECT 271.000 191.000 271.800 191.200 ;
        RECT 472.600 191.000 473.400 191.200 ;
        RECT 111.600 190.000 135.000 190.600 ;
        RECT 111.600 189.400 112.400 190.000 ;
        RECT 122.800 189.600 123.600 190.000 ;
        RECT 129.200 189.600 130.000 190.000 ;
        RECT 134.200 189.800 135.000 190.000 ;
        RECT 311.600 190.000 335.000 190.600 ;
        RECT 311.600 189.400 312.400 190.000 ;
        RECT 322.800 189.600 323.600 190.000 ;
        RECT 329.200 189.600 330.000 190.000 ;
        RECT 334.200 189.800 335.000 190.000 ;
        RECT 348.200 190.000 371.600 190.600 ;
        RECT 348.200 189.800 349.000 190.000 ;
        RECT 353.200 189.600 354.000 190.000 ;
        RECT 359.600 189.600 360.400 190.000 ;
        RECT 370.800 189.400 371.600 190.000 ;
        RECT 126.000 172.000 126.800 172.600 ;
        RECT 143.600 172.000 144.400 172.400 ;
        RECT 148.600 172.000 149.400 172.200 ;
        RECT 126.000 171.400 149.400 172.000 ;
        RECT 59.800 170.800 60.600 171.000 ;
        RECT 181.000 170.800 181.800 171.000 ;
        RECT 59.800 170.200 86.800 170.800 ;
        RECT 154.800 170.200 181.800 170.800 ;
        RECT 205.400 170.800 206.200 171.000 ;
        RECT 298.200 170.800 299.000 171.000 ;
        RECT 393.800 170.800 394.600 171.000 ;
        RECT 205.400 170.200 232.400 170.800 ;
        RECT 298.200 170.200 325.200 170.800 ;
        RECT 367.600 170.200 394.600 170.800 ;
        RECT 421.400 170.800 422.200 171.000 ;
        RECT 517.400 170.800 518.200 171.000 ;
        RECT 421.400 170.200 448.400 170.800 ;
        RECT 517.400 170.200 544.400 170.800 ;
        RECT 1.200 161.600 2.000 166.200 ;
        RECT 7.600 161.600 8.400 170.200 ;
        RECT 9.200 161.600 10.000 170.200 ;
        RECT 17.200 161.600 18.000 170.200 ;
        RECT 18.800 161.600 19.600 166.200 ;
        RECT 23.600 161.600 24.400 166.200 ;
        RECT 26.800 161.600 27.600 165.800 ;
        RECT 30.000 161.600 30.800 166.200 ;
        RECT 31.600 161.600 32.400 166.200 ;
        RECT 34.800 161.600 35.600 165.800 ;
        RECT 38.000 161.600 38.800 170.200 ;
        RECT 44.400 161.600 45.200 170.200 ;
        RECT 82.600 170.000 83.600 170.200 ;
        RECT 86.000 169.600 86.800 170.200 ;
        RECT 46.000 161.600 46.800 166.200 ;
        RECT 49.200 161.600 50.000 166.200 ;
        RECT 50.800 161.600 51.600 166.200 ;
        RECT 54.000 161.600 54.800 166.200 ;
        RECT 55.600 161.600 56.400 166.200 ;
        RECT 58.800 161.600 59.600 166.200 ;
        RECT 62.000 161.600 62.800 166.200 ;
        RECT 65.200 161.600 66.000 166.200 ;
        RECT 73.200 161.600 74.000 166.200 ;
        RECT 76.400 161.600 77.200 166.200 ;
        RECT 82.800 161.600 83.600 166.200 ;
        RECT 86.000 161.600 86.800 166.200 ;
        RECT 89.200 161.600 90.000 166.200 ;
        RECT 90.800 161.600 91.600 170.200 ;
        RECT 95.000 161.600 95.800 166.200 ;
        RECT 100.400 161.600 101.200 170.200 ;
        RECT 154.800 169.600 155.600 170.200 ;
        RECT 158.200 170.000 159.000 170.200 ;
        RECT 228.200 170.000 229.000 170.200 ;
        RECT 231.600 169.600 232.400 170.200 ;
        RECT 106.800 161.600 107.600 169.000 ;
        RECT 116.400 161.600 117.200 166.200 ;
        RECT 119.600 161.600 120.400 166.200 ;
        RECT 122.800 161.600 123.600 166.200 ;
        RECT 126.000 161.600 126.800 166.200 ;
        RECT 134.000 161.600 134.800 166.200 ;
        RECT 137.200 161.600 138.000 166.200 ;
        RECT 143.600 161.600 144.400 166.200 ;
        RECT 146.800 161.600 147.600 166.200 ;
        RECT 150.000 161.600 150.800 166.200 ;
        RECT 151.600 161.600 152.400 166.200 ;
        RECT 154.800 161.600 155.600 166.200 ;
        RECT 158.000 161.600 158.800 166.200 ;
        RECT 164.400 161.600 165.200 166.200 ;
        RECT 167.600 161.600 168.400 166.200 ;
        RECT 175.600 161.600 176.400 166.200 ;
        RECT 178.800 161.600 179.600 166.200 ;
        RECT 182.000 161.600 182.800 166.200 ;
        RECT 185.200 161.600 186.000 166.200 ;
        RECT 186.800 161.600 187.600 166.200 ;
        RECT 190.000 161.600 190.800 166.200 ;
        RECT 194.800 161.600 195.600 169.000 ;
        RECT 199.600 161.600 200.400 166.200 ;
        RECT 201.200 161.600 202.000 166.200 ;
        RECT 204.400 161.600 205.200 166.200 ;
        RECT 207.600 161.600 208.400 166.200 ;
        RECT 210.800 161.600 211.600 166.200 ;
        RECT 218.800 161.600 219.600 166.200 ;
        RECT 222.000 161.600 222.800 166.200 ;
        RECT 228.400 161.600 229.200 166.200 ;
        RECT 231.600 161.600 232.400 166.200 ;
        RECT 234.800 161.600 235.600 166.200 ;
        RECT 239.600 161.600 240.400 169.000 ;
        RECT 244.400 161.600 245.200 166.200 ;
        RECT 246.600 161.600 247.400 166.200 ;
        RECT 250.800 161.600 251.600 170.200 ;
        RECT 252.400 161.600 253.200 166.200 ;
        RECT 255.600 161.600 256.400 166.200 ;
        RECT 260.400 161.600 261.200 169.000 ;
        RECT 265.200 161.600 266.000 165.800 ;
        RECT 268.400 161.600 269.200 166.200 ;
        RECT 273.200 161.600 274.000 169.000 ;
        RECT 282.800 161.600 283.600 170.200 ;
        RECT 287.000 161.600 287.800 166.200 ;
        RECT 289.200 161.600 290.000 170.200 ;
        RECT 321.000 170.000 321.800 170.200 ;
        RECT 324.400 169.600 325.200 170.200 ;
        RECT 294.000 161.600 294.800 166.200 ;
        RECT 297.200 161.600 298.000 166.200 ;
        RECT 300.400 161.600 301.200 166.200 ;
        RECT 303.600 161.600 304.400 166.200 ;
        RECT 311.600 161.600 312.400 166.200 ;
        RECT 314.800 161.600 315.600 166.200 ;
        RECT 321.200 161.600 322.000 166.200 ;
        RECT 324.400 161.600 325.200 166.200 ;
        RECT 327.600 161.600 328.400 166.200 ;
        RECT 329.200 161.600 330.000 166.200 ;
        RECT 332.400 161.600 333.200 166.200 ;
        RECT 334.000 161.600 334.800 166.200 ;
        RECT 337.200 161.600 338.000 170.200 ;
        RECT 341.400 161.600 342.200 166.200 ;
        RECT 344.200 161.600 345.000 166.200 ;
        RECT 348.400 161.600 349.200 170.200 ;
        RECT 351.600 161.600 352.400 169.000 ;
        RECT 356.400 161.600 357.200 166.200 ;
        RECT 358.000 161.600 358.800 170.200 ;
        RECT 367.600 169.600 368.400 170.200 ;
        RECT 370.800 170.000 371.800 170.200 ;
        RECT 362.200 161.600 363.000 166.200 ;
        RECT 364.400 161.600 365.200 166.200 ;
        RECT 367.600 161.600 368.400 166.200 ;
        RECT 370.800 161.600 371.600 166.200 ;
        RECT 377.200 161.600 378.000 166.200 ;
        RECT 380.400 161.600 381.200 166.200 ;
        RECT 388.400 161.600 389.200 166.200 ;
        RECT 391.600 161.600 392.400 166.200 ;
        RECT 394.800 161.600 395.600 166.200 ;
        RECT 398.000 161.600 398.800 166.200 ;
        RECT 401.200 161.600 402.000 165.800 ;
        RECT 404.400 161.600 405.200 166.200 ;
        RECT 409.200 161.600 410.000 170.200 ;
        RECT 444.200 170.000 445.200 170.200 ;
        RECT 447.600 169.600 448.400 170.200 ;
        RECT 417.200 161.600 418.000 166.200 ;
        RECT 420.400 161.600 421.200 166.200 ;
        RECT 423.600 161.600 424.400 166.200 ;
        RECT 426.800 161.600 427.600 166.200 ;
        RECT 434.800 161.600 435.600 166.200 ;
        RECT 438.000 161.600 438.800 166.200 ;
        RECT 444.400 161.600 445.200 166.200 ;
        RECT 447.600 161.600 448.400 166.200 ;
        RECT 450.800 161.600 451.600 166.200 ;
        RECT 455.600 161.600 456.400 170.200 ;
        RECT 457.200 161.600 458.000 170.200 ;
        RECT 460.400 161.600 461.200 170.200 ;
        RECT 465.200 161.600 466.000 170.200 ;
        RECT 468.400 161.600 469.200 165.800 ;
        RECT 471.600 161.600 472.400 166.200 ;
        RECT 474.800 161.600 475.600 165.800 ;
        RECT 478.000 161.600 478.800 166.200 ;
        RECT 481.200 161.600 482.000 170.200 ;
        RECT 482.800 161.600 483.600 166.200 ;
        RECT 486.000 161.600 486.800 165.800 ;
        RECT 490.800 161.600 491.600 166.200 ;
        RECT 494.000 161.600 494.800 165.800 ;
        RECT 497.200 161.600 498.000 166.200 ;
        RECT 498.800 161.600 499.600 170.200 ;
        RECT 540.200 170.000 541.200 170.200 ;
        RECT 543.600 169.600 544.400 170.200 ;
        RECT 505.200 161.600 506.000 169.000 ;
        RECT 508.400 161.600 509.200 166.200 ;
        RECT 511.600 161.600 512.400 166.200 ;
        RECT 513.200 161.600 514.000 166.200 ;
        RECT 516.400 161.600 517.200 166.200 ;
        RECT 519.600 161.600 520.400 166.200 ;
        RECT 522.800 161.600 523.600 166.200 ;
        RECT 530.800 161.600 531.600 166.200 ;
        RECT 534.000 161.600 534.800 166.200 ;
        RECT 540.400 161.600 541.200 166.200 ;
        RECT 543.600 161.600 544.400 166.200 ;
        RECT 546.800 161.600 547.600 166.200 ;
        RECT 0.400 160.400 551.600 161.600 ;
        RECT 2.800 153.000 3.600 160.400 ;
        RECT 6.000 155.800 6.800 160.400 ;
        RECT 9.200 156.200 10.000 160.400 ;
        RECT 22.000 153.800 22.800 160.400 ;
        RECT 25.200 155.800 26.000 160.400 ;
        RECT 28.400 151.800 29.200 160.400 ;
        RECT 33.200 151.800 34.000 160.400 ;
        RECT 39.600 155.800 40.400 160.400 ;
        RECT 41.200 155.800 42.000 160.400 ;
        RECT 44.400 155.800 45.200 160.400 ;
        RECT 47.600 153.800 48.400 160.400 ;
        RECT 58.800 151.800 59.600 160.400 ;
        RECT 63.000 155.800 63.800 160.400 ;
        RECT 65.200 155.800 66.000 160.400 ;
        RECT 68.400 155.800 69.200 160.400 ;
        RECT 70.000 155.800 70.800 160.400 ;
        RECT 73.200 155.800 74.000 160.400 ;
        RECT 76.400 155.800 77.200 160.400 ;
        RECT 79.600 155.800 80.400 160.400 ;
        RECT 87.600 155.800 88.400 160.400 ;
        RECT 90.800 155.800 91.600 160.400 ;
        RECT 97.200 155.800 98.000 160.400 ;
        RECT 100.400 155.800 101.200 160.400 ;
        RECT 103.600 155.800 104.400 160.400 ;
        RECT 97.000 151.800 98.000 152.000 ;
        RECT 100.400 151.800 101.200 152.400 ;
        RECT 108.400 151.800 109.200 160.400 ;
        RECT 110.000 151.800 110.800 160.400 ;
        RECT 113.200 151.800 114.000 160.400 ;
        RECT 117.400 155.800 118.200 160.400 ;
        RECT 119.600 155.800 120.400 160.400 ;
        RECT 130.800 152.000 131.600 160.400 ;
        RECT 136.400 155.800 137.200 160.400 ;
        RECT 139.600 155.800 140.400 160.400 ;
        RECT 145.200 151.800 146.000 160.400 ;
        RECT 148.400 155.800 149.200 160.400 ;
        RECT 151.600 155.800 152.400 160.400 ;
        RECT 154.800 155.800 155.600 160.400 ;
        RECT 161.200 155.800 162.000 160.400 ;
        RECT 164.400 155.800 165.200 160.400 ;
        RECT 172.400 155.800 173.200 160.400 ;
        RECT 175.600 155.800 176.400 160.400 ;
        RECT 178.800 155.800 179.600 160.400 ;
        RECT 182.000 155.800 182.800 160.400 ;
        RECT 151.600 151.800 152.400 152.400 ;
        RECT 155.000 151.800 155.800 152.000 ;
        RECT 183.600 151.800 184.400 160.400 ;
        RECT 187.800 155.800 188.600 160.400 ;
        RECT 190.000 155.800 190.800 160.400 ;
        RECT 193.200 155.800 194.000 160.400 ;
        RECT 198.000 153.000 198.800 160.400 ;
        RECT 201.200 155.800 202.000 160.400 ;
        RECT 207.600 151.800 208.400 160.400 ;
        RECT 209.200 155.800 210.000 160.400 ;
        RECT 212.400 152.200 213.200 160.400 ;
        RECT 215.600 151.800 216.400 160.400 ;
        RECT 219.800 155.800 220.600 160.400 ;
        RECT 222.000 155.800 222.800 160.400 ;
        RECT 225.200 155.800 226.000 160.400 ;
        RECT 228.400 155.800 229.200 160.400 ;
        RECT 234.800 155.800 235.600 160.400 ;
        RECT 238.000 155.800 238.800 160.400 ;
        RECT 246.000 155.800 246.800 160.400 ;
        RECT 249.200 155.800 250.000 160.400 ;
        RECT 252.400 155.800 253.200 160.400 ;
        RECT 255.600 155.800 256.400 160.400 ;
        RECT 257.200 155.800 258.000 160.400 ;
        RECT 260.400 155.800 261.200 160.400 ;
        RECT 265.200 153.000 266.000 160.400 ;
        RECT 268.400 155.800 269.200 160.400 ;
        RECT 271.600 156.200 272.400 160.400 ;
        RECT 281.200 155.800 282.000 160.400 ;
        RECT 225.200 151.800 226.000 152.400 ;
        RECT 284.400 152.200 285.200 160.400 ;
        RECT 288.200 155.800 289.000 160.400 ;
        RECT 228.400 151.800 229.400 152.000 ;
        RECT 292.400 151.800 293.200 160.400 ;
        RECT 294.000 155.800 294.800 160.400 ;
        RECT 297.200 155.800 298.000 160.400 ;
        RECT 300.400 155.800 301.200 160.400 ;
        RECT 303.600 155.800 304.400 160.400 ;
        RECT 311.600 155.800 312.400 160.400 ;
        RECT 314.800 155.600 315.600 160.400 ;
        RECT 321.200 155.800 322.000 160.400 ;
        RECT 324.400 155.800 325.200 160.400 ;
        RECT 327.600 155.800 328.400 160.400 ;
        RECT 329.800 155.800 330.600 160.400 ;
        RECT 334.000 151.800 334.800 160.400 ;
        RECT 337.200 155.800 338.000 160.400 ;
        RECT 339.400 155.800 340.200 160.400 ;
        RECT 343.600 151.800 344.400 160.400 ;
        RECT 345.800 155.800 346.600 160.400 ;
        RECT 350.000 151.800 350.800 160.400 ;
        RECT 352.200 155.800 353.000 160.400 ;
        RECT 356.400 151.800 357.200 160.400 ;
        RECT 358.000 151.800 358.800 160.400 ;
        RECT 362.200 155.800 363.000 160.400 ;
        RECT 364.400 155.800 365.200 160.400 ;
        RECT 367.600 155.800 368.400 160.400 ;
        RECT 374.000 153.000 374.800 160.400 ;
        RECT 378.400 151.800 379.200 160.400 ;
        RECT 383.600 152.200 384.400 160.400 ;
        RECT 388.400 155.800 389.200 160.400 ;
        RECT 391.600 152.200 392.400 160.400 ;
        RECT 394.800 155.800 395.600 160.400 ;
        RECT 398.000 156.200 398.800 160.400 ;
        RECT 401.200 155.800 402.000 160.400 ;
        RECT 404.400 156.200 405.200 160.400 ;
        RECT 407.600 155.800 408.400 160.400 ;
        RECT 409.800 155.800 410.600 160.400 ;
        RECT 414.000 151.800 414.800 160.400 ;
        RECT 415.600 155.800 416.400 160.400 ;
        RECT 420.400 152.200 421.200 160.400 ;
        RECT 425.600 151.800 426.400 160.400 ;
        RECT 436.400 152.000 437.200 160.400 ;
        RECT 442.000 155.800 442.800 160.400 ;
        RECT 445.200 155.800 446.000 160.400 ;
        RECT 450.800 151.800 451.600 160.400 ;
        RECT 455.600 156.200 456.400 160.400 ;
        RECT 458.800 155.800 459.600 160.400 ;
        RECT 460.400 155.800 461.200 160.400 ;
        RECT 463.600 156.200 464.400 160.400 ;
        RECT 468.400 153.800 469.200 160.400 ;
        RECT 480.800 151.800 481.600 160.400 ;
        RECT 486.000 152.200 486.800 160.400 ;
        RECT 490.800 155.800 491.600 160.400 ;
        RECT 492.400 151.800 493.200 160.400 ;
        RECT 498.800 151.800 499.600 160.400 ;
        RECT 501.600 151.800 502.400 160.400 ;
        RECT 506.800 152.200 507.600 160.400 ;
        RECT 511.600 155.800 512.400 160.400 ;
        RECT 514.800 155.800 515.600 160.400 ;
        RECT 518.000 152.200 518.800 160.400 ;
        RECT 523.200 151.800 524.000 160.400 ;
        RECT 527.600 152.000 528.400 160.400 ;
        RECT 533.200 155.800 534.000 160.400 ;
        RECT 536.400 155.800 537.200 160.400 ;
        RECT 542.000 151.800 542.800 160.400 ;
        RECT 546.800 153.000 547.600 160.400 ;
        RECT 74.200 151.200 101.200 151.800 ;
        RECT 151.600 151.200 178.600 151.800 ;
        RECT 225.200 151.200 252.200 151.800 ;
        RECT 74.200 151.000 75.000 151.200 ;
        RECT 177.800 151.000 178.600 151.200 ;
        RECT 251.400 151.000 252.200 151.200 ;
        RECT 303.600 150.000 327.000 150.600 ;
        RECT 303.600 149.400 304.400 150.000 ;
        RECT 314.800 149.600 315.600 150.000 ;
        RECT 321.200 149.600 322.000 150.000 ;
        RECT 326.200 149.800 327.000 150.000 ;
        RECT 281.200 132.000 282.000 132.600 ;
        RECT 298.800 132.000 299.600 132.400 ;
        RECT 303.800 132.000 304.600 132.200 ;
        RECT 281.200 131.400 304.600 132.000 ;
        RECT 53.400 130.800 54.200 131.000 ;
        RECT 128.200 130.800 129.000 131.000 ;
        RECT 53.400 130.200 80.400 130.800 ;
        RECT 102.000 130.200 129.000 130.800 ;
        RECT 186.200 130.800 187.000 131.000 ;
        RECT 352.200 130.800 353.000 131.000 ;
        RECT 186.200 130.200 213.200 130.800 ;
        RECT 326.000 130.200 353.000 130.800 ;
        RECT 399.000 130.800 399.800 131.000 ;
        RECT 494.600 130.800 495.400 131.000 ;
        RECT 399.000 130.200 426.000 130.800 ;
        RECT 468.400 130.200 495.400 130.800 ;
        RECT 519.000 130.800 519.800 131.000 ;
        RECT 519.000 130.200 546.000 130.800 ;
        RECT 2.800 121.600 3.600 130.200 ;
        RECT 4.400 121.600 5.200 126.200 ;
        RECT 7.600 121.600 8.400 126.200 ;
        RECT 10.800 121.600 11.600 126.200 ;
        RECT 12.400 121.600 13.200 130.200 ;
        RECT 17.200 121.600 18.000 130.200 ;
        RECT 21.400 121.600 22.200 126.200 ;
        RECT 25.200 121.600 26.000 125.800 ;
        RECT 28.400 121.600 29.200 126.200 ;
        RECT 31.600 121.600 32.400 125.800 ;
        RECT 34.800 121.600 35.600 126.200 ;
        RECT 36.400 121.600 37.200 130.200 ;
        RECT 76.200 130.000 77.200 130.200 ;
        RECT 79.600 129.600 80.400 130.200 ;
        RECT 40.600 121.600 41.400 126.200 ;
        RECT 44.400 121.600 45.200 125.800 ;
        RECT 47.600 121.600 48.400 126.200 ;
        RECT 49.200 121.600 50.000 126.200 ;
        RECT 52.400 121.600 53.200 126.200 ;
        RECT 55.600 121.600 56.400 126.200 ;
        RECT 58.800 121.600 59.600 126.200 ;
        RECT 66.800 121.600 67.600 126.200 ;
        RECT 70.000 121.600 70.800 126.200 ;
        RECT 76.400 121.600 77.200 126.200 ;
        RECT 79.600 121.600 80.400 126.200 ;
        RECT 82.800 121.600 83.600 126.200 ;
        RECT 84.400 121.600 85.200 130.200 ;
        RECT 90.800 121.600 91.600 130.200 ;
        RECT 102.000 129.600 102.800 130.200 ;
        RECT 105.200 130.000 106.200 130.200 ;
        RECT 94.000 121.600 94.800 129.000 ;
        RECT 98.800 121.600 99.600 126.200 ;
        RECT 102.000 121.600 102.800 126.200 ;
        RECT 105.200 121.600 106.000 126.200 ;
        RECT 111.600 121.600 112.400 126.200 ;
        RECT 114.800 121.600 115.600 126.200 ;
        RECT 122.800 121.600 123.600 126.200 ;
        RECT 126.000 121.600 126.800 126.200 ;
        RECT 129.200 121.600 130.000 126.200 ;
        RECT 132.400 121.600 133.200 126.200 ;
        RECT 142.000 121.600 142.800 126.200 ;
        RECT 143.600 121.600 144.400 130.200 ;
        RECT 147.800 121.600 148.600 126.200 ;
        RECT 150.000 121.600 150.800 126.200 ;
        RECT 153.200 121.600 154.000 129.800 ;
        RECT 158.000 121.600 158.800 129.800 ;
        RECT 161.200 121.600 162.000 126.200 ;
        RECT 166.000 121.600 166.800 130.200 ;
        RECT 167.600 121.600 168.400 130.200 ;
        RECT 209.000 130.000 209.800 130.200 ;
        RECT 212.400 129.600 213.200 130.200 ;
        RECT 171.800 121.600 172.600 126.200 ;
        RECT 174.000 121.600 174.800 126.200 ;
        RECT 177.200 121.600 178.000 126.200 ;
        RECT 180.400 121.600 181.200 126.200 ;
        RECT 182.000 121.600 182.800 126.200 ;
        RECT 185.200 121.600 186.000 126.200 ;
        RECT 188.400 121.600 189.200 126.200 ;
        RECT 191.600 121.600 192.400 126.200 ;
        RECT 199.600 121.600 200.400 126.200 ;
        RECT 202.800 121.600 203.600 126.200 ;
        RECT 209.200 121.600 210.000 126.200 ;
        RECT 212.400 121.600 213.200 126.200 ;
        RECT 215.600 121.600 216.400 126.200 ;
        RECT 217.200 121.600 218.000 130.200 ;
        RECT 222.600 121.600 223.400 126.200 ;
        RECT 226.800 121.600 227.600 130.200 ;
        RECT 228.400 121.600 229.200 130.200 ;
        RECT 232.600 121.600 233.400 126.200 ;
        RECT 236.400 121.600 237.200 125.800 ;
        RECT 239.600 121.600 240.400 126.200 ;
        RECT 242.800 121.600 243.600 126.200 ;
        RECT 244.400 121.600 245.200 126.200 ;
        RECT 247.600 121.600 248.400 126.200 ;
        RECT 252.400 121.600 253.200 130.200 ;
        RECT 254.000 121.600 254.800 130.200 ;
        RECT 258.800 121.600 259.600 130.200 ;
        RECT 263.000 121.600 263.800 126.200 ;
        RECT 271.600 121.600 272.400 126.200 ;
        RECT 274.800 121.600 275.600 126.200 ;
        RECT 278.000 121.600 278.800 126.200 ;
        RECT 281.200 121.600 282.000 126.200 ;
        RECT 289.200 121.600 290.000 126.200 ;
        RECT 292.400 121.600 293.200 126.200 ;
        RECT 298.800 121.600 299.600 126.200 ;
        RECT 302.000 121.600 302.800 126.200 ;
        RECT 305.200 121.600 306.000 126.200 ;
        RECT 307.400 121.600 308.200 126.200 ;
        RECT 311.600 121.600 312.400 130.200 ;
        RECT 314.800 121.600 315.600 126.200 ;
        RECT 317.000 121.600 317.800 126.200 ;
        RECT 321.200 121.600 322.000 130.200 ;
        RECT 326.000 129.600 326.800 130.200 ;
        RECT 329.200 130.000 330.200 130.200 ;
        RECT 322.800 121.600 323.600 126.200 ;
        RECT 326.000 121.600 326.800 126.200 ;
        RECT 329.200 121.600 330.000 126.200 ;
        RECT 335.600 121.600 336.400 126.200 ;
        RECT 338.800 121.600 339.600 126.200 ;
        RECT 346.800 121.600 347.600 126.200 ;
        RECT 350.000 121.600 350.800 126.200 ;
        RECT 353.200 121.600 354.000 126.200 ;
        RECT 356.400 121.600 357.200 126.200 ;
        RECT 358.000 121.600 358.800 126.200 ;
        RECT 361.200 121.600 362.000 126.200 ;
        RECT 364.400 121.600 365.200 130.200 ;
        RECT 370.800 121.600 371.600 130.200 ;
        RECT 374.000 121.600 374.800 129.000 ;
        RECT 378.800 121.600 379.600 130.200 ;
        RECT 421.800 130.000 422.800 130.200 ;
        RECT 425.200 129.600 426.000 130.200 ;
        RECT 385.200 121.600 386.000 129.000 ;
        RECT 393.200 121.600 394.000 126.200 ;
        RECT 394.800 121.600 395.600 126.200 ;
        RECT 398.000 121.600 398.800 126.200 ;
        RECT 401.200 121.600 402.000 126.200 ;
        RECT 404.400 121.600 405.200 126.200 ;
        RECT 412.400 121.600 413.200 126.200 ;
        RECT 415.600 121.600 416.400 126.200 ;
        RECT 422.000 121.600 422.800 126.200 ;
        RECT 425.200 121.600 426.000 126.200 ;
        RECT 428.400 121.600 429.200 126.200 ;
        RECT 436.400 121.600 437.200 130.200 ;
        RECT 442.800 121.600 443.600 129.000 ;
        RECT 447.600 121.600 448.400 126.200 ;
        RECT 450.800 121.600 451.600 125.800 ;
        RECT 454.000 121.600 454.800 130.200 ;
        RECT 460.400 121.600 461.200 130.200 ;
        RECT 468.400 129.600 469.200 130.200 ;
        RECT 471.800 130.000 472.600 130.200 ;
        RECT 463.600 121.600 464.400 126.200 ;
        RECT 465.200 121.600 466.000 126.200 ;
        RECT 468.400 121.600 469.200 126.200 ;
        RECT 471.600 121.600 472.400 126.200 ;
        RECT 478.000 121.600 478.800 126.200 ;
        RECT 481.200 121.600 482.000 126.200 ;
        RECT 489.200 121.600 490.000 126.200 ;
        RECT 492.400 121.600 493.200 126.200 ;
        RECT 495.600 121.600 496.400 126.200 ;
        RECT 498.800 121.600 499.600 126.200 ;
        RECT 502.000 121.600 502.800 129.800 ;
        RECT 507.200 121.600 508.000 130.200 ;
        RECT 541.800 130.000 542.600 130.200 ;
        RECT 545.200 129.600 546.000 130.200 ;
        RECT 510.000 121.600 510.800 126.200 ;
        RECT 513.200 121.600 514.000 126.200 ;
        RECT 514.800 121.600 515.600 126.200 ;
        RECT 518.000 121.600 518.800 126.200 ;
        RECT 521.200 121.600 522.000 126.200 ;
        RECT 524.400 121.600 525.200 126.200 ;
        RECT 532.400 121.600 533.200 126.200 ;
        RECT 535.600 121.600 536.400 126.200 ;
        RECT 542.000 121.600 542.800 126.200 ;
        RECT 545.200 121.600 546.000 126.200 ;
        RECT 548.400 121.600 549.200 126.200 ;
        RECT 0.400 120.400 551.600 121.600 ;
        RECT 2.800 116.200 3.600 120.400 ;
        RECT 6.000 115.800 6.800 120.400 ;
        RECT 7.600 115.800 8.400 120.400 ;
        RECT 10.800 115.800 11.600 120.400 ;
        RECT 14.000 116.200 14.800 120.400 ;
        RECT 17.200 115.800 18.000 120.400 ;
        RECT 20.400 116.200 21.200 120.400 ;
        RECT 23.600 115.800 24.400 120.400 ;
        RECT 25.200 115.800 26.000 120.400 ;
        RECT 28.400 116.200 29.200 120.400 ;
        RECT 32.200 115.800 33.000 120.400 ;
        RECT 36.400 111.800 37.200 120.400 ;
        RECT 38.000 111.800 38.800 120.400 ;
        RECT 41.200 111.800 42.000 120.400 ;
        RECT 42.800 115.800 43.600 120.400 ;
        RECT 46.000 115.800 46.800 120.400 ;
        RECT 49.200 115.800 50.000 120.400 ;
        RECT 52.400 115.800 53.200 120.400 ;
        RECT 60.400 115.800 61.200 120.400 ;
        RECT 63.600 115.800 64.400 120.400 ;
        RECT 70.000 115.800 70.800 120.400 ;
        RECT 73.200 115.800 74.000 120.400 ;
        RECT 76.400 115.800 77.200 120.400 ;
        RECT 69.800 111.800 70.600 112.000 ;
        RECT 73.200 111.800 74.000 112.400 ;
        RECT 78.000 111.800 78.800 120.400 ;
        RECT 82.200 115.800 83.000 120.400 ;
        RECT 84.400 115.800 85.200 120.400 ;
        RECT 87.600 115.800 88.400 120.400 ;
        RECT 90.800 115.800 91.600 120.400 ;
        RECT 97.200 115.800 98.000 120.400 ;
        RECT 100.400 115.800 101.200 120.400 ;
        RECT 108.400 115.800 109.200 120.400 ;
        RECT 111.600 115.800 112.400 120.400 ;
        RECT 114.800 115.800 115.600 120.400 ;
        RECT 118.000 115.800 118.800 120.400 ;
        RECT 121.200 115.800 122.000 120.400 ;
        RECT 87.600 111.800 88.400 112.400 ;
        RECT 91.000 111.800 91.800 112.000 ;
        RECT 132.400 111.800 133.200 120.400 ;
        RECT 137.200 113.000 138.000 120.400 ;
        RECT 140.400 115.800 141.200 120.400 ;
        RECT 146.800 111.800 147.600 120.400 ;
        RECT 148.400 111.800 149.200 120.400 ;
        RECT 152.600 115.800 153.400 120.400 ;
        RECT 156.400 113.000 157.200 120.400 ;
        RECT 161.200 111.800 162.000 120.400 ;
        RECT 166.000 111.800 166.800 120.400 ;
        RECT 170.200 115.800 171.000 120.400 ;
        RECT 174.000 115.800 174.800 120.400 ;
        RECT 175.600 115.800 176.400 120.400 ;
        RECT 178.800 115.800 179.600 120.400 ;
        RECT 180.400 115.800 181.200 120.400 ;
        RECT 183.600 115.800 184.400 120.400 ;
        RECT 186.800 115.800 187.600 120.400 ;
        RECT 193.200 115.800 194.000 120.400 ;
        RECT 196.400 115.800 197.200 120.400 ;
        RECT 204.400 115.800 205.200 120.400 ;
        RECT 207.600 115.800 208.400 120.400 ;
        RECT 210.800 115.800 211.600 120.400 ;
        RECT 214.000 115.800 214.800 120.400 ;
        RECT 218.800 113.000 219.600 120.400 ;
        RECT 222.000 115.800 222.800 120.400 ;
        RECT 225.200 115.800 226.000 120.400 ;
        RECT 227.400 115.800 228.200 120.400 ;
        RECT 183.600 111.800 184.400 112.400 ;
        RECT 187.000 111.800 187.800 112.000 ;
        RECT 231.600 111.800 232.400 120.400 ;
        RECT 233.200 111.800 234.000 120.400 ;
        RECT 239.600 115.800 240.400 120.400 ;
        RECT 243.800 111.800 244.600 120.400 ;
        RECT 248.200 115.800 249.000 120.400 ;
        RECT 252.400 111.800 253.200 120.400 ;
        RECT 254.000 111.800 254.800 120.400 ;
        RECT 258.200 115.800 259.000 120.400 ;
        RECT 262.000 113.000 262.800 120.400 ;
        RECT 273.200 115.800 274.000 120.400 ;
        RECT 276.400 115.800 277.200 120.400 ;
        RECT 279.600 115.800 280.400 120.400 ;
        RECT 282.800 115.800 283.600 120.400 ;
        RECT 290.800 115.800 291.600 120.400 ;
        RECT 294.000 115.600 294.800 120.400 ;
        RECT 300.400 115.800 301.200 120.400 ;
        RECT 303.600 115.800 304.400 120.400 ;
        RECT 306.800 115.800 307.600 120.400 ;
        RECT 308.400 111.800 309.200 120.400 ;
        RECT 312.600 115.800 313.400 120.400 ;
        RECT 315.400 115.800 316.200 120.400 ;
        RECT 319.600 111.800 320.400 120.400 ;
        RECT 321.200 115.800 322.000 120.400 ;
        RECT 324.400 111.800 325.200 120.400 ;
        RECT 327.600 111.800 328.400 120.400 ;
        RECT 330.800 111.800 331.600 120.400 ;
        RECT 334.000 111.800 334.800 120.400 ;
        RECT 337.200 111.800 338.000 120.400 ;
        RECT 338.800 115.800 339.600 120.400 ;
        RECT 342.000 115.800 342.800 120.400 ;
        RECT 345.200 115.800 346.000 120.400 ;
        RECT 351.600 115.800 352.400 120.400 ;
        RECT 354.800 115.800 355.600 120.400 ;
        RECT 362.800 115.800 363.600 120.400 ;
        RECT 366.000 115.800 366.800 120.400 ;
        RECT 369.200 115.800 370.000 120.400 ;
        RECT 372.400 115.800 373.200 120.400 ;
        RECT 342.000 111.800 342.800 112.400 ;
        RECT 345.400 111.800 346.200 112.000 ;
        RECT 374.000 111.800 374.800 120.400 ;
        RECT 380.400 111.800 381.200 120.400 ;
        RECT 383.600 115.800 384.400 120.400 ;
        RECT 386.800 113.000 387.600 120.400 ;
        RECT 396.400 111.800 397.200 120.400 ;
        RECT 398.000 115.800 398.800 120.400 ;
        RECT 404.400 111.800 405.200 120.400 ;
        RECT 406.000 111.800 406.800 120.400 ;
        RECT 412.400 111.800 413.200 120.400 ;
        RECT 414.600 115.800 415.400 120.400 ;
        RECT 418.800 111.800 419.600 120.400 ;
        RECT 423.600 111.800 424.400 120.400 ;
        RECT 431.600 111.800 432.400 120.400 ;
        RECT 438.000 111.800 438.800 120.400 ;
        RECT 439.600 115.800 440.400 120.400 ;
        RECT 442.800 116.200 443.600 120.400 ;
        RECT 447.600 113.000 448.400 120.400 ;
        RECT 452.400 115.800 453.200 120.400 ;
        RECT 455.600 115.800 456.400 120.400 ;
        RECT 457.200 111.800 458.000 120.400 ;
        RECT 461.400 115.800 462.200 120.400 ;
        RECT 463.600 111.800 464.400 120.400 ;
        RECT 468.400 115.800 469.200 120.400 ;
        RECT 471.600 115.800 472.400 120.400 ;
        RECT 473.200 111.800 474.000 120.400 ;
        RECT 478.000 113.000 478.800 120.400 ;
        RECT 486.000 112.200 486.800 120.400 ;
        RECT 491.200 111.800 492.000 120.400 ;
        RECT 494.000 115.800 494.800 120.400 ;
        RECT 497.200 115.800 498.000 120.400 ;
        RECT 498.800 111.800 499.600 120.400 ;
        RECT 503.000 115.800 503.800 120.400 ;
        RECT 505.200 115.800 506.000 120.400 ;
        RECT 508.400 115.800 509.200 120.400 ;
        RECT 510.600 115.800 511.400 120.400 ;
        RECT 514.800 111.800 515.600 120.400 ;
        RECT 516.400 115.800 517.200 120.400 ;
        RECT 519.600 115.800 520.400 120.400 ;
        RECT 522.800 115.800 523.600 120.400 ;
        RECT 526.000 115.800 526.800 120.400 ;
        RECT 534.000 115.800 534.800 120.400 ;
        RECT 537.200 115.800 538.000 120.400 ;
        RECT 543.600 115.800 544.400 120.400 ;
        RECT 546.800 115.800 547.600 120.400 ;
        RECT 550.000 115.800 550.800 120.400 ;
        RECT 543.400 111.800 544.200 112.000 ;
        RECT 546.800 111.800 547.600 112.400 ;
        RECT 47.000 111.200 74.000 111.800 ;
        RECT 87.600 111.200 114.600 111.800 ;
        RECT 183.600 111.200 210.600 111.800 ;
        RECT 342.000 111.200 369.000 111.800 ;
        RECT 47.000 111.000 47.800 111.200 ;
        RECT 113.800 111.000 114.600 111.200 ;
        RECT 209.800 111.000 210.600 111.200 ;
        RECT 368.200 111.000 369.000 111.200 ;
        RECT 520.600 111.200 547.600 111.800 ;
        RECT 520.600 111.000 521.400 111.200 ;
        RECT 282.800 110.000 306.200 110.600 ;
        RECT 282.800 109.400 283.600 110.000 ;
        RECT 294.000 109.600 294.800 110.000 ;
        RECT 300.400 109.600 301.200 110.000 ;
        RECT 305.400 109.800 306.200 110.000 ;
        RECT 47.400 92.000 48.200 92.200 ;
        RECT 52.400 92.000 53.200 92.400 ;
        RECT 70.000 92.000 70.800 92.600 ;
        RECT 47.400 91.400 70.800 92.000 ;
        RECT 316.400 92.000 317.200 92.600 ;
        RECT 334.000 92.000 334.800 92.400 ;
        RECT 339.000 92.000 339.800 92.200 ;
        RECT 316.400 91.400 339.800 92.000 ;
        RECT 128.200 90.800 129.000 91.000 ;
        RECT 102.000 90.200 129.000 90.800 ;
        RECT 272.600 90.800 273.400 91.000 ;
        RECT 384.200 90.800 385.000 91.000 ;
        RECT 272.600 90.200 299.600 90.800 ;
        RECT 358.000 90.200 385.000 90.800 ;
        RECT 485.400 90.800 486.200 91.000 ;
        RECT 520.600 90.800 521.400 91.000 ;
        RECT 485.400 90.200 512.400 90.800 ;
        RECT 520.600 90.200 547.600 90.800 ;
        RECT 1.200 81.600 2.000 86.200 ;
        RECT 4.400 81.600 5.200 86.200 ;
        RECT 9.200 81.600 10.000 90.200 ;
        RECT 12.400 81.600 13.200 85.800 ;
        RECT 15.600 81.600 16.400 86.200 ;
        RECT 18.800 81.600 19.600 85.800 ;
        RECT 22.000 81.600 22.800 86.200 ;
        RECT 23.600 81.600 24.400 90.200 ;
        RECT 27.800 81.600 28.600 86.200 ;
        RECT 30.000 81.600 30.800 86.200 ;
        RECT 33.200 81.600 34.000 86.200 ;
        RECT 34.800 81.600 35.600 86.200 ;
        RECT 38.000 81.600 38.800 86.200 ;
        RECT 39.600 81.600 40.400 90.200 ;
        RECT 43.800 81.600 44.600 86.200 ;
        RECT 46.000 81.600 46.800 86.200 ;
        RECT 49.200 81.600 50.000 86.200 ;
        RECT 52.400 81.600 53.200 86.200 ;
        RECT 58.800 81.600 59.600 86.200 ;
        RECT 62.000 81.600 62.800 86.200 ;
        RECT 70.000 81.600 70.800 86.200 ;
        RECT 73.200 81.600 74.000 86.200 ;
        RECT 76.400 81.600 77.200 86.200 ;
        RECT 79.600 81.600 80.400 86.200 ;
        RECT 81.800 81.600 82.600 86.200 ;
        RECT 86.000 81.600 86.800 90.200 ;
        RECT 87.600 81.600 88.400 90.200 ;
        RECT 102.000 89.600 102.800 90.200 ;
        RECT 105.200 90.000 106.200 90.200 ;
        RECT 95.600 81.600 96.400 89.000 ;
        RECT 98.800 81.600 99.600 86.200 ;
        RECT 102.000 81.600 102.800 86.200 ;
        RECT 105.200 81.600 106.000 86.200 ;
        RECT 111.600 81.600 112.400 86.200 ;
        RECT 114.800 81.600 115.600 86.200 ;
        RECT 122.800 81.600 123.600 86.200 ;
        RECT 126.000 81.600 126.800 86.200 ;
        RECT 129.200 81.600 130.000 86.200 ;
        RECT 132.400 81.600 133.200 86.200 ;
        RECT 142.000 81.600 142.800 86.200 ;
        RECT 146.200 81.600 147.000 90.200 ;
        RECT 150.600 81.600 151.400 86.200 ;
        RECT 154.800 81.600 155.600 90.200 ;
        RECT 158.000 81.600 158.800 90.000 ;
        RECT 163.600 81.600 164.400 86.200 ;
        RECT 166.800 81.600 167.600 86.200 ;
        RECT 172.400 81.600 173.200 90.200 ;
        RECT 177.200 81.600 178.000 89.000 ;
        RECT 182.000 81.600 182.800 89.000 ;
        RECT 185.200 81.600 186.000 86.200 ;
        RECT 190.000 81.600 190.800 89.000 ;
        RECT 194.800 81.600 195.600 86.200 ;
        RECT 198.000 81.600 198.800 86.200 ;
        RECT 199.600 81.600 200.400 86.200 ;
        RECT 202.800 81.600 203.600 86.200 ;
        RECT 205.000 81.600 205.800 86.200 ;
        RECT 209.200 81.600 210.000 90.200 ;
        RECT 212.400 81.600 213.200 86.200 ;
        RECT 214.000 81.600 214.800 86.200 ;
        RECT 217.200 81.600 218.000 86.200 ;
        RECT 218.800 81.600 219.600 90.200 ;
        RECT 223.600 81.600 224.400 86.200 ;
        RECT 226.800 81.600 227.600 86.200 ;
        RECT 228.400 81.600 229.200 86.200 ;
        RECT 234.800 81.600 235.600 89.000 ;
        RECT 238.000 81.600 238.800 90.200 ;
        RECT 242.200 81.600 243.000 86.200 ;
        RECT 246.000 81.600 246.800 88.200 ;
        RECT 260.400 81.600 261.200 90.200 ;
        RECT 295.400 90.000 296.200 90.200 ;
        RECT 298.800 89.600 299.600 90.200 ;
        RECT 268.400 81.600 269.200 86.200 ;
        RECT 271.600 81.600 272.400 86.200 ;
        RECT 274.800 81.600 275.600 86.200 ;
        RECT 278.000 81.600 278.800 86.200 ;
        RECT 286.000 81.600 286.800 86.200 ;
        RECT 289.200 81.600 290.000 86.200 ;
        RECT 295.600 81.600 296.400 86.200 ;
        RECT 298.800 81.600 299.600 86.200 ;
        RECT 302.000 81.600 302.800 86.200 ;
        RECT 303.600 81.600 304.400 86.200 ;
        RECT 306.800 81.600 307.600 86.200 ;
        RECT 310.000 81.600 310.800 86.200 ;
        RECT 313.200 81.600 314.000 86.200 ;
        RECT 316.400 81.600 317.200 86.200 ;
        RECT 324.400 81.600 325.200 86.200 ;
        RECT 327.600 81.600 328.400 86.200 ;
        RECT 334.000 81.600 334.800 86.200 ;
        RECT 337.200 81.600 338.000 86.200 ;
        RECT 340.400 81.600 341.200 86.200 ;
        RECT 342.000 81.600 342.800 90.200 ;
        RECT 346.200 81.600 347.000 86.200 ;
        RECT 349.000 81.600 349.800 86.200 ;
        RECT 353.200 81.600 354.000 90.200 ;
        RECT 358.000 89.600 358.800 90.200 ;
        RECT 361.200 90.000 362.200 90.200 ;
        RECT 354.800 81.600 355.600 86.200 ;
        RECT 358.000 81.600 358.800 86.200 ;
        RECT 361.200 81.600 362.000 86.200 ;
        RECT 367.600 81.600 368.400 86.200 ;
        RECT 370.800 81.600 371.600 86.200 ;
        RECT 378.800 81.600 379.600 86.200 ;
        RECT 382.000 81.600 382.800 86.200 ;
        RECT 385.200 81.600 386.000 86.200 ;
        RECT 388.400 81.600 389.200 86.200 ;
        RECT 390.000 81.600 390.800 86.200 ;
        RECT 393.200 81.600 394.000 86.200 ;
        RECT 394.800 81.600 395.600 86.200 ;
        RECT 398.000 81.600 398.800 86.200 ;
        RECT 399.600 81.600 400.400 86.200 ;
        RECT 402.800 81.600 403.600 86.200 ;
        RECT 404.400 81.600 405.200 86.200 ;
        RECT 407.600 81.600 408.400 86.200 ;
        RECT 409.800 81.600 410.600 86.200 ;
        RECT 414.000 81.600 414.800 90.200 ;
        RECT 415.600 81.600 416.400 86.200 ;
        RECT 420.400 81.600 421.200 89.000 ;
        RECT 430.000 81.600 430.800 86.200 ;
        RECT 436.400 81.600 437.200 89.000 ;
        RECT 439.600 81.600 440.400 86.200 ;
        RECT 442.800 81.600 443.600 85.800 ;
        RECT 446.000 81.600 446.800 86.200 ;
        RECT 449.200 81.600 450.000 86.200 ;
        RECT 452.400 81.600 453.200 89.000 ;
        RECT 456.800 81.600 457.600 90.200 ;
        RECT 508.200 90.000 509.200 90.200 ;
        RECT 462.000 81.600 462.800 89.800 ;
        RECT 511.600 89.600 512.400 90.200 ;
        RECT 543.400 90.000 544.400 90.200 ;
        RECT 546.800 89.600 547.600 90.200 ;
        RECT 466.800 81.600 467.600 89.000 ;
        RECT 478.000 81.600 478.800 89.000 ;
        RECT 481.200 81.600 482.000 86.200 ;
        RECT 484.400 81.600 485.200 86.200 ;
        RECT 487.600 81.600 488.400 86.200 ;
        RECT 490.800 81.600 491.600 86.200 ;
        RECT 498.800 81.600 499.600 86.200 ;
        RECT 502.000 81.600 502.800 86.200 ;
        RECT 508.400 81.600 509.200 86.200 ;
        RECT 511.600 81.600 512.400 86.200 ;
        RECT 514.800 81.600 515.600 86.200 ;
        RECT 516.400 81.600 517.200 86.200 ;
        RECT 519.600 81.600 520.400 86.200 ;
        RECT 522.800 81.600 523.600 86.200 ;
        RECT 526.000 81.600 526.800 86.200 ;
        RECT 534.000 81.600 534.800 86.200 ;
        RECT 537.200 81.600 538.000 86.200 ;
        RECT 543.600 81.600 544.400 86.200 ;
        RECT 546.800 81.600 547.600 86.200 ;
        RECT 550.000 81.600 550.800 86.200 ;
        RECT 0.400 80.400 551.600 81.600 ;
        RECT 1.200 71.800 2.000 80.400 ;
        RECT 6.000 75.800 6.800 80.400 ;
        RECT 9.200 71.800 10.000 80.400 ;
        RECT 17.200 71.800 18.000 80.400 ;
        RECT 18.800 75.800 19.600 80.400 ;
        RECT 25.200 71.800 26.000 80.400 ;
        RECT 30.000 71.800 30.800 80.400 ;
        RECT 34.800 71.800 35.600 80.400 ;
        RECT 36.400 75.800 37.200 80.400 ;
        RECT 39.600 75.800 40.400 80.400 ;
        RECT 42.800 75.800 43.600 80.400 ;
        RECT 44.400 71.800 45.200 80.400 ;
        RECT 50.800 71.800 51.600 80.400 ;
        RECT 52.400 71.800 53.200 80.400 ;
        RECT 56.600 75.800 57.400 80.400 ;
        RECT 58.800 75.800 59.600 80.400 ;
        RECT 62.000 75.800 62.800 80.400 ;
        RECT 63.600 71.800 64.400 80.400 ;
        RECT 66.800 71.800 67.600 80.400 ;
        RECT 70.000 71.800 70.800 80.400 ;
        RECT 73.200 71.800 74.000 80.400 ;
        RECT 76.400 71.800 77.200 80.400 ;
        RECT 78.000 75.800 78.800 80.400 ;
        RECT 81.200 76.200 82.000 80.400 ;
        RECT 86.000 76.200 86.800 80.400 ;
        RECT 89.200 75.800 90.000 80.400 ;
        RECT 90.800 75.800 91.600 80.400 ;
        RECT 94.000 75.800 94.800 80.400 ;
        RECT 97.200 75.800 98.000 80.400 ;
        RECT 100.400 75.800 101.200 80.400 ;
        RECT 108.400 75.800 109.200 80.400 ;
        RECT 111.600 75.800 112.400 80.400 ;
        RECT 118.000 75.800 118.800 80.400 ;
        RECT 121.200 75.800 122.000 80.400 ;
        RECT 124.400 75.800 125.200 80.400 ;
        RECT 132.400 75.800 133.200 80.400 ;
        RECT 135.600 75.800 136.400 80.400 ;
        RECT 138.800 75.800 139.600 80.400 ;
        RECT 142.000 75.800 142.800 80.400 ;
        RECT 150.000 75.800 150.800 80.400 ;
        RECT 153.200 75.600 154.000 80.400 ;
        RECT 159.600 75.800 160.400 80.400 ;
        RECT 162.800 75.800 163.600 80.400 ;
        RECT 166.000 75.800 166.800 80.400 ;
        RECT 169.200 73.000 170.000 80.400 ;
        RECT 172.400 75.800 173.200 80.400 ;
        RECT 175.600 75.800 176.400 80.400 ;
        RECT 178.800 75.800 179.600 80.400 ;
        RECT 185.200 75.800 186.000 80.400 ;
        RECT 188.400 75.800 189.200 80.400 ;
        RECT 196.400 75.800 197.200 80.400 ;
        RECT 199.600 75.800 200.400 80.400 ;
        RECT 202.800 75.800 203.600 80.400 ;
        RECT 206.000 75.800 206.800 80.400 ;
        RECT 207.600 75.800 208.400 80.400 ;
        RECT 210.800 75.800 211.600 80.400 ;
        RECT 214.000 75.800 214.800 80.400 ;
        RECT 217.200 75.800 218.000 80.400 ;
        RECT 225.200 75.800 226.000 80.400 ;
        RECT 228.400 75.800 229.200 80.400 ;
        RECT 234.800 75.800 235.600 80.400 ;
        RECT 238.000 75.800 238.800 80.400 ;
        RECT 241.200 75.800 242.000 80.400 ;
        RECT 244.400 73.000 245.200 80.400 ;
        RECT 247.600 75.800 248.400 80.400 ;
        RECT 117.800 71.800 118.600 72.000 ;
        RECT 121.200 71.800 122.000 72.400 ;
        RECT 95.000 71.200 122.000 71.800 ;
        RECT 175.600 71.800 176.400 72.400 ;
        RECT 179.000 71.800 179.800 72.000 ;
        RECT 234.600 71.800 235.600 72.000 ;
        RECT 238.000 71.800 238.800 72.400 ;
        RECT 250.800 71.800 251.600 80.400 ;
        RECT 255.000 75.800 255.800 80.400 ;
        RECT 257.800 75.800 258.600 80.400 ;
        RECT 262.000 71.800 262.800 80.400 ;
        RECT 263.600 75.800 264.400 80.400 ;
        RECT 273.200 75.800 274.000 80.400 ;
        RECT 276.400 75.800 277.200 80.400 ;
        RECT 279.600 75.800 280.400 80.400 ;
        RECT 282.800 75.800 283.600 80.400 ;
        RECT 290.800 75.800 291.600 80.400 ;
        RECT 294.000 75.600 294.800 80.400 ;
        RECT 300.400 75.800 301.200 80.400 ;
        RECT 303.600 75.800 304.400 80.400 ;
        RECT 306.800 75.800 307.600 80.400 ;
        RECT 308.400 71.800 309.200 80.400 ;
        RECT 312.600 75.800 313.400 80.400 ;
        RECT 315.400 75.800 316.200 80.400 ;
        RECT 319.600 71.800 320.400 80.400 ;
        RECT 322.800 73.000 323.600 80.400 ;
        RECT 326.000 71.800 326.800 80.400 ;
        RECT 332.400 71.800 333.200 80.400 ;
        RECT 335.600 75.800 336.400 80.400 ;
        RECT 337.200 75.800 338.000 80.400 ;
        RECT 340.400 75.800 341.200 80.400 ;
        RECT 343.600 75.800 344.400 80.400 ;
        RECT 346.800 75.800 347.600 80.400 ;
        RECT 354.800 75.800 355.600 80.400 ;
        RECT 358.000 75.800 358.800 80.400 ;
        RECT 364.400 75.800 365.200 80.400 ;
        RECT 367.600 75.800 368.400 80.400 ;
        RECT 370.800 75.800 371.600 80.400 ;
        RECT 364.200 71.800 365.200 72.000 ;
        RECT 367.600 71.800 368.400 72.400 ;
        RECT 372.400 71.800 373.200 80.400 ;
        RECT 376.600 75.800 377.400 80.400 ;
        RECT 378.800 71.800 379.600 80.400 ;
        RECT 385.200 71.800 386.000 80.400 ;
        RECT 386.800 71.800 387.600 80.400 ;
        RECT 391.000 75.800 391.800 80.400 ;
        RECT 394.800 75.800 395.600 80.400 ;
        RECT 396.400 75.800 397.200 80.400 ;
        RECT 399.600 75.800 400.400 80.400 ;
        RECT 404.400 71.800 405.200 80.400 ;
        RECT 406.000 75.800 406.800 80.400 ;
        RECT 415.600 75.800 416.400 80.400 ;
        RECT 418.800 75.800 419.600 80.400 ;
        RECT 422.000 75.800 422.800 80.400 ;
        RECT 425.200 75.800 426.000 80.400 ;
        RECT 433.200 75.800 434.000 80.400 ;
        RECT 436.400 75.800 437.200 80.400 ;
        RECT 442.800 75.800 443.600 80.400 ;
        RECT 446.000 75.800 446.800 80.400 ;
        RECT 449.200 75.800 450.000 80.400 ;
        RECT 451.400 75.800 452.200 80.400 ;
        RECT 442.600 71.800 443.400 72.000 ;
        RECT 446.000 71.800 446.800 72.400 ;
        RECT 455.600 71.800 456.400 80.400 ;
        RECT 458.800 75.800 459.600 80.400 ;
        RECT 463.600 73.000 464.400 80.400 ;
        RECT 466.800 75.800 467.600 80.400 ;
        RECT 470.000 75.800 470.800 80.400 ;
        RECT 474.800 73.000 475.600 80.400 ;
        RECT 479.200 71.800 480.000 80.400 ;
        RECT 484.400 72.200 485.200 80.400 ;
        RECT 487.600 75.800 488.400 80.400 ;
        RECT 490.800 75.800 491.600 80.400 ;
        RECT 492.400 71.800 493.200 80.400 ;
        RECT 496.600 75.800 497.400 80.400 ;
        RECT 499.400 75.800 500.200 80.400 ;
        RECT 503.600 71.800 504.400 80.400 ;
        RECT 505.200 75.800 506.000 80.400 ;
        RECT 508.400 75.800 509.200 80.400 ;
        RECT 510.000 75.800 510.800 80.400 ;
        RECT 513.200 75.800 514.000 80.400 ;
        RECT 514.800 75.800 515.600 80.400 ;
        RECT 518.000 75.800 518.800 80.400 ;
        RECT 521.200 75.800 522.000 80.400 ;
        RECT 524.400 75.800 525.200 80.400 ;
        RECT 532.400 75.800 533.200 80.400 ;
        RECT 535.600 75.800 536.400 80.400 ;
        RECT 542.000 75.800 542.800 80.400 ;
        RECT 545.200 75.800 546.000 80.400 ;
        RECT 548.400 75.800 549.200 80.400 ;
        RECT 541.800 71.800 542.600 72.000 ;
        RECT 545.200 71.800 546.000 72.400 ;
        RECT 175.600 71.200 202.600 71.800 ;
        RECT 95.000 71.000 95.800 71.200 ;
        RECT 201.800 71.000 202.600 71.200 ;
        RECT 211.800 71.200 238.800 71.800 ;
        RECT 341.400 71.200 368.400 71.800 ;
        RECT 419.800 71.200 446.800 71.800 ;
        RECT 519.000 71.200 546.000 71.800 ;
        RECT 211.800 71.000 212.600 71.200 ;
        RECT 341.400 71.000 342.200 71.200 ;
        RECT 419.800 71.000 420.600 71.200 ;
        RECT 519.000 71.000 519.800 71.200 ;
        RECT 142.000 70.000 165.400 70.600 ;
        RECT 142.000 69.400 142.800 70.000 ;
        RECT 153.200 69.600 154.000 70.000 ;
        RECT 159.600 69.600 160.400 70.000 ;
        RECT 164.600 69.800 165.400 70.000 ;
        RECT 282.800 70.000 306.200 70.600 ;
        RECT 282.800 69.400 283.600 70.000 ;
        RECT 294.000 69.600 294.800 70.000 ;
        RECT 300.400 69.600 301.200 70.000 ;
        RECT 305.400 69.800 306.200 70.000 ;
        RECT 92.200 52.000 93.000 52.200 ;
        RECT 97.200 52.000 98.000 52.400 ;
        RECT 114.800 52.000 115.600 52.600 ;
        RECT 92.200 51.400 115.600 52.000 ;
        RECT 178.600 52.000 179.400 52.200 ;
        RECT 183.600 52.000 184.400 52.400 ;
        RECT 201.200 52.000 202.000 52.600 ;
        RECT 178.600 51.400 202.000 52.000 ;
        RECT 244.400 52.000 245.200 52.600 ;
        RECT 262.000 52.000 262.800 52.400 ;
        RECT 267.000 52.000 267.800 52.200 ;
        RECT 244.400 51.400 267.800 52.000 ;
        RECT 282.600 52.000 283.400 52.200 ;
        RECT 287.600 52.000 288.400 52.400 ;
        RECT 305.200 52.000 306.000 52.600 ;
        RECT 282.600 51.400 306.000 52.000 ;
        RECT 70.600 50.800 71.400 51.000 ;
        RECT 349.000 50.800 349.800 51.000 ;
        RECT 403.400 50.800 404.200 51.000 ;
        RECT 44.400 50.200 71.400 50.800 ;
        RECT 322.800 50.200 349.800 50.800 ;
        RECT 377.200 50.200 404.200 50.800 ;
        RECT 445.400 50.800 446.200 51.000 ;
        RECT 517.400 50.800 518.200 51.000 ;
        RECT 445.400 50.200 472.400 50.800 ;
        RECT 517.400 50.200 544.400 50.800 ;
        RECT 1.200 41.600 2.000 46.200 ;
        RECT 4.400 41.600 5.200 46.200 ;
        RECT 7.600 41.600 8.400 46.200 ;
        RECT 9.200 41.600 10.000 46.200 ;
        RECT 12.400 41.600 13.200 46.200 ;
        RECT 15.600 41.600 16.400 46.200 ;
        RECT 17.200 41.600 18.000 50.200 ;
        RECT 23.600 41.600 24.400 50.200 ;
        RECT 25.200 41.600 26.000 50.200 ;
        RECT 31.600 41.600 32.400 50.200 ;
        RECT 44.400 49.600 45.200 50.200 ;
        RECT 47.600 50.000 48.600 50.200 ;
        RECT 33.200 41.600 34.000 46.200 ;
        RECT 36.400 41.600 37.200 46.200 ;
        RECT 39.600 41.600 40.400 46.200 ;
        RECT 41.200 41.600 42.000 46.200 ;
        RECT 44.400 41.600 45.200 46.200 ;
        RECT 47.600 41.600 48.400 46.200 ;
        RECT 54.000 41.600 54.800 46.200 ;
        RECT 57.200 41.600 58.000 46.200 ;
        RECT 65.200 41.600 66.000 46.200 ;
        RECT 68.400 41.600 69.200 46.200 ;
        RECT 71.600 41.600 72.400 46.200 ;
        RECT 74.800 41.600 75.600 46.200 ;
        RECT 76.400 41.600 77.200 50.200 ;
        RECT 79.600 41.600 80.400 50.200 ;
        RECT 82.800 41.600 83.600 50.200 ;
        RECT 86.000 41.600 86.800 50.200 ;
        RECT 89.200 41.600 90.000 50.200 ;
        RECT 90.800 41.600 91.600 46.200 ;
        RECT 94.000 41.600 94.800 46.200 ;
        RECT 97.200 41.600 98.000 46.200 ;
        RECT 103.600 41.600 104.400 46.200 ;
        RECT 106.800 41.600 107.600 46.200 ;
        RECT 114.800 41.600 115.600 46.200 ;
        RECT 118.000 41.600 118.800 46.200 ;
        RECT 121.200 41.600 122.000 46.200 ;
        RECT 124.400 41.600 125.200 46.200 ;
        RECT 132.400 41.600 133.200 50.200 ;
        RECT 138.800 41.600 139.600 46.200 ;
        RECT 143.600 41.600 144.400 50.200 ;
        RECT 145.200 41.600 146.000 46.200 ;
        RECT 148.400 41.600 149.200 46.200 ;
        RECT 150.000 41.600 150.800 46.200 ;
        RECT 153.200 41.600 154.000 46.200 ;
        RECT 154.800 41.600 155.600 50.200 ;
        RECT 159.600 41.600 160.400 46.200 ;
        RECT 162.800 41.600 163.600 46.200 ;
        RECT 166.000 41.600 166.800 46.200 ;
        RECT 170.800 41.600 171.600 50.200 ;
        RECT 172.400 41.600 173.200 50.200 ;
        RECT 175.600 41.600 176.400 50.200 ;
        RECT 177.200 41.600 178.000 46.200 ;
        RECT 180.400 41.600 181.200 46.200 ;
        RECT 183.600 41.600 184.400 46.200 ;
        RECT 190.000 41.600 190.800 46.200 ;
        RECT 193.200 41.600 194.000 46.200 ;
        RECT 201.200 41.600 202.000 46.200 ;
        RECT 204.400 41.600 205.200 46.200 ;
        RECT 207.600 41.600 208.400 46.200 ;
        RECT 210.800 41.600 211.600 46.200 ;
        RECT 212.400 41.600 213.200 50.200 ;
        RECT 216.600 41.600 217.400 46.200 ;
        RECT 219.400 41.600 220.200 46.200 ;
        RECT 223.600 41.600 224.400 50.200 ;
        RECT 226.800 41.600 227.600 46.200 ;
        RECT 228.400 41.600 229.200 50.200 ;
        RECT 322.800 49.600 323.600 50.200 ;
        RECT 326.000 50.000 327.000 50.200 ;
        RECT 232.600 41.600 233.400 46.200 ;
        RECT 234.800 41.600 235.600 46.200 ;
        RECT 238.000 41.600 238.800 46.200 ;
        RECT 241.200 41.600 242.000 46.200 ;
        RECT 244.400 41.600 245.200 46.200 ;
        RECT 252.400 41.600 253.200 46.200 ;
        RECT 255.600 41.600 256.400 46.200 ;
        RECT 262.000 41.600 262.800 46.200 ;
        RECT 265.200 41.600 266.000 46.200 ;
        RECT 268.400 41.600 269.200 46.200 ;
        RECT 271.600 41.600 272.400 49.000 ;
        RECT 281.200 41.600 282.000 46.200 ;
        RECT 284.400 41.600 285.200 46.200 ;
        RECT 287.600 41.600 288.400 46.200 ;
        RECT 294.000 41.600 294.800 46.200 ;
        RECT 297.200 41.600 298.000 46.200 ;
        RECT 305.200 41.600 306.000 46.200 ;
        RECT 308.400 41.600 309.200 46.200 ;
        RECT 311.600 41.600 312.400 46.200 ;
        RECT 314.800 41.600 315.600 46.200 ;
        RECT 316.400 41.600 317.200 46.200 ;
        RECT 319.600 41.600 320.400 46.200 ;
        RECT 322.800 41.600 323.600 46.200 ;
        RECT 326.000 41.600 326.800 46.200 ;
        RECT 332.400 41.600 333.200 46.200 ;
        RECT 335.600 41.600 336.400 46.200 ;
        RECT 343.600 41.600 344.400 46.200 ;
        RECT 346.800 41.600 347.600 46.200 ;
        RECT 350.000 41.600 350.800 46.200 ;
        RECT 353.200 41.600 354.000 46.200 ;
        RECT 354.800 41.600 355.600 50.200 ;
        RECT 359.600 41.600 360.400 46.200 ;
        RECT 362.800 41.600 363.600 50.200 ;
        RECT 377.200 49.600 378.000 50.200 ;
        RECT 380.400 50.000 381.400 50.200 ;
        RECT 367.000 41.600 367.800 46.200 ;
        RECT 369.200 41.600 370.000 46.200 ;
        RECT 372.400 41.600 373.200 46.200 ;
        RECT 374.000 41.600 374.800 46.200 ;
        RECT 377.200 41.600 378.000 46.200 ;
        RECT 380.400 41.600 381.200 46.200 ;
        RECT 386.800 41.600 387.600 46.200 ;
        RECT 390.000 41.600 390.800 46.200 ;
        RECT 398.000 41.600 398.800 46.200 ;
        RECT 401.200 41.600 402.000 46.200 ;
        RECT 404.400 41.600 405.200 46.200 ;
        RECT 407.600 41.600 408.400 46.200 ;
        RECT 410.400 41.600 411.200 50.200 ;
        RECT 415.600 41.600 416.400 49.800 ;
        RECT 420.400 41.600 421.200 46.200 ;
        RECT 429.600 41.600 430.400 50.200 ;
        RECT 468.200 50.000 469.200 50.200 ;
        RECT 434.800 41.600 435.600 49.800 ;
        RECT 471.600 49.600 472.400 50.200 ;
        RECT 439.600 41.600 440.400 46.200 ;
        RECT 441.200 41.600 442.000 46.200 ;
        RECT 444.400 41.600 445.200 46.200 ;
        RECT 447.600 41.600 448.400 46.200 ;
        RECT 450.800 41.600 451.600 46.200 ;
        RECT 458.800 41.600 459.600 46.200 ;
        RECT 462.000 41.600 462.800 46.200 ;
        RECT 468.400 41.600 469.200 46.200 ;
        RECT 471.600 41.600 472.400 46.200 ;
        RECT 474.800 41.600 475.600 46.200 ;
        RECT 476.400 41.600 477.200 46.200 ;
        RECT 479.600 41.600 480.400 46.200 ;
        RECT 482.400 41.600 483.200 50.200 ;
        RECT 487.600 41.600 488.400 49.800 ;
        RECT 492.400 41.600 493.200 49.800 ;
        RECT 497.600 41.600 498.400 50.200 ;
        RECT 500.400 41.600 501.200 50.200 ;
        RECT 504.600 41.600 505.400 46.200 ;
        RECT 506.800 41.600 507.600 50.200 ;
        RECT 540.200 50.000 541.200 50.200 ;
        RECT 543.600 49.600 544.400 50.200 ;
        RECT 511.000 41.600 511.800 46.200 ;
        RECT 513.200 41.600 514.000 46.200 ;
        RECT 516.400 41.600 517.200 46.200 ;
        RECT 519.600 41.600 520.400 46.200 ;
        RECT 522.800 41.600 523.600 46.200 ;
        RECT 530.800 41.600 531.600 46.200 ;
        RECT 534.000 41.600 534.800 46.200 ;
        RECT 540.400 41.600 541.200 46.200 ;
        RECT 543.600 41.600 544.400 46.200 ;
        RECT 546.800 41.600 547.600 46.200 ;
        RECT 0.400 40.400 551.600 41.600 ;
        RECT 1.200 35.800 2.000 40.400 ;
        RECT 4.400 35.800 5.200 40.400 ;
        RECT 7.600 35.800 8.400 40.400 ;
        RECT 10.800 35.800 11.600 40.400 ;
        RECT 18.800 35.800 19.600 40.400 ;
        RECT 22.000 35.800 22.800 40.400 ;
        RECT 28.400 35.800 29.200 40.400 ;
        RECT 31.600 35.800 32.400 40.400 ;
        RECT 34.800 35.800 35.600 40.400 ;
        RECT 36.400 35.800 37.200 40.400 ;
        RECT 39.600 35.800 40.400 40.400 ;
        RECT 42.800 35.800 43.600 40.400 ;
        RECT 46.000 35.800 46.800 40.400 ;
        RECT 54.000 35.800 54.800 40.400 ;
        RECT 57.200 35.800 58.000 40.400 ;
        RECT 63.600 35.800 64.400 40.400 ;
        RECT 66.800 35.800 67.600 40.400 ;
        RECT 70.000 35.800 70.800 40.400 ;
        RECT 73.200 33.000 74.000 40.400 ;
        RECT 28.200 31.800 29.000 32.000 ;
        RECT 31.600 31.800 32.400 32.400 ;
        RECT 63.400 31.800 64.200 32.000 ;
        RECT 66.800 31.800 67.600 32.400 ;
        RECT 76.400 31.800 77.200 40.400 ;
        RECT 79.600 31.800 80.400 40.400 ;
        RECT 82.800 31.800 83.600 40.400 ;
        RECT 86.000 31.800 86.800 40.400 ;
        RECT 89.200 31.800 90.000 40.400 ;
        RECT 90.800 35.800 91.600 40.400 ;
        RECT 94.000 35.800 94.800 40.400 ;
        RECT 97.200 35.800 98.000 40.400 ;
        RECT 103.600 35.800 104.400 40.400 ;
        RECT 106.800 35.800 107.600 40.400 ;
        RECT 114.800 35.800 115.600 40.400 ;
        RECT 118.000 35.800 118.800 40.400 ;
        RECT 121.200 35.800 122.000 40.400 ;
        RECT 124.400 35.800 125.200 40.400 ;
        RECT 132.400 35.800 133.200 40.400 ;
        RECT 135.600 35.800 136.400 40.400 ;
        RECT 138.800 35.800 139.600 40.400 ;
        RECT 142.000 35.800 142.800 40.400 ;
        RECT 150.000 35.800 150.800 40.400 ;
        RECT 153.200 35.600 154.000 40.400 ;
        RECT 159.600 35.800 160.400 40.400 ;
        RECT 162.800 35.800 163.600 40.400 ;
        RECT 166.000 35.800 166.800 40.400 ;
        RECT 167.600 35.800 168.400 40.400 ;
        RECT 170.800 35.800 171.600 40.400 ;
        RECT 174.000 35.800 174.800 40.400 ;
        RECT 177.200 35.800 178.000 40.400 ;
        RECT 185.200 35.800 186.000 40.400 ;
        RECT 188.400 35.600 189.200 40.400 ;
        RECT 194.800 35.800 195.600 40.400 ;
        RECT 198.000 35.800 198.800 40.400 ;
        RECT 201.200 35.800 202.000 40.400 ;
        RECT 202.800 35.800 203.600 40.400 ;
        RECT 206.000 35.800 206.800 40.400 ;
        RECT 208.200 35.800 209.000 40.400 ;
        RECT 94.000 31.800 94.800 32.400 ;
        RECT 97.200 31.800 98.200 32.000 ;
        RECT 212.400 31.800 213.200 40.400 ;
        RECT 214.000 35.800 214.800 40.400 ;
        RECT 217.200 31.800 218.000 40.400 ;
        RECT 221.400 35.800 222.200 40.400 ;
        RECT 223.600 31.800 224.400 40.400 ;
        RECT 227.800 35.800 228.600 40.400 ;
        RECT 230.000 35.800 230.800 40.400 ;
        RECT 233.200 35.800 234.000 40.400 ;
        RECT 236.400 35.800 237.200 40.400 ;
        RECT 239.600 35.800 240.400 40.400 ;
        RECT 247.600 35.800 248.400 40.400 ;
        RECT 250.800 35.600 251.600 40.400 ;
        RECT 257.200 35.800 258.000 40.400 ;
        RECT 260.400 35.800 261.200 40.400 ;
        RECT 263.600 35.800 264.400 40.400 ;
        RECT 265.200 35.800 266.000 40.400 ;
        RECT 268.400 31.800 269.200 40.400 ;
        RECT 272.600 35.800 273.400 40.400 ;
        RECT 281.800 35.800 282.600 40.400 ;
        RECT 286.000 31.800 286.800 40.400 ;
        RECT 287.600 35.800 288.400 40.400 ;
        RECT 290.800 35.800 291.600 40.400 ;
        RECT 294.000 35.800 294.800 40.400 ;
        RECT 297.200 35.800 298.000 40.400 ;
        RECT 305.200 35.800 306.000 40.400 ;
        RECT 308.400 35.600 309.200 40.400 ;
        RECT 314.800 35.800 315.600 40.400 ;
        RECT 318.000 35.800 318.800 40.400 ;
        RECT 321.200 35.800 322.000 40.400 ;
        RECT 322.800 35.800 323.600 40.400 ;
        RECT 326.000 35.800 326.800 40.400 ;
        RECT 329.200 35.800 330.000 40.400 ;
        RECT 332.400 35.800 333.200 40.400 ;
        RECT 340.400 35.800 341.200 40.400 ;
        RECT 343.600 35.800 344.400 40.400 ;
        RECT 350.000 35.800 350.800 40.400 ;
        RECT 353.200 35.800 354.000 40.400 ;
        RECT 356.400 35.800 357.200 40.400 ;
        RECT 349.800 31.800 350.800 32.000 ;
        RECT 353.200 31.800 354.000 32.400 ;
        RECT 358.000 31.800 358.800 40.400 ;
        RECT 361.200 31.800 362.000 40.400 ;
        RECT 364.400 31.800 365.200 40.400 ;
        RECT 367.600 31.800 368.400 40.400 ;
        RECT 370.800 31.800 371.600 40.400 ;
        RECT 372.400 35.800 373.200 40.400 ;
        RECT 375.600 35.800 376.400 40.400 ;
        RECT 378.800 35.800 379.600 40.400 ;
        RECT 385.200 35.800 386.000 40.400 ;
        RECT 388.400 35.800 389.200 40.400 ;
        RECT 396.400 35.800 397.200 40.400 ;
        RECT 399.600 35.800 400.400 40.400 ;
        RECT 402.800 35.800 403.600 40.400 ;
        RECT 406.000 35.800 406.800 40.400 ;
        RECT 407.600 35.800 408.400 40.400 ;
        RECT 417.200 35.800 418.000 40.400 ;
        RECT 420.400 35.800 421.200 40.400 ;
        RECT 423.600 35.800 424.400 40.400 ;
        RECT 430.000 35.800 430.800 40.400 ;
        RECT 433.200 35.800 434.000 40.400 ;
        RECT 441.200 35.800 442.000 40.400 ;
        RECT 444.400 35.800 445.200 40.400 ;
        RECT 447.600 35.800 448.400 40.400 ;
        RECT 450.800 35.800 451.600 40.400 ;
        RECT 375.600 31.800 376.400 32.400 ;
        RECT 379.000 31.800 379.800 32.000 ;
        RECT 420.400 31.800 421.200 32.400 ;
        RECT 423.800 31.800 424.600 32.000 ;
        RECT 454.000 31.800 454.800 40.400 ;
        RECT 459.600 35.800 460.400 40.400 ;
        RECT 462.800 35.800 463.600 40.400 ;
        RECT 468.400 32.000 469.200 40.400 ;
        RECT 471.600 35.800 472.400 40.400 ;
        RECT 474.800 31.800 475.600 40.400 ;
        RECT 479.000 35.800 479.800 40.400 ;
        RECT 481.200 35.800 482.000 40.400 ;
        RECT 484.400 35.800 485.200 40.400 ;
        RECT 487.600 35.800 488.400 40.400 ;
        RECT 490.800 35.800 491.600 40.400 ;
        RECT 498.800 35.800 499.600 40.400 ;
        RECT 502.000 35.800 502.800 40.400 ;
        RECT 508.400 35.800 509.200 40.400 ;
        RECT 511.600 35.800 512.400 40.400 ;
        RECT 514.800 35.800 515.600 40.400 ;
        RECT 508.200 31.800 509.200 32.000 ;
        RECT 511.600 31.800 512.400 32.400 ;
        RECT 517.600 31.800 518.400 40.400 ;
        RECT 522.800 32.200 523.600 40.400 ;
        RECT 527.600 32.200 528.400 40.400 ;
        RECT 532.800 31.800 533.600 40.400 ;
        RECT 535.600 31.800 536.400 40.400 ;
        RECT 538.800 31.800 539.600 40.400 ;
        RECT 542.000 31.800 542.800 40.400 ;
        RECT 545.200 31.800 546.000 40.400 ;
        RECT 548.400 31.800 549.200 40.400 ;
        RECT 5.400 31.200 32.400 31.800 ;
        RECT 40.600 31.200 67.600 31.800 ;
        RECT 94.000 31.200 121.000 31.800 ;
        RECT 5.400 31.000 6.200 31.200 ;
        RECT 40.600 31.000 41.400 31.200 ;
        RECT 120.200 31.000 121.000 31.200 ;
        RECT 327.000 31.200 354.000 31.800 ;
        RECT 375.600 31.200 402.600 31.800 ;
        RECT 420.400 31.200 447.400 31.800 ;
        RECT 327.000 31.000 327.800 31.200 ;
        RECT 401.800 31.000 402.600 31.200 ;
        RECT 446.600 31.000 447.400 31.200 ;
        RECT 485.400 31.200 512.400 31.800 ;
        RECT 485.400 31.000 486.200 31.200 ;
        RECT 142.000 30.000 165.400 30.600 ;
        RECT 142.000 29.400 142.800 30.000 ;
        RECT 153.200 29.600 154.000 30.000 ;
        RECT 159.600 29.600 160.400 30.000 ;
        RECT 164.600 29.800 165.400 30.000 ;
        RECT 177.200 30.000 200.600 30.600 ;
        RECT 177.200 29.400 178.000 30.000 ;
        RECT 188.400 29.600 189.200 30.000 ;
        RECT 194.800 29.600 195.600 30.000 ;
        RECT 199.800 29.800 200.600 30.000 ;
        RECT 239.600 30.000 263.000 30.600 ;
        RECT 239.600 29.400 240.400 30.000 ;
        RECT 250.800 29.600 251.600 30.000 ;
        RECT 257.200 29.600 258.000 30.000 ;
        RECT 262.200 29.800 263.000 30.000 ;
        RECT 297.200 30.000 320.600 30.600 ;
        RECT 297.200 29.400 298.000 30.000 ;
        RECT 308.400 29.600 309.200 30.000 ;
        RECT 314.800 29.600 315.600 30.000 ;
        RECT 319.800 29.800 320.600 30.000 ;
        RECT 183.400 12.000 184.200 12.200 ;
        RECT 188.400 12.000 189.200 12.400 ;
        RECT 206.000 12.000 206.800 12.600 ;
        RECT 183.400 11.400 206.800 12.000 ;
        RECT 298.800 12.000 299.600 12.600 ;
        RECT 316.400 12.000 317.200 12.400 ;
        RECT 321.400 12.000 322.200 12.200 ;
        RECT 298.800 11.400 322.200 12.000 ;
        RECT 5.400 10.800 6.200 11.000 ;
        RECT 65.800 10.800 66.600 11.000 ;
        RECT 113.800 10.800 114.600 11.000 ;
        RECT 5.400 10.200 32.400 10.800 ;
        RECT 28.200 10.000 29.000 10.200 ;
        RECT 31.600 9.600 32.400 10.200 ;
        RECT 39.600 10.200 66.600 10.800 ;
        RECT 87.600 10.200 114.600 10.800 ;
        RECT 141.400 10.800 142.200 11.000 ;
        RECT 341.400 10.800 342.200 11.000 ;
        RECT 425.800 10.800 426.600 11.000 ;
        RECT 496.200 10.800 497.000 11.000 ;
        RECT 534.600 10.800 535.400 11.000 ;
        RECT 141.400 10.200 168.400 10.800 ;
        RECT 341.400 10.200 368.400 10.800 ;
        RECT 399.600 10.200 426.600 10.800 ;
        RECT 470.000 10.200 497.000 10.800 ;
        RECT 508.400 10.200 535.400 10.800 ;
        RECT 39.600 9.600 40.400 10.200 ;
        RECT 42.800 10.000 43.800 10.200 ;
        RECT 1.200 1.600 2.000 6.200 ;
        RECT 4.400 1.600 5.200 6.200 ;
        RECT 7.600 1.600 8.400 6.200 ;
        RECT 10.800 1.600 11.600 6.200 ;
        RECT 18.800 1.600 19.600 6.200 ;
        RECT 22.000 1.600 22.800 6.200 ;
        RECT 28.400 1.600 29.200 6.200 ;
        RECT 31.600 1.600 32.400 6.200 ;
        RECT 34.800 1.600 35.600 6.200 ;
        RECT 36.400 1.600 37.200 6.200 ;
        RECT 39.600 1.600 40.400 6.200 ;
        RECT 42.800 1.600 43.600 6.200 ;
        RECT 49.200 1.600 50.000 6.200 ;
        RECT 52.400 1.600 53.200 6.200 ;
        RECT 60.400 1.600 61.200 6.200 ;
        RECT 63.600 1.600 64.400 6.200 ;
        RECT 66.800 1.600 67.600 6.200 ;
        RECT 70.000 1.600 70.800 6.200 ;
        RECT 73.200 1.600 74.000 9.800 ;
        RECT 76.400 1.600 77.200 6.200 ;
        RECT 78.000 1.600 78.800 6.200 ;
        RECT 81.200 1.600 82.000 9.800 ;
        RECT 87.600 9.600 88.400 10.200 ;
        RECT 91.000 10.000 91.800 10.200 ;
        RECT 84.400 1.600 85.200 6.200 ;
        RECT 87.600 1.600 88.400 6.200 ;
        RECT 90.800 1.600 91.600 6.200 ;
        RECT 97.200 1.600 98.000 6.200 ;
        RECT 100.400 1.600 101.200 6.200 ;
        RECT 108.400 1.600 109.200 6.200 ;
        RECT 111.600 1.600 112.400 6.200 ;
        RECT 114.800 1.600 115.600 6.200 ;
        RECT 118.000 1.600 118.800 6.200 ;
        RECT 119.600 1.600 120.400 10.200 ;
        RECT 131.400 1.600 132.200 6.200 ;
        RECT 135.600 1.600 136.400 10.200 ;
        RECT 164.200 10.000 165.200 10.200 ;
        RECT 167.600 9.600 168.400 10.200 ;
        RECT 137.200 1.600 138.000 6.200 ;
        RECT 140.400 1.600 141.200 6.200 ;
        RECT 143.600 1.600 144.400 6.200 ;
        RECT 146.800 1.600 147.600 6.200 ;
        RECT 154.800 1.600 155.600 6.200 ;
        RECT 158.000 1.600 158.800 6.200 ;
        RECT 164.400 1.600 165.200 6.200 ;
        RECT 167.600 1.600 168.400 6.200 ;
        RECT 170.800 1.600 171.600 6.200 ;
        RECT 174.000 1.600 174.800 9.000 ;
        RECT 178.800 1.600 179.600 9.000 ;
        RECT 182.000 1.600 182.800 6.200 ;
        RECT 185.200 1.600 186.000 6.200 ;
        RECT 188.400 1.600 189.200 6.200 ;
        RECT 194.800 1.600 195.600 6.200 ;
        RECT 198.000 1.600 198.800 6.200 ;
        RECT 206.000 1.600 206.800 6.200 ;
        RECT 209.200 1.600 210.000 6.200 ;
        RECT 212.400 1.600 213.200 6.200 ;
        RECT 215.600 1.600 216.400 6.200 ;
        RECT 217.200 1.600 218.000 6.200 ;
        RECT 220.400 1.600 221.200 10.200 ;
        RECT 224.600 1.600 225.400 6.200 ;
        RECT 226.800 1.600 227.600 10.200 ;
        RECT 231.000 1.600 231.800 6.200 ;
        RECT 233.200 1.600 234.000 6.200 ;
        RECT 236.400 1.600 237.200 6.200 ;
        RECT 238.000 1.600 238.800 10.200 ;
        RECT 242.200 1.600 243.000 6.200 ;
        RECT 244.400 1.600 245.200 10.200 ;
        RECT 248.600 1.600 249.400 6.200 ;
        RECT 251.400 1.600 252.200 6.200 ;
        RECT 255.600 1.600 256.400 10.200 ;
        RECT 257.800 1.600 258.600 6.200 ;
        RECT 262.000 1.600 262.800 10.200 ;
        RECT 265.200 1.600 266.000 6.200 ;
        RECT 266.800 1.600 267.600 6.200 ;
        RECT 270.000 1.600 270.800 10.200 ;
        RECT 274.200 1.600 275.000 6.200 ;
        RECT 282.800 1.600 283.600 10.200 ;
        RECT 364.200 10.000 365.200 10.200 ;
        RECT 287.000 1.600 287.800 6.200 ;
        RECT 289.200 1.600 290.000 6.200 ;
        RECT 292.400 1.600 293.200 6.200 ;
        RECT 295.600 1.600 296.400 6.200 ;
        RECT 298.800 1.600 299.600 6.200 ;
        RECT 306.800 1.600 307.600 6.200 ;
        RECT 310.000 1.600 310.800 6.200 ;
        RECT 316.400 1.600 317.200 6.200 ;
        RECT 319.600 1.600 320.400 6.200 ;
        RECT 322.800 1.600 323.600 6.200 ;
        RECT 324.400 1.600 325.200 6.200 ;
        RECT 327.600 1.600 328.400 9.800 ;
        RECT 330.800 1.600 331.600 6.200 ;
        RECT 334.000 1.600 334.800 9.800 ;
        RECT 367.600 9.600 368.400 10.200 ;
        RECT 337.200 1.600 338.000 6.200 ;
        RECT 340.400 1.600 341.200 6.200 ;
        RECT 343.600 1.600 344.400 6.200 ;
        RECT 346.800 1.600 347.600 6.200 ;
        RECT 354.800 1.600 355.600 6.200 ;
        RECT 358.000 1.600 358.800 6.200 ;
        RECT 364.400 1.600 365.200 6.200 ;
        RECT 367.600 1.600 368.400 6.200 ;
        RECT 370.800 1.600 371.600 6.200 ;
        RECT 374.000 1.600 374.800 9.000 ;
        RECT 378.800 1.600 379.600 10.200 ;
        RECT 384.400 1.600 385.200 6.200 ;
        RECT 387.600 1.600 388.400 6.200 ;
        RECT 393.200 1.600 394.000 10.000 ;
        RECT 399.600 9.600 400.400 10.200 ;
        RECT 403.000 10.000 403.800 10.200 ;
        RECT 396.400 1.600 397.200 6.200 ;
        RECT 399.600 1.600 400.400 6.200 ;
        RECT 402.800 1.600 403.600 6.200 ;
        RECT 409.200 1.600 410.000 6.200 ;
        RECT 412.400 1.600 413.200 6.200 ;
        RECT 420.400 1.600 421.200 6.200 ;
        RECT 423.600 1.600 424.400 6.200 ;
        RECT 426.800 1.600 427.600 6.200 ;
        RECT 430.000 1.600 430.800 6.200 ;
        RECT 439.600 1.600 440.400 10.000 ;
        RECT 445.200 1.600 446.000 6.200 ;
        RECT 448.400 1.600 449.200 6.200 ;
        RECT 454.000 1.600 454.800 10.200 ;
        RECT 470.000 9.600 470.800 10.200 ;
        RECT 473.400 10.000 474.200 10.200 ;
        RECT 508.400 9.600 509.200 10.200 ;
        RECT 511.800 10.000 512.600 10.200 ;
        RECT 458.800 1.600 459.600 9.000 ;
        RECT 463.600 1.600 464.400 9.000 ;
        RECT 466.800 1.600 467.600 6.200 ;
        RECT 470.000 1.600 470.800 6.200 ;
        RECT 473.200 1.600 474.000 6.200 ;
        RECT 479.600 1.600 480.400 6.200 ;
        RECT 482.800 1.600 483.600 6.200 ;
        RECT 490.800 1.600 491.600 6.200 ;
        RECT 494.000 1.600 494.800 6.200 ;
        RECT 497.200 1.600 498.000 6.200 ;
        RECT 500.400 1.600 501.200 6.200 ;
        RECT 502.000 1.600 502.800 6.200 ;
        RECT 505.200 1.600 506.000 6.200 ;
        RECT 508.400 1.600 509.200 6.200 ;
        RECT 511.600 1.600 512.400 6.200 ;
        RECT 518.000 1.600 518.800 6.200 ;
        RECT 521.200 1.600 522.000 6.200 ;
        RECT 529.200 1.600 530.000 6.200 ;
        RECT 532.400 1.600 533.200 6.200 ;
        RECT 535.600 1.600 536.400 6.200 ;
        RECT 538.800 1.600 539.600 6.200 ;
        RECT 542.000 1.600 542.800 9.000 ;
        RECT 546.800 1.600 547.600 9.000 ;
        RECT 0.400 0.400 551.600 1.600 ;
      LAYER via1 ;
        RECT 372.400 371.600 373.200 372.400 ;
        RECT 98.800 370.000 99.600 370.800 ;
        RECT 31.600 363.600 32.400 364.400 ;
        RECT 42.800 363.600 43.600 364.400 ;
        RECT 98.800 365.400 99.600 366.200 ;
        RECT 143.600 363.600 144.400 364.400 ;
        RECT 154.800 363.600 155.600 364.400 ;
        RECT 190.000 363.600 190.800 364.400 ;
        RECT 282.800 363.600 283.600 364.400 ;
        RECT 372.400 365.400 373.200 366.200 ;
        RECT 538.800 370.000 539.600 370.800 ;
        RECT 398.000 363.600 398.800 364.400 ;
        RECT 466.800 363.600 467.600 364.400 ;
        RECT 478.000 365.400 478.800 366.200 ;
        RECT 538.800 363.600 539.600 364.400 ;
        RECT 121.900 360.600 122.700 361.400 ;
        RECT 122.900 360.600 123.700 361.400 ;
        RECT 123.900 360.600 124.700 361.400 ;
        RECT 124.900 360.600 125.700 361.400 ;
        RECT 125.900 360.600 126.700 361.400 ;
        RECT 126.900 360.600 127.700 361.400 ;
        RECT 422.700 360.600 423.500 361.400 ;
        RECT 423.700 360.600 424.500 361.400 ;
        RECT 424.700 360.600 425.500 361.400 ;
        RECT 425.700 360.600 426.500 361.400 ;
        RECT 426.700 360.600 427.500 361.400 ;
        RECT 427.700 360.600 428.500 361.400 ;
        RECT 31.600 357.600 32.400 358.400 ;
        RECT 31.600 351.600 32.400 352.400 ;
        RECT 65.200 351.200 66.000 352.000 ;
        RECT 143.600 357.600 144.400 358.400 ;
        RECT 268.400 357.600 269.200 358.400 ;
        RECT 105.200 351.200 106.000 352.000 ;
        RECT 143.600 351.600 144.400 352.400 ;
        RECT 202.800 351.200 203.600 352.000 ;
        RECT 238.000 351.200 238.800 352.000 ;
        RECT 268.400 351.600 269.200 352.400 ;
        RECT 545.200 357.600 546.000 358.400 ;
        RECT 545.200 351.600 546.000 352.400 ;
        RECT 34.800 323.600 35.600 324.400 ;
        RECT 121.200 330.000 122.000 330.800 ;
        RECT 121.200 325.400 122.000 326.200 ;
        RECT 142.000 323.600 142.800 324.400 ;
        RECT 246.000 330.000 246.800 330.800 ;
        RECT 246.000 325.400 246.800 326.200 ;
        RECT 278.000 323.600 278.800 324.400 ;
        RECT 316.400 325.400 317.200 326.200 ;
        RECT 462.000 323.600 462.800 324.400 ;
        RECT 121.900 320.600 122.700 321.400 ;
        RECT 122.900 320.600 123.700 321.400 ;
        RECT 123.900 320.600 124.700 321.400 ;
        RECT 124.900 320.600 125.700 321.400 ;
        RECT 125.900 320.600 126.700 321.400 ;
        RECT 126.900 320.600 127.700 321.400 ;
        RECT 422.700 320.600 423.500 321.400 ;
        RECT 423.700 320.600 424.500 321.400 ;
        RECT 424.700 320.600 425.500 321.400 ;
        RECT 425.700 320.600 426.500 321.400 ;
        RECT 426.700 320.600 427.500 321.400 ;
        RECT 427.700 320.600 428.500 321.400 ;
        RECT 279.600 317.600 280.400 318.400 ;
        RECT 279.600 311.600 280.400 312.400 ;
        RECT 444.400 317.600 445.200 318.400 ;
        RECT 444.400 311.600 445.200 312.400 ;
        RECT 65.200 290.000 66.000 290.800 ;
        RECT 100.400 290.000 101.200 290.800 ;
        RECT 65.200 285.400 66.000 286.200 ;
        RECT 100.400 283.600 101.200 284.400 ;
        RECT 302.000 290.000 302.800 290.800 ;
        RECT 302.000 285.400 302.800 286.200 ;
        RECT 478.000 290.000 478.800 290.800 ;
        RECT 478.000 285.400 478.800 286.200 ;
        RECT 540.400 290.000 541.200 290.800 ;
        RECT 540.400 285.400 541.200 286.200 ;
        RECT 121.900 280.600 122.700 281.400 ;
        RECT 122.900 280.600 123.700 281.400 ;
        RECT 123.900 280.600 124.700 281.400 ;
        RECT 124.900 280.600 125.700 281.400 ;
        RECT 125.900 280.600 126.700 281.400 ;
        RECT 126.900 280.600 127.700 281.400 ;
        RECT 422.700 280.600 423.500 281.400 ;
        RECT 423.700 280.600 424.500 281.400 ;
        RECT 424.700 280.600 425.500 281.400 ;
        RECT 425.700 280.600 426.500 281.400 ;
        RECT 426.700 280.600 427.500 281.400 ;
        RECT 427.700 280.600 428.500 281.400 ;
        RECT 31.600 277.600 32.400 278.400 ;
        RECT 31.600 271.600 32.400 272.400 ;
        RECT 97.200 271.200 98.000 272.000 ;
        RECT 390.000 271.200 390.800 272.000 ;
        RECT 482.800 277.600 483.600 278.400 ;
        RECT 518.000 277.600 518.800 278.400 ;
        RECT 482.800 271.600 483.600 272.400 ;
        RECT 518.000 271.600 518.800 272.400 ;
        RECT 255.600 251.600 256.400 252.400 ;
        RECT 297.200 251.600 298.000 252.400 ;
        RECT 106.800 250.000 107.600 250.800 ;
        RECT 106.800 245.400 107.600 246.200 ;
        RECT 151.600 245.400 152.400 246.200 ;
        RECT 236.400 243.600 237.200 244.400 ;
        RECT 255.600 245.400 256.400 246.200 ;
        RECT 297.200 245.400 298.000 246.200 ;
        RECT 415.600 250.000 416.400 250.800 ;
        RECT 460.400 250.000 461.200 250.800 ;
        RECT 356.400 245.400 357.200 246.200 ;
        RECT 415.600 243.600 416.400 244.400 ;
        RECT 460.400 245.400 461.200 246.200 ;
        RECT 486.000 245.400 486.800 246.200 ;
        RECT 121.900 240.600 122.700 241.400 ;
        RECT 122.900 240.600 123.700 241.400 ;
        RECT 123.900 240.600 124.700 241.400 ;
        RECT 124.900 240.600 125.700 241.400 ;
        RECT 125.900 240.600 126.700 241.400 ;
        RECT 126.900 240.600 127.700 241.400 ;
        RECT 422.700 240.600 423.500 241.400 ;
        RECT 423.700 240.600 424.500 241.400 ;
        RECT 424.700 240.600 425.500 241.400 ;
        RECT 425.700 240.600 426.500 241.400 ;
        RECT 426.700 240.600 427.500 241.400 ;
        RECT 427.700 240.600 428.500 241.400 ;
        RECT 31.600 237.600 32.400 238.400 ;
        RECT 31.600 231.600 32.400 232.400 ;
        RECT 130.800 231.200 131.600 232.000 ;
        RECT 234.800 237.600 235.600 238.400 ;
        RECT 234.800 231.600 235.600 232.400 ;
        RECT 266.800 231.200 267.600 232.000 ;
        RECT 404.400 231.200 405.200 232.000 ;
        RECT 526.000 237.600 526.800 238.400 ;
        RECT 526.000 231.600 526.800 232.400 ;
        RECT 300.400 211.600 301.200 212.400 ;
        RECT 119.600 203.600 120.400 204.400 ;
        RECT 273.200 210.000 274.000 210.800 ;
        RECT 273.200 203.600 274.000 204.400 ;
        RECT 300.400 205.400 301.200 206.200 ;
        RECT 510.000 203.600 510.800 204.400 ;
        RECT 521.200 205.400 522.000 206.200 ;
        RECT 121.900 200.600 122.700 201.400 ;
        RECT 122.900 200.600 123.700 201.400 ;
        RECT 123.900 200.600 124.700 201.400 ;
        RECT 124.900 200.600 125.700 201.400 ;
        RECT 125.900 200.600 126.700 201.400 ;
        RECT 126.900 200.600 127.700 201.400 ;
        RECT 422.700 200.600 423.500 201.400 ;
        RECT 423.700 200.600 424.500 201.400 ;
        RECT 424.700 200.600 425.500 201.400 ;
        RECT 425.700 200.600 426.500 201.400 ;
        RECT 426.700 200.600 427.500 201.400 ;
        RECT 427.700 200.600 428.500 201.400 ;
        RECT 146.800 197.600 147.600 198.400 ;
        RECT 73.200 191.200 74.000 192.000 ;
        RECT 146.800 191.600 147.600 192.400 ;
        RECT 212.400 197.600 213.200 198.400 ;
        RECT 212.400 191.600 213.200 192.400 ;
        RECT 294.000 191.200 294.800 192.000 ;
        RECT 498.800 197.600 499.600 198.400 ;
        RECT 498.800 191.600 499.600 192.400 ;
        RECT 126.000 171.600 126.800 172.400 ;
        RECT 82.800 170.000 83.600 170.800 ;
        RECT 82.800 163.600 83.600 164.400 ;
        RECT 126.000 165.400 126.800 166.200 ;
        RECT 154.800 163.600 155.600 164.400 ;
        RECT 231.600 163.600 232.400 164.400 ;
        RECT 324.400 163.600 325.200 164.400 ;
        RECT 370.800 163.600 371.600 164.400 ;
        RECT 444.400 170.000 445.200 170.800 ;
        RECT 444.400 165.400 445.200 166.200 ;
        RECT 540.400 170.000 541.200 170.800 ;
        RECT 540.400 165.400 541.200 166.200 ;
        RECT 121.900 160.600 122.700 161.400 ;
        RECT 122.900 160.600 123.700 161.400 ;
        RECT 123.900 160.600 124.700 161.400 ;
        RECT 124.900 160.600 125.700 161.400 ;
        RECT 125.900 160.600 126.700 161.400 ;
        RECT 126.900 160.600 127.700 161.400 ;
        RECT 422.700 160.600 423.500 161.400 ;
        RECT 423.700 160.600 424.500 161.400 ;
        RECT 424.700 160.600 425.500 161.400 ;
        RECT 425.700 160.600 426.500 161.400 ;
        RECT 426.700 160.600 427.500 161.400 ;
        RECT 427.700 160.600 428.500 161.400 ;
        RECT 97.200 151.200 98.000 152.000 ;
        RECT 151.600 157.600 152.400 158.400 ;
        RECT 151.600 151.600 152.400 152.400 ;
        RECT 228.400 151.200 229.200 152.000 ;
        RECT 281.200 131.600 282.000 132.400 ;
        RECT 76.400 130.000 77.200 130.800 ;
        RECT 76.400 123.600 77.200 124.400 ;
        RECT 105.200 125.400 106.000 126.200 ;
        RECT 212.400 123.600 213.200 124.400 ;
        RECT 281.200 125.400 282.000 126.200 ;
        RECT 329.200 123.600 330.000 124.400 ;
        RECT 422.000 130.000 422.800 130.800 ;
        RECT 422.000 125.400 422.800 126.200 ;
        RECT 468.400 123.600 469.200 124.400 ;
        RECT 545.200 123.600 546.000 124.400 ;
        RECT 121.900 120.600 122.700 121.400 ;
        RECT 122.900 120.600 123.700 121.400 ;
        RECT 123.900 120.600 124.700 121.400 ;
        RECT 124.900 120.600 125.700 121.400 ;
        RECT 125.900 120.600 126.700 121.400 ;
        RECT 126.900 120.600 127.700 121.400 ;
        RECT 422.700 120.600 423.500 121.400 ;
        RECT 423.700 120.600 424.500 121.400 ;
        RECT 424.700 120.600 425.500 121.400 ;
        RECT 425.700 120.600 426.500 121.400 ;
        RECT 426.700 120.600 427.500 121.400 ;
        RECT 427.700 120.600 428.500 121.400 ;
        RECT 73.200 117.600 74.000 118.400 ;
        RECT 73.200 111.600 74.000 112.400 ;
        RECT 87.600 117.600 88.400 118.400 ;
        RECT 87.600 111.600 88.400 112.400 ;
        RECT 183.600 117.600 184.400 118.400 ;
        RECT 183.600 111.600 184.400 112.400 ;
        RECT 342.000 117.600 342.800 118.400 ;
        RECT 342.000 111.600 342.800 112.400 ;
        RECT 546.800 117.600 547.600 118.400 ;
        RECT 546.800 111.600 547.600 112.400 ;
        RECT 70.000 91.600 70.800 92.400 ;
        RECT 316.400 91.600 317.200 92.400 ;
        RECT 70.000 85.400 70.800 86.200 ;
        RECT 105.200 85.400 106.000 86.200 ;
        RECT 298.800 83.600 299.600 84.400 ;
        RECT 316.400 85.400 317.200 86.200 ;
        RECT 361.200 83.600 362.000 84.400 ;
        RECT 508.400 90.000 509.200 90.800 ;
        RECT 543.600 90.000 544.400 90.800 ;
        RECT 508.400 85.400 509.200 86.200 ;
        RECT 543.600 83.600 544.400 84.400 ;
        RECT 121.900 80.600 122.700 81.400 ;
        RECT 122.900 80.600 123.700 81.400 ;
        RECT 123.900 80.600 124.700 81.400 ;
        RECT 124.900 80.600 125.700 81.400 ;
        RECT 125.900 80.600 126.700 81.400 ;
        RECT 126.900 80.600 127.700 81.400 ;
        RECT 422.700 80.600 423.500 81.400 ;
        RECT 423.700 80.600 424.500 81.400 ;
        RECT 424.700 80.600 425.500 81.400 ;
        RECT 425.700 80.600 426.500 81.400 ;
        RECT 426.700 80.600 427.500 81.400 ;
        RECT 427.700 80.600 428.500 81.400 ;
        RECT 121.200 77.600 122.000 78.400 ;
        RECT 175.600 77.600 176.400 78.400 ;
        RECT 121.200 71.600 122.000 72.400 ;
        RECT 175.600 71.600 176.400 72.400 ;
        RECT 234.800 71.200 235.600 72.000 ;
        RECT 364.400 71.200 365.200 72.000 ;
        RECT 446.000 77.600 446.800 78.400 ;
        RECT 446.000 71.600 446.800 72.400 ;
        RECT 545.200 77.600 546.000 78.400 ;
        RECT 545.200 71.600 546.000 72.400 ;
        RECT 114.800 51.600 115.600 52.400 ;
        RECT 201.200 51.600 202.000 52.400 ;
        RECT 244.400 51.600 245.200 52.400 ;
        RECT 305.200 51.600 306.000 52.400 ;
        RECT 47.600 43.600 48.400 44.400 ;
        RECT 114.800 45.400 115.600 46.200 ;
        RECT 201.200 45.400 202.000 46.200 ;
        RECT 244.400 45.400 245.200 46.200 ;
        RECT 305.200 45.400 306.000 46.200 ;
        RECT 326.000 45.400 326.800 46.200 ;
        RECT 380.400 45.400 381.200 46.200 ;
        RECT 468.400 50.000 469.200 50.800 ;
        RECT 468.400 45.400 469.200 46.200 ;
        RECT 540.400 50.000 541.200 50.800 ;
        RECT 540.400 45.400 541.200 46.200 ;
        RECT 121.900 40.600 122.700 41.400 ;
        RECT 122.900 40.600 123.700 41.400 ;
        RECT 123.900 40.600 124.700 41.400 ;
        RECT 124.900 40.600 125.700 41.400 ;
        RECT 125.900 40.600 126.700 41.400 ;
        RECT 126.900 40.600 127.700 41.400 ;
        RECT 422.700 40.600 423.500 41.400 ;
        RECT 423.700 40.600 424.500 41.400 ;
        RECT 424.700 40.600 425.500 41.400 ;
        RECT 425.700 40.600 426.500 41.400 ;
        RECT 426.700 40.600 427.500 41.400 ;
        RECT 427.700 40.600 428.500 41.400 ;
        RECT 31.600 37.600 32.400 38.400 ;
        RECT 66.800 37.600 67.600 38.400 ;
        RECT 31.600 31.600 32.400 32.400 ;
        RECT 66.800 31.600 67.600 32.400 ;
        RECT 97.200 31.200 98.000 32.000 ;
        RECT 350.000 31.200 350.800 32.000 ;
        RECT 375.600 37.600 376.400 38.400 ;
        RECT 420.400 37.600 421.200 38.400 ;
        RECT 375.600 31.600 376.400 32.400 ;
        RECT 420.400 31.600 421.200 32.400 ;
        RECT 508.400 31.200 509.200 32.000 ;
        RECT 206.000 11.600 206.800 12.400 ;
        RECT 298.800 11.600 299.600 12.400 ;
        RECT 31.600 3.600 32.400 4.400 ;
        RECT 42.800 3.600 43.600 4.400 ;
        RECT 87.600 3.600 88.400 4.400 ;
        RECT 164.400 10.000 165.200 10.800 ;
        RECT 164.400 3.600 165.200 4.400 ;
        RECT 206.000 5.400 206.800 6.200 ;
        RECT 364.400 10.000 365.200 10.800 ;
        RECT 298.800 5.400 299.600 6.200 ;
        RECT 364.400 5.400 365.200 6.200 ;
        RECT 399.600 3.600 400.400 4.400 ;
        RECT 470.000 3.600 470.800 4.400 ;
        RECT 508.400 3.600 509.200 4.400 ;
        RECT 121.900 0.600 122.700 1.400 ;
        RECT 122.900 0.600 123.700 1.400 ;
        RECT 123.900 0.600 124.700 1.400 ;
        RECT 124.900 0.600 125.700 1.400 ;
        RECT 125.900 0.600 126.700 1.400 ;
        RECT 126.900 0.600 127.700 1.400 ;
        RECT 422.700 0.600 423.500 1.400 ;
        RECT 423.700 0.600 424.500 1.400 ;
        RECT 424.700 0.600 425.500 1.400 ;
        RECT 425.700 0.600 426.500 1.400 ;
        RECT 426.700 0.600 427.500 1.400 ;
        RECT 427.700 0.600 428.500 1.400 ;
      LAYER metal2 ;
        RECT 372.400 371.600 373.200 372.400 ;
        RECT 31.600 369.600 32.400 370.400 ;
        RECT 42.800 370.000 43.600 370.800 ;
        RECT 98.800 370.000 99.600 370.800 ;
        RECT 31.700 364.400 32.300 369.600 ;
        RECT 42.900 364.400 43.500 370.000 ;
        RECT 98.900 366.200 99.500 370.000 ;
        RECT 143.600 369.600 144.400 370.400 ;
        RECT 154.800 370.000 155.600 370.800 ;
        RECT 190.000 370.000 190.800 370.800 ;
        RECT 98.800 365.400 99.600 366.200 ;
        RECT 143.700 364.400 144.300 369.600 ;
        RECT 154.900 364.400 155.500 370.000 ;
        RECT 190.100 364.400 190.700 370.000 ;
        RECT 282.800 369.600 283.600 370.400 ;
        RECT 282.900 364.400 283.500 369.600 ;
        RECT 372.500 366.200 373.100 371.600 ;
        RECT 398.000 369.600 398.800 370.400 ;
        RECT 466.800 369.600 467.600 370.400 ;
        RECT 478.000 370.000 478.800 370.800 ;
        RECT 538.800 370.000 539.600 370.800 ;
        RECT 372.400 365.400 373.200 366.200 ;
        RECT 398.100 364.400 398.700 369.600 ;
        RECT 466.900 364.400 467.500 369.600 ;
        RECT 478.100 366.200 478.700 370.000 ;
        RECT 478.000 365.400 478.800 366.200 ;
        RECT 538.900 364.400 539.500 370.000 ;
        RECT 31.600 363.600 32.400 364.400 ;
        RECT 42.800 363.600 43.600 364.400 ;
        RECT 143.600 363.600 144.400 364.400 ;
        RECT 154.800 363.600 155.600 364.400 ;
        RECT 190.000 363.600 190.800 364.400 ;
        RECT 282.800 363.600 283.600 364.400 ;
        RECT 398.000 363.600 398.800 364.400 ;
        RECT 466.800 363.600 467.600 364.400 ;
        RECT 538.800 363.600 539.600 364.400 ;
        RECT 124.200 361.400 125.400 361.600 ;
        RECT 425.000 361.400 426.200 361.600 ;
        RECT 121.900 360.600 127.700 361.400 ;
        RECT 422.700 360.600 428.500 361.400 ;
        RECT 124.200 360.400 125.400 360.600 ;
        RECT 425.000 360.400 426.200 360.600 ;
        RECT 31.600 357.600 32.400 358.400 ;
        RECT 143.600 357.600 144.400 358.400 ;
        RECT 268.400 357.600 269.200 358.400 ;
        RECT 545.200 357.600 546.000 358.400 ;
        RECT 31.700 352.400 32.300 357.600 ;
        RECT 65.200 355.800 66.000 356.600 ;
        RECT 105.200 355.800 106.000 356.600 ;
        RECT 31.600 351.600 32.400 352.400 ;
        RECT 65.300 352.000 65.900 355.800 ;
        RECT 105.300 352.000 105.900 355.800 ;
        RECT 143.700 352.400 144.300 357.600 ;
        RECT 202.800 355.800 203.600 356.600 ;
        RECT 238.000 355.800 238.800 356.600 ;
        RECT 65.200 351.200 66.000 352.000 ;
        RECT 105.200 351.200 106.000 352.000 ;
        RECT 143.600 351.600 144.400 352.400 ;
        RECT 202.900 352.000 203.500 355.800 ;
        RECT 238.100 352.000 238.700 355.800 ;
        RECT 268.500 352.400 269.100 357.600 ;
        RECT 545.300 352.400 545.900 357.600 ;
        RECT 202.800 351.200 203.600 352.000 ;
        RECT 238.000 351.200 238.800 352.000 ;
        RECT 268.400 351.600 269.200 352.400 ;
        RECT 545.200 351.600 546.000 352.400 ;
        RECT 34.800 329.600 35.600 330.400 ;
        RECT 121.200 330.000 122.000 330.800 ;
        RECT 142.000 330.000 142.800 330.800 ;
        RECT 246.000 330.000 246.800 330.800 ;
        RECT 34.900 324.400 35.500 329.600 ;
        RECT 121.300 326.200 121.900 330.000 ;
        RECT 121.200 325.400 122.000 326.200 ;
        RECT 142.100 324.400 142.700 330.000 ;
        RECT 246.100 326.200 246.700 330.000 ;
        RECT 278.000 329.600 278.800 330.400 ;
        RECT 316.400 330.000 317.200 330.800 ;
        RECT 246.000 325.400 246.800 326.200 ;
        RECT 278.100 324.400 278.700 329.600 ;
        RECT 316.500 326.200 317.100 330.000 ;
        RECT 462.000 329.600 462.800 330.400 ;
        RECT 316.400 325.400 317.200 326.200 ;
        RECT 462.100 324.400 462.700 329.600 ;
        RECT 34.800 323.600 35.600 324.400 ;
        RECT 142.000 323.600 142.800 324.400 ;
        RECT 278.000 323.600 278.800 324.400 ;
        RECT 462.000 323.600 462.800 324.400 ;
        RECT 124.200 321.400 125.400 321.600 ;
        RECT 425.000 321.400 426.200 321.600 ;
        RECT 121.900 320.600 127.700 321.400 ;
        RECT 422.700 320.600 428.500 321.400 ;
        RECT 124.200 320.400 125.400 320.600 ;
        RECT 425.000 320.400 426.200 320.600 ;
        RECT 279.600 317.600 280.400 318.400 ;
        RECT 444.400 317.600 445.200 318.400 ;
        RECT 279.700 312.400 280.300 317.600 ;
        RECT 311.600 315.600 312.400 316.400 ;
        RECT 279.600 311.600 280.400 312.400 ;
        RECT 311.700 310.400 312.300 315.600 ;
        RECT 444.500 312.400 445.100 317.600 ;
        RECT 444.400 311.600 445.200 312.400 ;
        RECT 311.600 309.600 312.400 310.400 ;
        RECT 65.200 290.000 66.000 290.800 ;
        RECT 100.400 290.000 101.200 290.800 ;
        RECT 302.000 290.000 302.800 290.800 ;
        RECT 478.000 290.000 478.800 290.800 ;
        RECT 540.400 290.000 541.200 290.800 ;
        RECT 65.300 286.200 65.900 290.000 ;
        RECT 65.200 285.400 66.000 286.200 ;
        RECT 100.500 284.400 101.100 290.000 ;
        RECT 302.100 286.200 302.700 290.000 ;
        RECT 478.100 286.200 478.700 290.000 ;
        RECT 540.500 286.200 541.100 290.000 ;
        RECT 302.000 285.400 302.800 286.200 ;
        RECT 478.000 285.400 478.800 286.200 ;
        RECT 540.400 285.400 541.200 286.200 ;
        RECT 100.400 283.600 101.200 284.400 ;
        RECT 124.200 281.400 125.400 281.600 ;
        RECT 425.000 281.400 426.200 281.600 ;
        RECT 121.900 280.600 127.700 281.400 ;
        RECT 422.700 280.600 428.500 281.400 ;
        RECT 124.200 280.400 125.400 280.600 ;
        RECT 425.000 280.400 426.200 280.600 ;
        RECT 31.600 277.600 32.400 278.400 ;
        RECT 482.800 277.600 483.600 278.400 ;
        RECT 518.000 277.600 518.800 278.400 ;
        RECT 31.700 272.400 32.300 277.600 ;
        RECT 97.200 275.800 98.000 276.600 ;
        RECT 31.600 271.600 32.400 272.400 ;
        RECT 97.300 272.000 97.900 275.800 ;
        RECT 289.200 275.600 290.000 276.400 ;
        RECT 316.400 275.600 317.200 276.400 ;
        RECT 361.200 275.600 362.000 276.400 ;
        RECT 390.000 275.800 390.800 276.600 ;
        RECT 97.200 271.200 98.000 272.000 ;
        RECT 289.300 270.400 289.900 275.600 ;
        RECT 316.500 270.400 317.100 275.600 ;
        RECT 361.300 270.400 361.900 275.600 ;
        RECT 390.100 272.000 390.700 275.800 ;
        RECT 482.900 272.400 483.500 277.600 ;
        RECT 518.100 272.400 518.700 277.600 ;
        RECT 390.000 271.200 390.800 272.000 ;
        RECT 482.800 271.600 483.600 272.400 ;
        RECT 518.000 271.600 518.800 272.400 ;
        RECT 289.200 269.600 290.000 270.400 ;
        RECT 316.400 269.600 317.200 270.400 ;
        RECT 361.200 269.600 362.000 270.400 ;
        RECT 255.600 251.600 256.400 252.400 ;
        RECT 297.200 251.600 298.000 252.400 ;
        RECT 106.800 250.000 107.600 250.800 ;
        RECT 151.600 250.000 152.400 250.800 ;
        RECT 106.900 246.200 107.500 250.000 ;
        RECT 151.700 246.200 152.300 250.000 ;
        RECT 236.400 249.600 237.200 250.400 ;
        RECT 106.800 245.400 107.600 246.200 ;
        RECT 151.600 245.400 152.400 246.200 ;
        RECT 236.500 244.400 237.100 249.600 ;
        RECT 255.700 246.200 256.300 251.600 ;
        RECT 297.300 246.200 297.900 251.600 ;
        RECT 356.400 250.000 357.200 250.800 ;
        RECT 415.600 250.000 416.400 250.800 ;
        RECT 460.400 250.000 461.200 250.800 ;
        RECT 486.000 250.000 486.800 250.800 ;
        RECT 356.500 246.200 357.100 250.000 ;
        RECT 255.600 245.400 256.400 246.200 ;
        RECT 297.200 245.400 298.000 246.200 ;
        RECT 356.400 245.400 357.200 246.200 ;
        RECT 415.700 244.400 416.300 250.000 ;
        RECT 460.500 246.200 461.100 250.000 ;
        RECT 486.100 246.200 486.700 250.000 ;
        RECT 460.400 245.400 461.200 246.200 ;
        RECT 486.000 245.400 486.800 246.200 ;
        RECT 236.400 243.600 237.200 244.400 ;
        RECT 415.600 243.600 416.400 244.400 ;
        RECT 124.200 241.400 125.400 241.600 ;
        RECT 425.000 241.400 426.200 241.600 ;
        RECT 121.900 240.600 127.700 241.400 ;
        RECT 422.700 240.600 428.500 241.400 ;
        RECT 124.200 240.400 125.400 240.600 ;
        RECT 425.000 240.400 426.200 240.600 ;
        RECT 31.600 237.600 32.400 238.400 ;
        RECT 234.800 237.600 235.600 238.400 ;
        RECT 526.000 237.600 526.800 238.400 ;
        RECT 31.700 232.400 32.300 237.600 ;
        RECT 130.800 235.800 131.600 236.600 ;
        RECT 31.600 231.600 32.400 232.400 ;
        RECT 130.900 232.000 131.500 235.800 ;
        RECT 234.900 232.400 235.500 237.600 ;
        RECT 266.800 235.800 267.600 236.600 ;
        RECT 130.800 231.200 131.600 232.000 ;
        RECT 234.800 231.600 235.600 232.400 ;
        RECT 266.900 232.000 267.500 235.800 ;
        RECT 305.200 235.600 306.000 236.400 ;
        RECT 404.400 235.800 405.200 236.600 ;
        RECT 266.800 231.200 267.600 232.000 ;
        RECT 305.300 230.400 305.900 235.600 ;
        RECT 404.500 232.000 405.100 235.800 ;
        RECT 526.100 232.400 526.700 237.600 ;
        RECT 404.400 231.200 405.200 232.000 ;
        RECT 526.000 231.600 526.800 232.400 ;
        RECT 305.200 229.600 306.000 230.400 ;
        RECT 300.400 211.600 301.200 212.400 ;
        RECT 119.600 209.600 120.400 210.400 ;
        RECT 273.200 210.000 274.000 210.800 ;
        RECT 119.700 204.400 120.300 209.600 ;
        RECT 273.300 204.400 273.900 210.000 ;
        RECT 300.500 206.200 301.100 211.600 ;
        RECT 510.000 209.600 510.800 210.400 ;
        RECT 521.200 210.000 522.000 210.800 ;
        RECT 300.400 205.400 301.200 206.200 ;
        RECT 510.100 204.400 510.700 209.600 ;
        RECT 521.300 206.200 521.900 210.000 ;
        RECT 521.200 205.400 522.000 206.200 ;
        RECT 119.600 203.600 120.400 204.400 ;
        RECT 273.200 203.600 274.000 204.400 ;
        RECT 510.000 203.600 510.800 204.400 ;
        RECT 124.200 201.400 125.400 201.600 ;
        RECT 425.000 201.400 426.200 201.600 ;
        RECT 121.900 200.600 127.700 201.400 ;
        RECT 422.700 200.600 428.500 201.400 ;
        RECT 124.200 200.400 125.400 200.600 ;
        RECT 425.000 200.400 426.200 200.600 ;
        RECT 146.800 197.600 147.600 198.400 ;
        RECT 212.400 197.600 213.200 198.400 ;
        RECT 498.800 197.600 499.600 198.400 ;
        RECT 73.200 195.800 74.000 196.600 ;
        RECT 73.300 192.000 73.900 195.800 ;
        RECT 122.800 195.600 123.600 196.400 ;
        RECT 73.200 191.200 74.000 192.000 ;
        RECT 122.900 190.400 123.500 195.600 ;
        RECT 146.900 192.400 147.500 197.600 ;
        RECT 212.500 192.400 213.100 197.600 ;
        RECT 294.000 195.800 294.800 196.600 ;
        RECT 146.800 191.600 147.600 192.400 ;
        RECT 212.400 191.600 213.200 192.400 ;
        RECT 294.100 192.000 294.700 195.800 ;
        RECT 322.800 195.600 323.600 196.400 ;
        RECT 359.600 195.600 360.400 196.400 ;
        RECT 294.000 191.200 294.800 192.000 ;
        RECT 322.900 190.400 323.500 195.600 ;
        RECT 359.700 190.400 360.300 195.600 ;
        RECT 498.900 192.400 499.500 197.600 ;
        RECT 498.800 191.600 499.600 192.400 ;
        RECT 122.800 189.600 123.600 190.400 ;
        RECT 322.800 189.600 323.600 190.400 ;
        RECT 359.600 189.600 360.400 190.400 ;
        RECT 126.000 171.600 126.800 172.400 ;
        RECT 82.800 170.000 83.600 170.800 ;
        RECT 82.900 164.400 83.500 170.000 ;
        RECT 126.100 166.200 126.700 171.600 ;
        RECT 154.800 169.600 155.600 170.400 ;
        RECT 231.600 169.600 232.400 170.400 ;
        RECT 324.400 169.600 325.200 170.400 ;
        RECT 370.800 170.000 371.600 170.800 ;
        RECT 444.400 170.000 445.200 170.800 ;
        RECT 540.400 170.000 541.200 170.800 ;
        RECT 126.000 165.400 126.800 166.200 ;
        RECT 154.900 164.400 155.500 169.600 ;
        RECT 231.700 164.400 232.300 169.600 ;
        RECT 324.500 164.400 325.100 169.600 ;
        RECT 370.900 164.400 371.500 170.000 ;
        RECT 444.500 166.200 445.100 170.000 ;
        RECT 540.500 166.200 541.100 170.000 ;
        RECT 444.400 165.400 445.200 166.200 ;
        RECT 540.400 165.400 541.200 166.200 ;
        RECT 82.800 163.600 83.600 164.400 ;
        RECT 154.800 163.600 155.600 164.400 ;
        RECT 231.600 163.600 232.400 164.400 ;
        RECT 324.400 163.600 325.200 164.400 ;
        RECT 370.800 163.600 371.600 164.400 ;
        RECT 124.200 161.400 125.400 161.600 ;
        RECT 425.000 161.400 426.200 161.600 ;
        RECT 121.900 160.600 127.700 161.400 ;
        RECT 422.700 160.600 428.500 161.400 ;
        RECT 124.200 160.400 125.400 160.600 ;
        RECT 425.000 160.400 426.200 160.600 ;
        RECT 151.600 157.600 152.400 158.400 ;
        RECT 97.200 155.800 98.000 156.600 ;
        RECT 97.300 152.000 97.900 155.800 ;
        RECT 151.700 152.400 152.300 157.600 ;
        RECT 228.400 155.800 229.200 156.600 ;
        RECT 97.200 151.200 98.000 152.000 ;
        RECT 151.600 151.600 152.400 152.400 ;
        RECT 228.500 152.000 229.100 155.800 ;
        RECT 314.800 155.600 315.600 156.400 ;
        RECT 228.400 151.200 229.200 152.000 ;
        RECT 314.900 150.400 315.500 155.600 ;
        RECT 314.800 149.600 315.600 150.400 ;
        RECT 281.200 131.600 282.000 132.400 ;
        RECT 76.400 130.000 77.200 130.800 ;
        RECT 105.200 130.000 106.000 130.800 ;
        RECT 76.500 124.400 77.100 130.000 ;
        RECT 105.300 126.200 105.900 130.000 ;
        RECT 212.400 129.600 213.200 130.400 ;
        RECT 105.200 125.400 106.000 126.200 ;
        RECT 212.500 124.400 213.100 129.600 ;
        RECT 281.300 126.200 281.900 131.600 ;
        RECT 329.200 130.000 330.000 130.800 ;
        RECT 422.000 130.000 422.800 130.800 ;
        RECT 281.200 125.400 282.000 126.200 ;
        RECT 329.300 124.400 329.900 130.000 ;
        RECT 422.100 126.200 422.700 130.000 ;
        RECT 468.400 129.600 469.200 130.400 ;
        RECT 545.200 129.600 546.000 130.400 ;
        RECT 422.000 125.400 422.800 126.200 ;
        RECT 468.500 124.400 469.100 129.600 ;
        RECT 545.300 124.400 545.900 129.600 ;
        RECT 76.400 123.600 77.200 124.400 ;
        RECT 212.400 123.600 213.200 124.400 ;
        RECT 329.200 123.600 330.000 124.400 ;
        RECT 468.400 123.600 469.200 124.400 ;
        RECT 545.200 123.600 546.000 124.400 ;
        RECT 124.200 121.400 125.400 121.600 ;
        RECT 425.000 121.400 426.200 121.600 ;
        RECT 121.900 120.600 127.700 121.400 ;
        RECT 422.700 120.600 428.500 121.400 ;
        RECT 124.200 120.400 125.400 120.600 ;
        RECT 425.000 120.400 426.200 120.600 ;
        RECT 73.200 117.600 74.000 118.400 ;
        RECT 87.600 117.600 88.400 118.400 ;
        RECT 183.600 117.600 184.400 118.400 ;
        RECT 342.000 117.600 342.800 118.400 ;
        RECT 546.800 117.600 547.600 118.400 ;
        RECT 73.300 112.400 73.900 117.600 ;
        RECT 87.700 112.400 88.300 117.600 ;
        RECT 183.700 112.400 184.300 117.600 ;
        RECT 294.000 115.600 294.800 116.400 ;
        RECT 73.200 111.600 74.000 112.400 ;
        RECT 87.600 111.600 88.400 112.400 ;
        RECT 183.600 111.600 184.400 112.400 ;
        RECT 294.100 110.400 294.700 115.600 ;
        RECT 342.100 112.400 342.700 117.600 ;
        RECT 546.900 112.400 547.500 117.600 ;
        RECT 342.000 111.600 342.800 112.400 ;
        RECT 546.800 111.600 547.600 112.400 ;
        RECT 294.000 109.600 294.800 110.400 ;
        RECT 70.000 91.600 70.800 92.400 ;
        RECT 316.400 91.600 317.200 92.400 ;
        RECT 70.100 86.200 70.700 91.600 ;
        RECT 105.200 90.000 106.000 90.800 ;
        RECT 105.300 86.200 105.900 90.000 ;
        RECT 298.800 89.600 299.600 90.400 ;
        RECT 70.000 85.400 70.800 86.200 ;
        RECT 105.200 85.400 106.000 86.200 ;
        RECT 298.900 84.400 299.500 89.600 ;
        RECT 316.500 86.200 317.100 91.600 ;
        RECT 361.200 90.000 362.000 90.800 ;
        RECT 508.400 90.000 509.200 90.800 ;
        RECT 543.600 90.000 544.400 90.800 ;
        RECT 316.400 85.400 317.200 86.200 ;
        RECT 361.300 84.400 361.900 90.000 ;
        RECT 508.500 86.200 509.100 90.000 ;
        RECT 508.400 85.400 509.200 86.200 ;
        RECT 543.700 84.400 544.300 90.000 ;
        RECT 298.800 83.600 299.600 84.400 ;
        RECT 361.200 83.600 362.000 84.400 ;
        RECT 543.600 83.600 544.400 84.400 ;
        RECT 124.200 81.400 125.400 81.600 ;
        RECT 425.000 81.400 426.200 81.600 ;
        RECT 121.900 80.600 127.700 81.400 ;
        RECT 422.700 80.600 428.500 81.400 ;
        RECT 124.200 80.400 125.400 80.600 ;
        RECT 425.000 80.400 426.200 80.600 ;
        RECT 121.200 77.600 122.000 78.400 ;
        RECT 175.600 77.600 176.400 78.400 ;
        RECT 446.000 77.600 446.800 78.400 ;
        RECT 545.200 77.600 546.000 78.400 ;
        RECT 121.300 72.400 121.900 77.600 ;
        RECT 153.200 75.600 154.000 76.400 ;
        RECT 121.200 71.600 122.000 72.400 ;
        RECT 153.300 70.400 153.900 75.600 ;
        RECT 175.700 72.400 176.300 77.600 ;
        RECT 234.800 75.800 235.600 76.600 ;
        RECT 175.600 71.600 176.400 72.400 ;
        RECT 234.900 72.000 235.500 75.800 ;
        RECT 294.000 75.600 294.800 76.400 ;
        RECT 364.400 75.800 365.200 76.600 ;
        RECT 234.800 71.200 235.600 72.000 ;
        RECT 294.100 70.400 294.700 75.600 ;
        RECT 364.500 72.000 365.100 75.800 ;
        RECT 446.100 72.400 446.700 77.600 ;
        RECT 545.300 72.400 545.900 77.600 ;
        RECT 364.400 71.200 365.200 72.000 ;
        RECT 446.000 71.600 446.800 72.400 ;
        RECT 545.200 71.600 546.000 72.400 ;
        RECT 153.200 69.600 154.000 70.400 ;
        RECT 294.000 69.600 294.800 70.400 ;
        RECT 114.800 51.600 115.600 52.400 ;
        RECT 201.200 51.600 202.000 52.400 ;
        RECT 244.400 51.600 245.200 52.400 ;
        RECT 305.200 51.600 306.000 52.400 ;
        RECT 47.600 50.000 48.400 50.800 ;
        RECT 47.700 44.400 48.300 50.000 ;
        RECT 114.900 46.200 115.500 51.600 ;
        RECT 201.300 46.200 201.900 51.600 ;
        RECT 244.500 46.200 245.100 51.600 ;
        RECT 305.300 46.200 305.900 51.600 ;
        RECT 326.000 50.000 326.800 50.800 ;
        RECT 380.400 50.000 381.200 50.800 ;
        RECT 468.400 50.000 469.200 50.800 ;
        RECT 540.400 50.000 541.200 50.800 ;
        RECT 326.100 46.200 326.700 50.000 ;
        RECT 380.500 46.200 381.100 50.000 ;
        RECT 468.500 46.200 469.100 50.000 ;
        RECT 540.500 46.200 541.100 50.000 ;
        RECT 114.800 45.400 115.600 46.200 ;
        RECT 201.200 45.400 202.000 46.200 ;
        RECT 244.400 45.400 245.200 46.200 ;
        RECT 305.200 45.400 306.000 46.200 ;
        RECT 326.000 45.400 326.800 46.200 ;
        RECT 380.400 45.400 381.200 46.200 ;
        RECT 468.400 45.400 469.200 46.200 ;
        RECT 540.400 45.400 541.200 46.200 ;
        RECT 47.600 43.600 48.400 44.400 ;
        RECT 124.200 41.400 125.400 41.600 ;
        RECT 425.000 41.400 426.200 41.600 ;
        RECT 121.900 40.600 127.700 41.400 ;
        RECT 422.700 40.600 428.500 41.400 ;
        RECT 124.200 40.400 125.400 40.600 ;
        RECT 425.000 40.400 426.200 40.600 ;
        RECT 31.600 37.600 32.400 38.400 ;
        RECT 66.800 37.600 67.600 38.400 ;
        RECT 375.600 37.600 376.400 38.400 ;
        RECT 420.400 37.600 421.200 38.400 ;
        RECT 31.700 32.400 32.300 37.600 ;
        RECT 66.900 32.400 67.500 37.600 ;
        RECT 97.200 35.800 98.000 36.600 ;
        RECT 31.600 31.600 32.400 32.400 ;
        RECT 66.800 31.600 67.600 32.400 ;
        RECT 97.300 32.000 97.900 35.800 ;
        RECT 153.200 35.600 154.000 36.400 ;
        RECT 188.400 35.600 189.200 36.400 ;
        RECT 250.800 35.600 251.600 36.400 ;
        RECT 308.400 35.600 309.200 36.400 ;
        RECT 350.000 35.800 350.800 36.600 ;
        RECT 97.200 31.200 98.000 32.000 ;
        RECT 153.300 30.400 153.900 35.600 ;
        RECT 188.500 30.400 189.100 35.600 ;
        RECT 250.900 30.400 251.500 35.600 ;
        RECT 308.500 30.400 309.100 35.600 ;
        RECT 350.100 32.000 350.700 35.800 ;
        RECT 375.700 32.400 376.300 37.600 ;
        RECT 420.500 32.400 421.100 37.600 ;
        RECT 508.400 35.800 509.200 36.600 ;
        RECT 350.000 31.200 350.800 32.000 ;
        RECT 375.600 31.600 376.400 32.400 ;
        RECT 420.400 31.600 421.200 32.400 ;
        RECT 508.500 32.000 509.100 35.800 ;
        RECT 508.400 31.200 509.200 32.000 ;
        RECT 153.200 29.600 154.000 30.400 ;
        RECT 188.400 29.600 189.200 30.400 ;
        RECT 250.800 29.600 251.600 30.400 ;
        RECT 308.400 29.600 309.200 30.400 ;
        RECT 206.000 11.600 206.800 12.400 ;
        RECT 298.800 11.600 299.600 12.400 ;
        RECT 31.600 9.600 32.400 10.400 ;
        RECT 42.800 10.000 43.600 10.800 ;
        RECT 31.700 4.400 32.300 9.600 ;
        RECT 42.900 4.400 43.500 10.000 ;
        RECT 87.600 9.600 88.400 10.400 ;
        RECT 164.400 10.000 165.200 10.800 ;
        RECT 87.700 4.400 88.300 9.600 ;
        RECT 164.500 4.400 165.100 10.000 ;
        RECT 206.100 6.200 206.700 11.600 ;
        RECT 298.900 6.200 299.500 11.600 ;
        RECT 364.400 10.000 365.200 10.800 ;
        RECT 364.500 6.200 365.100 10.000 ;
        RECT 399.600 9.600 400.400 10.400 ;
        RECT 470.000 9.600 470.800 10.400 ;
        RECT 508.400 9.600 509.200 10.400 ;
        RECT 206.000 5.400 206.800 6.200 ;
        RECT 298.800 5.400 299.600 6.200 ;
        RECT 364.400 5.400 365.200 6.200 ;
        RECT 399.700 4.400 400.300 9.600 ;
        RECT 470.100 4.400 470.700 9.600 ;
        RECT 508.500 4.400 509.100 9.600 ;
        RECT 31.600 3.600 32.400 4.400 ;
        RECT 42.800 3.600 43.600 4.400 ;
        RECT 87.600 3.600 88.400 4.400 ;
        RECT 164.400 3.600 165.200 4.400 ;
        RECT 399.600 3.600 400.400 4.400 ;
        RECT 470.000 3.600 470.800 4.400 ;
        RECT 508.400 3.600 509.200 4.400 ;
        RECT 124.200 1.400 125.400 1.600 ;
        RECT 425.000 1.400 426.200 1.600 ;
        RECT 121.900 0.600 127.700 1.400 ;
        RECT 422.700 0.600 428.500 1.400 ;
        RECT 124.200 0.400 125.400 0.600 ;
        RECT 425.000 0.400 426.200 0.600 ;
      LAYER via2 ;
        RECT 122.900 360.600 123.700 361.400 ;
        RECT 123.900 360.600 124.700 361.400 ;
        RECT 124.900 360.600 125.700 361.400 ;
        RECT 125.900 360.600 126.700 361.400 ;
        RECT 126.900 360.600 127.700 361.400 ;
        RECT 423.700 360.600 424.500 361.400 ;
        RECT 424.700 360.600 425.500 361.400 ;
        RECT 425.700 360.600 426.500 361.400 ;
        RECT 426.700 360.600 427.500 361.400 ;
        RECT 427.700 360.600 428.500 361.400 ;
        RECT 122.900 320.600 123.700 321.400 ;
        RECT 123.900 320.600 124.700 321.400 ;
        RECT 124.900 320.600 125.700 321.400 ;
        RECT 125.900 320.600 126.700 321.400 ;
        RECT 126.900 320.600 127.700 321.400 ;
        RECT 423.700 320.600 424.500 321.400 ;
        RECT 424.700 320.600 425.500 321.400 ;
        RECT 425.700 320.600 426.500 321.400 ;
        RECT 426.700 320.600 427.500 321.400 ;
        RECT 427.700 320.600 428.500 321.400 ;
        RECT 122.900 280.600 123.700 281.400 ;
        RECT 123.900 280.600 124.700 281.400 ;
        RECT 124.900 280.600 125.700 281.400 ;
        RECT 125.900 280.600 126.700 281.400 ;
        RECT 126.900 280.600 127.700 281.400 ;
        RECT 423.700 280.600 424.500 281.400 ;
        RECT 424.700 280.600 425.500 281.400 ;
        RECT 425.700 280.600 426.500 281.400 ;
        RECT 426.700 280.600 427.500 281.400 ;
        RECT 427.700 280.600 428.500 281.400 ;
        RECT 122.900 240.600 123.700 241.400 ;
        RECT 123.900 240.600 124.700 241.400 ;
        RECT 124.900 240.600 125.700 241.400 ;
        RECT 125.900 240.600 126.700 241.400 ;
        RECT 126.900 240.600 127.700 241.400 ;
        RECT 423.700 240.600 424.500 241.400 ;
        RECT 424.700 240.600 425.500 241.400 ;
        RECT 425.700 240.600 426.500 241.400 ;
        RECT 426.700 240.600 427.500 241.400 ;
        RECT 427.700 240.600 428.500 241.400 ;
        RECT 122.900 200.600 123.700 201.400 ;
        RECT 123.900 200.600 124.700 201.400 ;
        RECT 124.900 200.600 125.700 201.400 ;
        RECT 125.900 200.600 126.700 201.400 ;
        RECT 126.900 200.600 127.700 201.400 ;
        RECT 423.700 200.600 424.500 201.400 ;
        RECT 424.700 200.600 425.500 201.400 ;
        RECT 425.700 200.600 426.500 201.400 ;
        RECT 426.700 200.600 427.500 201.400 ;
        RECT 427.700 200.600 428.500 201.400 ;
        RECT 122.900 160.600 123.700 161.400 ;
        RECT 123.900 160.600 124.700 161.400 ;
        RECT 124.900 160.600 125.700 161.400 ;
        RECT 125.900 160.600 126.700 161.400 ;
        RECT 126.900 160.600 127.700 161.400 ;
        RECT 423.700 160.600 424.500 161.400 ;
        RECT 424.700 160.600 425.500 161.400 ;
        RECT 425.700 160.600 426.500 161.400 ;
        RECT 426.700 160.600 427.500 161.400 ;
        RECT 427.700 160.600 428.500 161.400 ;
        RECT 122.900 120.600 123.700 121.400 ;
        RECT 123.900 120.600 124.700 121.400 ;
        RECT 124.900 120.600 125.700 121.400 ;
        RECT 125.900 120.600 126.700 121.400 ;
        RECT 126.900 120.600 127.700 121.400 ;
        RECT 423.700 120.600 424.500 121.400 ;
        RECT 424.700 120.600 425.500 121.400 ;
        RECT 425.700 120.600 426.500 121.400 ;
        RECT 426.700 120.600 427.500 121.400 ;
        RECT 427.700 120.600 428.500 121.400 ;
        RECT 122.900 80.600 123.700 81.400 ;
        RECT 123.900 80.600 124.700 81.400 ;
        RECT 124.900 80.600 125.700 81.400 ;
        RECT 125.900 80.600 126.700 81.400 ;
        RECT 126.900 80.600 127.700 81.400 ;
        RECT 423.700 80.600 424.500 81.400 ;
        RECT 424.700 80.600 425.500 81.400 ;
        RECT 425.700 80.600 426.500 81.400 ;
        RECT 426.700 80.600 427.500 81.400 ;
        RECT 427.700 80.600 428.500 81.400 ;
        RECT 122.900 40.600 123.700 41.400 ;
        RECT 123.900 40.600 124.700 41.400 ;
        RECT 124.900 40.600 125.700 41.400 ;
        RECT 125.900 40.600 126.700 41.400 ;
        RECT 126.900 40.600 127.700 41.400 ;
        RECT 423.700 40.600 424.500 41.400 ;
        RECT 424.700 40.600 425.500 41.400 ;
        RECT 425.700 40.600 426.500 41.400 ;
        RECT 426.700 40.600 427.500 41.400 ;
        RECT 427.700 40.600 428.500 41.400 ;
        RECT 122.900 0.600 123.700 1.400 ;
        RECT 123.900 0.600 124.700 1.400 ;
        RECT 124.900 0.600 125.700 1.400 ;
        RECT 125.900 0.600 126.700 1.400 ;
        RECT 126.900 0.600 127.700 1.400 ;
        RECT 423.700 0.600 424.500 1.400 ;
        RECT 424.700 0.600 425.500 1.400 ;
        RECT 425.700 0.600 426.500 1.400 ;
        RECT 426.700 0.600 427.500 1.400 ;
        RECT 427.700 0.600 428.500 1.400 ;
      LAYER metal3 ;
        RECT 121.800 360.400 127.800 361.600 ;
        RECT 422.600 360.400 428.600 361.600 ;
        RECT 121.800 320.400 127.800 321.600 ;
        RECT 422.600 320.400 428.600 321.600 ;
        RECT 121.800 280.400 127.800 281.600 ;
        RECT 422.600 280.400 428.600 281.600 ;
        RECT 121.800 240.400 127.800 241.600 ;
        RECT 422.600 240.400 428.600 241.600 ;
        RECT 121.800 200.400 127.800 201.600 ;
        RECT 422.600 200.400 428.600 201.600 ;
        RECT 121.800 160.400 127.800 161.600 ;
        RECT 422.600 160.400 428.600 161.600 ;
        RECT 121.800 120.400 127.800 121.600 ;
        RECT 422.600 120.400 428.600 121.600 ;
        RECT 121.800 80.400 127.800 81.600 ;
        RECT 422.600 80.400 428.600 81.600 ;
        RECT 121.800 40.400 127.800 41.600 ;
        RECT 422.600 40.400 428.600 41.600 ;
        RECT 121.800 0.400 127.800 1.600 ;
        RECT 422.600 0.400 428.600 1.600 ;
      LAYER via3 ;
        RECT 122.000 360.600 122.800 361.400 ;
        RECT 123.200 360.600 124.000 361.400 ;
        RECT 124.400 360.600 125.200 361.400 ;
        RECT 125.600 360.600 126.400 361.400 ;
        RECT 126.800 360.600 127.600 361.400 ;
        RECT 422.800 360.600 423.600 361.400 ;
        RECT 424.000 360.600 424.800 361.400 ;
        RECT 425.200 360.600 426.000 361.400 ;
        RECT 426.400 360.600 427.200 361.400 ;
        RECT 427.600 360.600 428.400 361.400 ;
        RECT 122.000 320.600 122.800 321.400 ;
        RECT 123.200 320.600 124.000 321.400 ;
        RECT 124.400 320.600 125.200 321.400 ;
        RECT 125.600 320.600 126.400 321.400 ;
        RECT 126.800 320.600 127.600 321.400 ;
        RECT 422.800 320.600 423.600 321.400 ;
        RECT 424.000 320.600 424.800 321.400 ;
        RECT 425.200 320.600 426.000 321.400 ;
        RECT 426.400 320.600 427.200 321.400 ;
        RECT 427.600 320.600 428.400 321.400 ;
        RECT 122.000 280.600 122.800 281.400 ;
        RECT 123.200 280.600 124.000 281.400 ;
        RECT 124.400 280.600 125.200 281.400 ;
        RECT 125.600 280.600 126.400 281.400 ;
        RECT 126.800 280.600 127.600 281.400 ;
        RECT 422.800 280.600 423.600 281.400 ;
        RECT 424.000 280.600 424.800 281.400 ;
        RECT 425.200 280.600 426.000 281.400 ;
        RECT 426.400 280.600 427.200 281.400 ;
        RECT 427.600 280.600 428.400 281.400 ;
        RECT 122.000 240.600 122.800 241.400 ;
        RECT 123.200 240.600 124.000 241.400 ;
        RECT 124.400 240.600 125.200 241.400 ;
        RECT 125.600 240.600 126.400 241.400 ;
        RECT 126.800 240.600 127.600 241.400 ;
        RECT 422.800 240.600 423.600 241.400 ;
        RECT 424.000 240.600 424.800 241.400 ;
        RECT 425.200 240.600 426.000 241.400 ;
        RECT 426.400 240.600 427.200 241.400 ;
        RECT 427.600 240.600 428.400 241.400 ;
        RECT 122.000 200.600 122.800 201.400 ;
        RECT 123.200 200.600 124.000 201.400 ;
        RECT 124.400 200.600 125.200 201.400 ;
        RECT 125.600 200.600 126.400 201.400 ;
        RECT 126.800 200.600 127.600 201.400 ;
        RECT 422.800 200.600 423.600 201.400 ;
        RECT 424.000 200.600 424.800 201.400 ;
        RECT 425.200 200.600 426.000 201.400 ;
        RECT 426.400 200.600 427.200 201.400 ;
        RECT 427.600 200.600 428.400 201.400 ;
        RECT 122.000 160.600 122.800 161.400 ;
        RECT 123.200 160.600 124.000 161.400 ;
        RECT 124.400 160.600 125.200 161.400 ;
        RECT 125.600 160.600 126.400 161.400 ;
        RECT 126.800 160.600 127.600 161.400 ;
        RECT 422.800 160.600 423.600 161.400 ;
        RECT 424.000 160.600 424.800 161.400 ;
        RECT 425.200 160.600 426.000 161.400 ;
        RECT 426.400 160.600 427.200 161.400 ;
        RECT 427.600 160.600 428.400 161.400 ;
        RECT 122.000 120.600 122.800 121.400 ;
        RECT 123.200 120.600 124.000 121.400 ;
        RECT 124.400 120.600 125.200 121.400 ;
        RECT 125.600 120.600 126.400 121.400 ;
        RECT 126.800 120.600 127.600 121.400 ;
        RECT 422.800 120.600 423.600 121.400 ;
        RECT 424.000 120.600 424.800 121.400 ;
        RECT 425.200 120.600 426.000 121.400 ;
        RECT 426.400 120.600 427.200 121.400 ;
        RECT 427.600 120.600 428.400 121.400 ;
        RECT 122.000 80.600 122.800 81.400 ;
        RECT 123.200 80.600 124.000 81.400 ;
        RECT 124.400 80.600 125.200 81.400 ;
        RECT 125.600 80.600 126.400 81.400 ;
        RECT 126.800 80.600 127.600 81.400 ;
        RECT 422.800 80.600 423.600 81.400 ;
        RECT 424.000 80.600 424.800 81.400 ;
        RECT 425.200 80.600 426.000 81.400 ;
        RECT 426.400 80.600 427.200 81.400 ;
        RECT 427.600 80.600 428.400 81.400 ;
        RECT 122.000 40.600 122.800 41.400 ;
        RECT 123.200 40.600 124.000 41.400 ;
        RECT 124.400 40.600 125.200 41.400 ;
        RECT 125.600 40.600 126.400 41.400 ;
        RECT 126.800 40.600 127.600 41.400 ;
        RECT 422.800 40.600 423.600 41.400 ;
        RECT 424.000 40.600 424.800 41.400 ;
        RECT 425.200 40.600 426.000 41.400 ;
        RECT 426.400 40.600 427.200 41.400 ;
        RECT 427.600 40.600 428.400 41.400 ;
        RECT 122.000 0.600 122.800 1.400 ;
        RECT 123.200 0.600 124.000 1.400 ;
        RECT 124.400 0.600 125.200 1.400 ;
        RECT 125.600 0.600 126.400 1.400 ;
        RECT 126.800 0.600 127.600 1.400 ;
        RECT 422.800 0.600 423.600 1.400 ;
        RECT 424.000 0.600 424.800 1.400 ;
        RECT 425.200 0.600 426.000 1.400 ;
        RECT 426.400 0.600 427.200 1.400 ;
        RECT 427.600 0.600 428.400 1.400 ;
      LAYER metal4 ;
        RECT 121.600 -1.000 128.000 381.600 ;
        RECT 422.400 -1.000 428.800 381.600 ;
    END
  END vdd
  PIN arst_i
    PORT
      LAYER metal1 ;
        RECT 174.000 331.600 174.800 333.200 ;
        RECT 206.000 331.600 206.800 333.200 ;
        RECT 433.200 291.600 434.000 293.200 ;
        RECT 185.200 228.800 186.000 230.400 ;
        RECT 364.400 228.800 365.200 230.400 ;
        RECT 450.800 188.800 451.600 190.400 ;
        RECT 175.600 91.600 176.400 93.200 ;
        RECT 180.400 91.600 181.200 93.200 ;
        RECT 422.000 91.600 422.800 93.200 ;
        RECT 449.200 92.300 450.000 92.400 ;
        RECT 450.800 92.300 451.600 93.200 ;
        RECT 449.200 91.700 451.600 92.300 ;
        RECT 449.200 91.600 450.000 91.700 ;
        RECT 450.800 91.600 451.600 91.700 ;
        RECT 170.800 68.800 171.600 70.400 ;
      LAYER via1 ;
        RECT 185.200 229.600 186.000 230.400 ;
        RECT 364.400 229.600 365.200 230.400 ;
        RECT 450.800 189.600 451.600 190.400 ;
        RECT 170.800 69.600 171.600 70.400 ;
      LAYER metal2 ;
        RECT 206.100 382.400 206.700 386.300 ;
        RECT 206.000 381.600 206.800 382.400 ;
        RECT 174.000 331.600 174.800 332.400 ;
        RECT 206.000 331.600 206.800 332.400 ;
        RECT 433.200 291.600 434.000 292.400 ;
        RECT 185.200 239.600 186.000 240.400 ;
        RECT 185.300 230.400 185.900 239.600 ;
        RECT 364.400 237.600 365.200 238.400 ;
        RECT 364.500 230.400 365.100 237.600 ;
        RECT 185.200 229.600 186.000 230.400 ;
        RECT 364.400 229.600 365.200 230.400 ;
        RECT 450.800 225.600 451.600 226.400 ;
        RECT 450.900 190.400 451.500 225.600 ;
        RECT 450.800 189.600 451.600 190.400 ;
        RECT 450.900 150.400 451.500 189.600 ;
        RECT 450.800 149.600 451.600 150.400 ;
        RECT 170.800 91.600 171.600 92.400 ;
        RECT 175.600 91.600 176.400 92.400 ;
        RECT 180.400 91.600 181.200 92.400 ;
        RECT 422.000 91.600 422.800 92.400 ;
        RECT 449.200 91.600 450.000 92.400 ;
        RECT 170.900 70.400 171.500 91.600 ;
        RECT 170.800 69.600 171.600 70.400 ;
      LAYER metal3 ;
        RECT 206.000 382.300 206.800 382.400 ;
        RECT 209.200 382.300 210.000 382.400 ;
        RECT 206.000 381.700 210.000 382.300 ;
        RECT 206.000 381.600 206.800 381.700 ;
        RECT 209.200 381.600 210.000 381.700 ;
        RECT 174.000 332.300 174.800 332.400 ;
        RECT 206.000 332.300 206.800 332.400 ;
        RECT 209.200 332.300 210.000 332.400 ;
        RECT 174.000 331.700 210.000 332.300 ;
        RECT 174.000 331.600 174.800 331.700 ;
        RECT 206.000 331.600 206.800 331.700 ;
        RECT 209.200 331.600 210.000 331.700 ;
        RECT 433.200 292.300 434.000 292.400 ;
        RECT 442.800 292.300 443.600 292.400 ;
        RECT 433.200 291.700 443.600 292.300 ;
        RECT 433.200 291.600 434.000 291.700 ;
        RECT 442.800 291.600 443.600 291.700 ;
        RECT 366.000 248.300 366.800 248.400 ;
        RECT 442.800 248.300 443.600 248.400 ;
        RECT 366.000 247.700 443.600 248.300 ;
        RECT 366.000 247.600 366.800 247.700 ;
        RECT 442.800 247.600 443.600 247.700 ;
        RECT 170.800 240.300 171.600 240.400 ;
        RECT 185.200 240.300 186.000 240.400 ;
        RECT 209.200 240.300 210.000 240.400 ;
        RECT 170.800 239.700 307.500 240.300 ;
        RECT 170.800 239.600 171.600 239.700 ;
        RECT 185.200 239.600 186.000 239.700 ;
        RECT 209.200 239.600 210.000 239.700 ;
        RECT 306.900 238.300 307.500 239.700 ;
        RECT 364.400 238.300 365.200 238.400 ;
        RECT 366.000 238.300 366.800 238.400 ;
        RECT 306.900 237.700 366.800 238.300 ;
        RECT 364.400 237.600 365.200 237.700 ;
        RECT 366.000 237.600 366.800 237.700 ;
        RECT 442.800 226.300 443.600 226.400 ;
        RECT 450.800 226.300 451.600 226.400 ;
        RECT 442.800 225.700 451.600 226.300 ;
        RECT 442.800 225.600 443.600 225.700 ;
        RECT 450.800 225.600 451.600 225.700 ;
        RECT 449.200 150.300 450.000 150.400 ;
        RECT 450.800 150.300 451.600 150.400 ;
        RECT 449.200 149.700 451.600 150.300 ;
        RECT 449.200 149.600 450.000 149.700 ;
        RECT 450.800 149.600 451.600 149.700 ;
        RECT 170.800 92.300 171.600 92.400 ;
        RECT 175.600 92.300 176.400 92.400 ;
        RECT 180.400 92.300 181.200 92.400 ;
        RECT 170.800 91.700 181.200 92.300 ;
        RECT 170.800 91.600 171.600 91.700 ;
        RECT 175.600 91.600 176.400 91.700 ;
        RECT 180.400 91.600 181.200 91.700 ;
        RECT 422.000 92.300 422.800 92.400 ;
        RECT 449.200 92.300 450.000 92.400 ;
        RECT 422.000 91.700 450.000 92.300 ;
        RECT 422.000 91.600 422.800 91.700 ;
        RECT 449.200 91.600 450.000 91.700 ;
      LAYER metal4 ;
        RECT 170.600 91.400 171.800 240.600 ;
        RECT 209.000 239.400 210.200 382.600 ;
        RECT 365.800 237.400 367.000 248.600 ;
        RECT 442.600 225.400 443.800 292.600 ;
        RECT 449.000 91.400 450.200 150.600 ;
    END
  END arst_i
  PIN scl_pad_i
    PORT
      LAYER metal1 ;
        RECT 326.400 13.800 327.200 14.000 ;
        RECT 326.200 13.200 327.200 13.800 ;
        RECT 326.200 12.400 326.800 13.200 ;
        RECT 326.000 11.600 326.800 12.400 ;
      LAYER metal2 ;
        RECT 326.000 11.600 326.800 12.400 ;
        RECT 326.100 4.400 326.700 11.600 ;
        RECT 326.000 3.600 326.800 4.400 ;
        RECT 329.200 3.600 330.000 4.400 ;
        RECT 329.300 -2.300 329.900 3.600 ;
      LAYER metal3 ;
        RECT 326.000 4.300 326.800 4.400 ;
        RECT 329.200 4.300 330.000 4.400 ;
        RECT 326.000 3.700 330.000 4.300 ;
        RECT 326.000 3.600 326.800 3.700 ;
        RECT 329.200 3.600 330.000 3.700 ;
    END
  END scl_pad_i
  PIN scl_pad_o
    PORT
      LAYER metal1 ;
        RECT 172.400 12.400 173.200 19.800 ;
        RECT 172.400 10.200 173.000 12.400 ;
        RECT 172.400 2.200 173.200 10.200 ;
      LAYER via1 ;
        RECT 172.400 3.600 173.200 4.400 ;
      LAYER metal2 ;
        RECT 172.400 3.600 173.200 4.400 ;
        RECT 172.500 -1.700 173.100 3.600 ;
        RECT 172.500 -2.300 174.700 -1.700 ;
    END
  END scl_pad_o
  PIN scl_padoen_o
    PORT
      LAYER metal1 ;
        RECT 1.200 151.800 2.000 159.800 ;
        RECT 1.200 149.600 1.800 151.800 ;
        RECT 1.200 142.200 2.000 149.600 ;
      LAYER via1 ;
        RECT 1.200 147.600 2.000 148.400 ;
      LAYER metal2 ;
        RECT 1.200 149.600 2.000 150.400 ;
        RECT 1.300 148.400 1.900 149.600 ;
        RECT 1.200 147.600 2.000 148.400 ;
      LAYER metal3 ;
        RECT 1.200 150.300 2.000 150.400 ;
        RECT -3.500 149.700 2.000 150.300 ;
        RECT 1.200 149.600 2.000 149.700 ;
    END
  END scl_padoen_o
  PIN sda_pad_i
    PORT
      LAYER metal1 ;
        RECT 74.400 13.800 75.200 14.000 ;
        RECT 74.400 13.200 75.400 13.800 ;
        RECT 74.800 12.400 75.400 13.200 ;
        RECT 74.800 11.600 75.600 12.400 ;
      LAYER metal2 ;
        RECT 74.800 11.600 75.600 12.400 ;
        RECT 74.900 -1.700 75.500 11.600 ;
        RECT 74.900 -2.300 77.100 -1.700 ;
    END
  END sda_pad_i
  PIN sda_pad_o
    PORT
      LAYER metal1 ;
        RECT 180.400 12.400 181.200 19.800 ;
        RECT 180.600 10.200 181.200 12.400 ;
        RECT 180.400 2.200 181.200 10.200 ;
      LAYER via1 ;
        RECT 180.400 3.600 181.200 4.400 ;
      LAYER metal2 ;
        RECT 180.400 3.600 181.200 4.400 ;
        RECT 180.500 -1.700 181.100 3.600 ;
        RECT 178.900 -2.300 181.100 -1.700 ;
    END
  END sda_pad_o
  PIN sda_padoen_o
    PORT
      LAYER metal1 ;
        RECT 71.600 31.800 72.400 39.800 ;
        RECT 71.600 29.600 72.200 31.800 ;
        RECT 71.600 22.200 72.400 29.600 ;
      LAYER via1 ;
        RECT 71.600 23.600 72.400 24.400 ;
      LAYER metal2 ;
        RECT 71.600 23.600 72.400 24.400 ;
        RECT 71.700 -1.700 72.300 23.600 ;
        RECT 71.700 -2.300 73.900 -1.700 ;
    END
  END sda_padoen_o
  PIN wb_ack_o
    PORT
      LAYER metal1 ;
        RECT 550.000 238.300 550.800 239.800 ;
        RECT 551.600 238.300 552.400 238.400 ;
        RECT 550.000 237.700 552.400 238.300 ;
        RECT 550.000 231.800 550.800 237.700 ;
        RECT 551.600 237.600 552.400 237.700 ;
        RECT 550.200 229.600 550.800 231.800 ;
        RECT 550.000 222.200 550.800 229.600 ;
      LAYER metal2 ;
        RECT 551.600 239.600 552.400 240.400 ;
        RECT 551.700 238.400 552.300 239.600 ;
        RECT 551.600 237.600 552.400 238.400 ;
      LAYER metal3 ;
        RECT 551.600 240.300 552.400 240.400 ;
        RECT 551.600 239.700 555.500 240.300 ;
        RECT 551.600 239.600 552.400 239.700 ;
    END
  END wb_ack_o
  PIN wb_adr_i[2]
    PORT
      LAYER metal1 ;
        RECT 449.200 190.800 450.000 192.400 ;
        RECT 457.200 173.600 458.000 175.200 ;
        RECT 494.800 171.600 496.400 172.400 ;
        RECT 482.800 169.600 483.600 171.200 ;
        RECT 462.000 149.600 463.600 150.400 ;
        RECT 470.000 147.600 471.600 148.400 ;
      LAYER via1 ;
        RECT 449.200 191.600 450.000 192.400 ;
        RECT 495.600 171.600 496.400 172.400 ;
      LAYER metal2 ;
        RECT 449.200 191.600 450.000 192.400 ;
        RECT 449.300 180.400 449.900 191.600 ;
        RECT 449.200 179.600 450.000 180.400 ;
        RECT 457.200 179.600 458.000 180.400 ;
        RECT 457.300 174.400 457.900 179.600 ;
        RECT 457.200 173.600 458.000 174.400 ;
        RECT 457.300 170.400 457.900 173.600 ;
        RECT 495.600 171.600 496.400 172.400 ;
        RECT 495.700 170.400 496.300 171.600 ;
        RECT 457.200 169.600 458.000 170.400 ;
        RECT 470.000 169.600 470.800 170.400 ;
        RECT 482.800 169.600 483.600 170.400 ;
        RECT 495.600 169.600 496.400 170.400 ;
        RECT 470.100 152.400 470.700 169.600 ;
        RECT 462.000 151.600 462.800 152.400 ;
        RECT 470.000 151.600 470.800 152.400 ;
        RECT 462.100 150.400 462.700 151.600 ;
        RECT 462.000 149.600 462.800 150.400 ;
        RECT 470.100 148.400 470.700 151.600 ;
        RECT 470.000 147.600 470.800 148.400 ;
      LAYER metal3 ;
        RECT 449.200 180.300 450.000 180.400 ;
        RECT 457.200 180.300 458.000 180.400 ;
        RECT 449.200 179.700 458.000 180.300 ;
        RECT 449.200 179.600 450.000 179.700 ;
        RECT 457.200 179.600 458.000 179.700 ;
        RECT 532.400 176.300 533.200 176.400 ;
        RECT 532.400 175.700 555.500 176.300 ;
        RECT 532.400 175.600 533.200 175.700 ;
        RECT 457.200 170.300 458.000 170.400 ;
        RECT 470.000 170.300 470.800 170.400 ;
        RECT 482.800 170.300 483.600 170.400 ;
        RECT 495.600 170.300 496.400 170.400 ;
        RECT 532.400 170.300 533.200 170.400 ;
        RECT 457.200 169.700 533.200 170.300 ;
        RECT 457.200 169.600 458.000 169.700 ;
        RECT 470.000 169.600 470.800 169.700 ;
        RECT 482.800 169.600 483.600 169.700 ;
        RECT 495.600 169.600 496.400 169.700 ;
        RECT 532.400 169.600 533.200 169.700 ;
        RECT 462.000 152.300 462.800 152.400 ;
        RECT 470.000 152.300 470.800 152.400 ;
        RECT 462.000 151.700 470.800 152.300 ;
        RECT 462.000 151.600 462.800 151.700 ;
        RECT 470.000 151.600 470.800 151.700 ;
      LAYER metal4 ;
        RECT 532.200 169.400 533.400 176.600 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[1]
    PORT
      LAYER metal1 ;
        RECT 490.800 175.600 491.600 177.200 ;
        RECT 462.000 170.800 462.800 172.400 ;
        RECT 475.600 171.600 477.200 172.400 ;
        RECT 458.800 152.300 459.600 152.400 ;
        RECT 460.400 152.300 461.200 152.400 ;
        RECT 458.800 151.700 461.200 152.300 ;
        RECT 458.800 150.800 459.600 151.700 ;
        RECT 460.400 150.800 461.200 151.700 ;
        RECT 468.400 145.600 470.200 146.400 ;
      LAYER via1 ;
        RECT 462.000 171.600 462.800 172.400 ;
        RECT 476.400 171.600 477.200 172.400 ;
        RECT 460.400 151.600 461.200 152.400 ;
      LAYER metal2 ;
        RECT 490.800 179.600 491.600 180.400 ;
        RECT 490.900 176.400 491.500 179.600 ;
        RECT 490.800 175.600 491.600 176.400 ;
        RECT 462.000 171.600 462.800 172.400 ;
        RECT 476.400 171.600 477.200 172.400 ;
        RECT 462.100 164.400 462.700 171.600 ;
        RECT 476.500 166.400 477.100 171.600 ;
        RECT 490.900 166.400 491.500 175.600 ;
        RECT 476.400 165.600 477.200 166.400 ;
        RECT 490.800 165.600 491.600 166.400 ;
        RECT 462.000 164.300 462.800 164.400 ;
        RECT 460.500 163.700 462.800 164.300 ;
        RECT 460.500 152.400 461.100 163.700 ;
        RECT 462.000 163.600 462.800 163.700 ;
        RECT 468.400 163.600 469.200 164.400 ;
        RECT 460.400 151.600 461.200 152.400 ;
        RECT 468.500 146.400 469.100 163.600 ;
        RECT 468.400 145.600 469.200 146.400 ;
      LAYER metal3 ;
        RECT 490.800 180.300 491.600 180.400 ;
        RECT 490.800 179.700 537.900 180.300 ;
        RECT 490.800 179.600 491.600 179.700 ;
        RECT 537.300 178.300 537.900 179.700 ;
        RECT 554.900 178.300 555.500 180.300 ;
        RECT 537.300 177.700 555.500 178.300 ;
        RECT 476.400 166.300 477.200 166.400 ;
        RECT 490.800 166.300 491.600 166.400 ;
        RECT 476.400 165.700 491.600 166.300 ;
        RECT 476.400 165.600 477.200 165.700 ;
        RECT 490.800 165.600 491.600 165.700 ;
        RECT 462.000 164.300 462.800 164.400 ;
        RECT 468.400 164.300 469.200 164.400 ;
        RECT 476.500 164.300 477.100 165.600 ;
        RECT 462.000 163.700 477.100 164.300 ;
        RECT 462.000 163.600 462.800 163.700 ;
        RECT 468.400 163.600 469.200 163.700 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[0]
    PORT
      LAYER metal1 ;
        RECT 465.200 175.600 466.000 177.200 ;
        RECT 481.200 173.600 482.000 175.200 ;
        RECT 471.600 169.600 472.400 171.200 ;
        RECT 478.000 169.600 478.800 172.400 ;
        RECT 497.200 169.600 498.000 171.200 ;
      LAYER via1 ;
        RECT 478.000 171.600 478.800 172.400 ;
      LAYER metal2 ;
        RECT 465.200 175.600 466.000 176.400 ;
        RECT 465.300 172.400 465.900 175.600 ;
        RECT 481.200 173.600 482.000 174.400 ;
        RECT 481.300 172.400 481.900 173.600 ;
        RECT 465.200 171.600 466.000 172.400 ;
        RECT 471.600 171.600 472.400 172.400 ;
        RECT 478.000 171.600 478.800 172.400 ;
        RECT 481.200 171.600 482.000 172.400 ;
        RECT 497.200 171.600 498.000 172.400 ;
        RECT 471.700 170.400 472.300 171.600 ;
        RECT 497.300 170.400 497.900 171.600 ;
        RECT 471.600 169.600 472.400 170.400 ;
        RECT 497.200 169.600 498.000 170.400 ;
        RECT 497.300 168.400 497.900 169.600 ;
        RECT 497.200 167.600 498.000 168.400 ;
      LAYER metal3 ;
        RECT 465.200 172.300 466.000 172.400 ;
        RECT 471.600 172.300 472.400 172.400 ;
        RECT 478.000 172.300 478.800 172.400 ;
        RECT 481.200 172.300 482.000 172.400 ;
        RECT 497.200 172.300 498.000 172.400 ;
        RECT 465.200 171.700 498.000 172.300 ;
        RECT 465.200 171.600 466.000 171.700 ;
        RECT 471.600 171.600 472.400 171.700 ;
        RECT 478.000 171.600 478.800 171.700 ;
        RECT 481.200 171.600 482.000 171.700 ;
        RECT 497.200 171.600 498.000 171.700 ;
        RECT 537.300 169.700 555.500 170.300 ;
        RECT 497.200 168.300 498.000 168.400 ;
        RECT 537.300 168.300 537.900 169.700 ;
        RECT 497.200 167.700 537.900 168.300 ;
        RECT 497.200 167.600 498.000 167.700 ;
    END
  END wb_adr_i[0]
  PIN wb_clk_i
    PORT
      LAYER metal1 ;
        RECT 254.000 333.800 254.800 334.400 ;
        RECT 254.000 333.000 255.800 333.800 ;
        RECT 78.000 308.200 79.800 309.000 ;
        RECT 145.200 308.200 147.000 309.000 ;
        RECT 491.400 308.200 493.200 309.000 ;
        RECT 78.000 307.600 78.800 308.200 ;
        RECT 145.200 307.600 146.000 308.200 ;
        RECT 492.400 307.600 493.200 308.200 ;
        RECT 322.800 293.800 323.600 294.400 ;
        RECT 321.800 293.000 323.600 293.800 ;
        RECT 514.800 253.800 515.600 254.400 ;
        RECT 514.800 253.000 516.600 253.800 ;
        RECT 336.200 108.200 338.000 109.000 ;
        RECT 337.200 107.600 338.000 108.200 ;
        RECT 75.400 68.200 77.200 69.000 ;
        RECT 76.400 67.600 77.200 68.200 ;
        RECT 76.400 53.800 77.200 54.400 ;
        RECT 76.400 53.000 78.200 53.800 ;
        RECT 76.400 28.200 78.200 29.000 ;
        RECT 369.800 28.200 371.600 29.000 ;
        RECT 76.400 27.600 77.200 28.200 ;
        RECT 370.800 27.600 371.600 28.200 ;
        RECT 535.600 28.200 537.400 29.000 ;
        RECT 535.600 27.600 536.400 28.200 ;
      LAYER via1 ;
        RECT 254.000 333.600 254.800 334.400 ;
        RECT 322.800 293.600 323.600 294.400 ;
        RECT 514.800 253.600 515.600 254.400 ;
        RECT 76.400 53.600 77.200 54.400 ;
      LAYER metal2 ;
        RECT 254.000 333.600 254.800 334.400 ;
        RECT 254.100 310.400 254.700 333.600 ;
        RECT 254.000 309.600 254.800 310.400 ;
        RECT 322.800 309.600 323.600 310.400 ;
        RECT 78.000 307.600 78.800 308.400 ;
        RECT 145.200 307.600 146.000 308.400 ;
        RECT 322.900 302.400 323.500 309.600 ;
        RECT 492.400 307.600 493.200 308.400 ;
        RECT 492.500 302.400 493.100 307.600 ;
        RECT 322.800 301.600 323.600 302.400 ;
        RECT 492.400 301.600 493.200 302.400 ;
        RECT 322.900 294.400 323.500 301.600 ;
        RECT 322.800 293.600 323.600 294.400 ;
        RECT 322.900 292.400 323.500 293.600 ;
        RECT 322.800 291.600 323.600 292.400 ;
        RECT 514.800 255.600 515.600 256.400 ;
        RECT 514.900 254.400 515.500 255.600 ;
        RECT 514.800 253.600 515.600 254.400 ;
        RECT 337.200 123.600 338.000 124.400 ;
        RECT 337.300 108.400 337.900 123.600 ;
        RECT 337.200 107.600 338.000 108.400 ;
        RECT 337.300 102.300 337.900 107.600 ;
        RECT 337.300 101.700 339.500 102.300 ;
        RECT 76.400 67.600 77.200 68.400 ;
        RECT 76.500 54.400 77.100 67.600 ;
        RECT 338.900 66.400 339.500 101.700 ;
        RECT 338.800 65.600 339.600 66.400 ;
        RECT 370.800 65.600 371.600 66.400 ;
        RECT 76.400 53.600 77.200 54.400 ;
        RECT 76.500 28.400 77.100 53.600 ;
        RECT 370.900 28.400 371.500 65.600 ;
        RECT 76.400 27.600 77.200 28.400 ;
        RECT 370.800 27.600 371.600 28.400 ;
        RECT 535.600 27.600 536.400 28.400 ;
        RECT 370.900 4.400 371.500 27.600 ;
        RECT 535.700 4.400 536.300 27.600 ;
        RECT 370.800 3.600 371.600 4.400 ;
        RECT 516.400 3.600 517.200 4.400 ;
        RECT 535.600 3.600 536.400 4.400 ;
        RECT 516.500 -2.300 517.100 3.600 ;
      LAYER metal3 ;
        RECT 254.000 310.300 254.800 310.400 ;
        RECT 322.800 310.300 323.600 310.400 ;
        RECT 254.000 309.700 323.600 310.300 ;
        RECT 254.000 309.600 254.800 309.700 ;
        RECT 322.800 309.600 323.600 309.700 ;
        RECT 78.000 308.300 78.800 308.400 ;
        RECT 145.200 308.300 146.000 308.400 ;
        RECT 254.100 308.300 254.700 309.600 ;
        RECT 78.000 307.700 254.700 308.300 ;
        RECT 78.000 307.600 78.800 307.700 ;
        RECT 145.200 307.600 146.000 307.700 ;
        RECT 322.800 302.300 323.600 302.400 ;
        RECT 492.400 302.300 493.200 302.400 ;
        RECT 494.000 302.300 494.800 302.400 ;
        RECT 322.800 301.700 494.800 302.300 ;
        RECT 322.800 301.600 323.600 301.700 ;
        RECT 492.400 301.600 493.200 301.700 ;
        RECT 494.000 301.600 494.800 301.700 ;
        RECT 321.200 292.300 322.000 292.400 ;
        RECT 322.800 292.300 323.600 292.400 ;
        RECT 321.200 291.700 323.600 292.300 ;
        RECT 321.200 291.600 322.000 291.700 ;
        RECT 322.800 291.600 323.600 291.700 ;
        RECT 494.000 256.300 494.800 256.400 ;
        RECT 514.800 256.300 515.600 256.400 ;
        RECT 494.000 255.700 515.600 256.300 ;
        RECT 494.000 255.600 494.800 255.700 ;
        RECT 514.800 255.600 515.600 255.700 ;
        RECT 318.000 246.300 318.800 246.400 ;
        RECT 321.200 246.300 322.000 246.400 ;
        RECT 318.000 245.700 322.000 246.300 ;
        RECT 318.000 245.600 318.800 245.700 ;
        RECT 321.200 245.600 322.000 245.700 ;
        RECT 318.000 124.300 318.800 124.400 ;
        RECT 337.200 124.300 338.000 124.400 ;
        RECT 318.000 123.700 338.000 124.300 ;
        RECT 318.000 123.600 318.800 123.700 ;
        RECT 337.200 123.600 338.000 123.700 ;
        RECT 76.400 68.300 77.200 68.400 ;
        RECT 78.000 68.300 78.800 68.400 ;
        RECT 76.400 67.700 78.800 68.300 ;
        RECT 76.400 67.600 77.200 67.700 ;
        RECT 78.000 67.600 78.800 67.700 ;
        RECT 338.800 66.300 339.600 66.400 ;
        RECT 370.800 66.300 371.600 66.400 ;
        RECT 338.800 65.700 371.600 66.300 ;
        RECT 338.800 65.600 339.600 65.700 ;
        RECT 370.800 65.600 371.600 65.700 ;
        RECT 370.800 4.300 371.600 4.400 ;
        RECT 516.400 4.300 517.200 4.400 ;
        RECT 535.600 4.300 536.400 4.400 ;
        RECT 370.800 3.700 536.400 4.300 ;
        RECT 370.800 3.600 371.600 3.700 ;
        RECT 516.400 3.600 517.200 3.700 ;
        RECT 535.600 3.600 536.400 3.700 ;
      LAYER metal4 ;
        RECT 77.800 67.400 79.000 308.600 ;
        RECT 317.800 123.400 319.000 246.600 ;
        RECT 321.000 245.400 322.200 292.600 ;
        RECT 493.800 255.400 495.000 302.600 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    PORT
      LAYER metal1 ;
        RECT 542.000 311.600 542.800 313.200 ;
      LAYER metal2 ;
        RECT 542.000 311.600 542.800 312.400 ;
      LAYER metal3 ;
        RECT 542.000 312.300 542.800 312.400 ;
        RECT 542.000 311.700 555.500 312.300 ;
        RECT 542.000 311.600 542.800 311.700 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[7]
    PORT
      LAYER metal1 ;
        RECT 369.200 228.800 370.000 230.400 ;
        RECT 494.000 226.800 494.800 228.400 ;
        RECT 338.800 211.600 339.600 213.200 ;
      LAYER via1 ;
        RECT 369.200 229.600 370.000 230.400 ;
        RECT 494.000 227.600 494.800 228.400 ;
      LAYER metal2 ;
        RECT 494.000 233.600 494.800 234.400 ;
        RECT 369.200 229.600 370.000 230.400 ;
        RECT 369.300 220.400 369.900 229.600 ;
        RECT 494.100 228.400 494.700 233.600 ;
        RECT 494.000 227.600 494.800 228.400 ;
        RECT 494.100 220.400 494.700 227.600 ;
        RECT 338.800 219.600 339.600 220.400 ;
        RECT 369.200 219.600 370.000 220.400 ;
        RECT 494.000 219.600 494.800 220.400 ;
        RECT 338.900 212.400 339.500 219.600 ;
        RECT 338.800 211.600 339.600 212.400 ;
      LAYER metal3 ;
        RECT 494.000 234.300 494.800 234.400 ;
        RECT 554.900 234.300 555.500 236.300 ;
        RECT 494.000 233.700 555.500 234.300 ;
        RECT 494.000 233.600 494.800 233.700 ;
        RECT 338.800 220.300 339.600 220.400 ;
        RECT 369.200 220.300 370.000 220.400 ;
        RECT 494.000 220.300 494.800 220.400 ;
        RECT 338.800 219.700 494.800 220.300 ;
        RECT 338.800 219.600 339.600 219.700 ;
        RECT 369.200 219.600 370.000 219.700 ;
        RECT 494.000 219.600 494.800 219.700 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_i[6]
    PORT
      LAYER metal1 ;
        RECT 343.600 291.600 344.400 293.200 ;
        RECT 342.000 228.800 342.800 230.400 ;
        RECT 372.400 226.800 373.200 228.400 ;
      LAYER via1 ;
        RECT 342.000 229.600 342.800 230.400 ;
        RECT 372.400 227.600 373.200 228.400 ;
      LAYER metal2 ;
        RECT 343.700 380.400 344.300 386.300 ;
        RECT 343.600 379.600 344.400 380.400 ;
        RECT 350.000 379.600 350.800 380.400 ;
        RECT 343.600 291.600 344.400 292.400 ;
        RECT 343.700 286.400 344.300 291.600 ;
        RECT 350.100 286.400 350.700 379.600 ;
        RECT 343.600 285.600 344.400 286.400 ;
        RECT 350.000 285.600 350.800 286.400 ;
        RECT 342.000 229.600 342.800 230.400 ;
        RECT 342.100 226.400 342.700 229.600 ;
        RECT 350.100 226.400 350.700 285.600 ;
        RECT 372.400 227.600 373.200 228.400 ;
        RECT 372.500 226.400 373.100 227.600 ;
        RECT 342.000 225.600 342.800 226.400 ;
        RECT 350.000 225.600 350.800 226.400 ;
        RECT 372.400 225.600 373.200 226.400 ;
      LAYER metal3 ;
        RECT 343.600 380.300 344.400 380.400 ;
        RECT 350.000 380.300 350.800 380.400 ;
        RECT 343.600 379.700 350.800 380.300 ;
        RECT 343.600 379.600 344.400 379.700 ;
        RECT 350.000 379.600 350.800 379.700 ;
        RECT 343.600 286.300 344.400 286.400 ;
        RECT 350.000 286.300 350.800 286.400 ;
        RECT 343.600 285.700 350.800 286.300 ;
        RECT 343.600 285.600 344.400 285.700 ;
        RECT 350.000 285.600 350.800 285.700 ;
        RECT 342.000 226.300 342.800 226.400 ;
        RECT 350.000 226.300 350.800 226.400 ;
        RECT 372.400 226.300 373.200 226.400 ;
        RECT 342.000 225.700 373.200 226.300 ;
        RECT 342.000 225.600 342.800 225.700 ;
        RECT 350.000 225.600 350.800 225.700 ;
        RECT 372.400 225.600 373.200 225.700 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[5]
    PORT
      LAYER metal1 ;
        RECT 332.400 252.300 333.200 253.200 ;
        RECT 335.600 252.300 336.400 252.400 ;
        RECT 332.400 251.700 336.400 252.300 ;
        RECT 332.400 251.600 333.200 251.700 ;
        RECT 335.600 251.600 336.400 251.700 ;
        RECT 335.600 228.800 336.400 230.400 ;
        RECT 486.000 226.800 486.800 228.400 ;
      LAYER via1 ;
        RECT 335.600 229.600 336.400 230.400 ;
        RECT 486.000 227.600 486.800 228.400 ;
      LAYER metal2 ;
        RECT 335.600 251.600 336.400 252.400 ;
        RECT 335.700 234.400 336.300 251.600 ;
        RECT 486.000 235.600 486.800 236.400 ;
        RECT 335.600 233.600 336.400 234.400 ;
        RECT 335.700 230.400 336.300 233.600 ;
        RECT 335.600 229.600 336.400 230.400 ;
        RECT 486.100 228.400 486.700 235.600 ;
        RECT 486.000 227.600 486.800 228.400 ;
      LAYER metal3 ;
        RECT 486.000 236.300 486.800 236.400 ;
        RECT 551.600 236.300 552.400 236.400 ;
        RECT 430.100 235.700 552.400 236.300 ;
        RECT 335.600 234.300 336.400 234.400 ;
        RECT 430.100 234.300 430.700 235.700 ;
        RECT 486.000 235.600 486.800 235.700 ;
        RECT 551.600 235.600 552.400 235.700 ;
        RECT 335.600 233.700 430.700 234.300 ;
        RECT 335.600 233.600 336.400 233.700 ;
        RECT 551.600 228.300 552.400 228.400 ;
        RECT 551.600 227.700 555.500 228.300 ;
        RECT 551.600 227.600 552.400 227.700 ;
      LAYER metal4 ;
        RECT 551.400 227.400 552.600 236.600 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[4]
    PORT
      LAYER metal1 ;
        RECT 348.400 148.800 349.200 150.400 ;
        RECT 364.400 146.800 365.200 148.400 ;
        RECT 319.600 131.600 320.400 133.200 ;
      LAYER via1 ;
        RECT 348.400 149.600 349.200 150.400 ;
        RECT 364.400 147.600 365.200 148.400 ;
      LAYER metal2 ;
        RECT 348.400 149.600 349.200 150.400 ;
        RECT 348.500 148.400 349.100 149.600 ;
        RECT 348.400 147.600 349.200 148.400 ;
        RECT 364.400 147.600 365.200 148.400 ;
        RECT 348.500 136.400 349.100 147.600 ;
        RECT 319.600 135.600 320.400 136.400 ;
        RECT 348.400 135.600 349.200 136.400 ;
        RECT 319.700 132.400 320.300 135.600 ;
        RECT 319.600 131.600 320.400 132.400 ;
        RECT 319.700 100.400 320.300 131.600 ;
        RECT 319.600 99.600 320.400 100.400 ;
        RECT 326.000 1.600 326.800 2.400 ;
        RECT 326.100 -2.300 326.700 1.600 ;
      LAYER metal3 ;
        RECT 348.400 148.300 349.200 148.400 ;
        RECT 364.400 148.300 365.200 148.400 ;
        RECT 348.400 147.700 365.200 148.300 ;
        RECT 348.400 147.600 349.200 147.700 ;
        RECT 364.400 147.600 365.200 147.700 ;
        RECT 319.600 136.300 320.400 136.400 ;
        RECT 348.400 136.300 349.200 136.400 ;
        RECT 319.600 135.700 349.200 136.300 ;
        RECT 319.600 135.600 320.400 135.700 ;
        RECT 348.400 135.600 349.200 135.700 ;
        RECT 319.600 100.300 320.400 100.400 ;
        RECT 321.200 100.300 322.000 100.400 ;
        RECT 319.600 99.700 322.000 100.300 ;
        RECT 319.600 99.600 320.400 99.700 ;
        RECT 321.200 99.600 322.000 99.700 ;
        RECT 321.200 2.300 322.000 2.400 ;
        RECT 326.000 2.300 326.800 2.400 ;
        RECT 321.200 1.700 326.800 2.300 ;
        RECT 321.200 1.600 322.000 1.700 ;
        RECT 326.000 1.600 326.800 1.700 ;
      LAYER metal4 ;
        RECT 321.000 1.400 322.200 100.600 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[3]
    PORT
      LAYER metal1 ;
        RECT 406.000 184.800 406.800 186.400 ;
        RECT 346.800 172.300 347.600 173.200 ;
        RECT 348.400 172.300 349.200 172.400 ;
        RECT 346.800 171.700 349.200 172.300 ;
        RECT 346.800 171.600 347.600 171.700 ;
        RECT 348.400 171.600 349.200 171.700 ;
        RECT 342.000 148.800 342.800 150.400 ;
        RECT 466.800 108.300 467.600 108.400 ;
        RECT 468.400 108.300 469.200 108.400 ;
        RECT 466.800 107.700 469.200 108.300 ;
        RECT 466.800 107.600 467.600 107.700 ;
        RECT 468.400 106.800 469.200 107.700 ;
      LAYER via1 ;
        RECT 406.000 185.600 406.800 186.400 ;
        RECT 342.000 149.600 342.800 150.400 ;
      LAYER metal2 ;
        RECT 406.000 185.600 406.800 186.400 ;
        RECT 348.400 171.600 349.200 172.400 ;
        RECT 348.500 170.400 349.100 171.600 ;
        RECT 342.000 169.600 342.800 170.400 ;
        RECT 348.400 169.600 349.200 170.400 ;
        RECT 342.100 150.400 342.700 169.600 ;
        RECT 342.000 149.600 342.800 150.400 ;
        RECT 466.800 107.600 467.600 108.400 ;
        RECT 466.900 100.400 467.500 107.600 ;
        RECT 466.800 99.600 467.600 100.400 ;
        RECT 470.000 1.600 470.800 2.400 ;
        RECT 470.100 -2.300 470.700 1.600 ;
      LAYER metal3 ;
        RECT 406.000 186.300 406.800 186.400 ;
        RECT 407.600 186.300 408.400 186.400 ;
        RECT 406.000 185.700 408.400 186.300 ;
        RECT 406.000 185.600 406.800 185.700 ;
        RECT 407.600 185.600 408.400 185.700 ;
        RECT 342.000 170.300 342.800 170.400 ;
        RECT 348.400 170.300 349.200 170.400 ;
        RECT 407.600 170.300 408.400 170.400 ;
        RECT 342.000 169.700 408.400 170.300 ;
        RECT 342.000 169.600 342.800 169.700 ;
        RECT 348.400 169.600 349.200 169.700 ;
        RECT 407.600 169.600 408.400 169.700 ;
        RECT 407.600 106.300 408.400 106.400 ;
        RECT 452.400 106.300 453.200 106.400 ;
        RECT 407.600 105.700 453.200 106.300 ;
        RECT 407.600 105.600 408.400 105.700 ;
        RECT 452.400 105.600 453.200 105.700 ;
        RECT 452.400 100.300 453.200 100.400 ;
        RECT 466.800 100.300 467.600 100.400 ;
        RECT 452.400 99.700 467.600 100.300 ;
        RECT 452.400 99.600 453.200 99.700 ;
        RECT 466.800 99.600 467.600 99.700 ;
        RECT 452.400 2.300 453.200 2.400 ;
        RECT 470.000 2.300 470.800 2.400 ;
        RECT 452.400 1.700 470.800 2.300 ;
        RECT 452.400 1.600 453.200 1.700 ;
        RECT 470.000 1.600 470.800 1.700 ;
      LAYER metal4 ;
        RECT 407.400 105.400 408.600 186.600 ;
        RECT 452.200 1.400 453.400 106.600 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[2]
    PORT
      LAYER metal1 ;
        RECT 310.000 108.800 310.800 110.400 ;
        RECT 260.400 68.800 261.200 70.400 ;
        RECT 316.400 55.600 317.200 57.200 ;
      LAYER via1 ;
        RECT 310.000 109.600 310.800 110.400 ;
        RECT 260.400 69.600 261.200 70.400 ;
      LAYER metal2 ;
        RECT 310.000 109.600 310.800 110.400 ;
        RECT 310.100 82.400 310.700 109.600 ;
        RECT 260.400 81.600 261.200 82.400 ;
        RECT 310.000 81.600 310.800 82.400 ;
        RECT 316.400 81.600 317.200 82.400 ;
        RECT 260.500 70.400 261.100 81.600 ;
        RECT 260.400 69.600 261.200 70.400 ;
        RECT 316.500 56.400 317.100 81.600 ;
        RECT 316.400 55.600 317.200 56.400 ;
        RECT 316.500 -2.300 317.100 55.600 ;
      LAYER metal3 ;
        RECT 260.400 82.300 261.200 82.400 ;
        RECT 310.000 82.300 310.800 82.400 ;
        RECT 316.400 82.300 317.200 82.400 ;
        RECT 260.400 81.700 317.200 82.300 ;
        RECT 260.400 81.600 261.200 81.700 ;
        RECT 310.000 81.600 310.800 81.700 ;
        RECT 316.400 81.600 317.200 81.700 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[1]
    PORT
      LAYER metal1 ;
        RECT 354.800 150.300 355.600 150.400 ;
        RECT 358.000 150.300 358.800 150.400 ;
        RECT 354.800 149.700 358.800 150.300 ;
        RECT 354.800 148.800 355.600 149.700 ;
        RECT 358.000 149.600 358.800 149.700 ;
        RECT 358.000 135.600 358.800 137.200 ;
        RECT 351.600 91.600 352.400 93.200 ;
      LAYER metal2 ;
        RECT 358.000 149.600 358.800 150.400 ;
        RECT 358.100 136.400 358.700 149.600 ;
        RECT 358.000 135.600 358.800 136.400 ;
        RECT 358.100 120.400 358.700 135.600 ;
        RECT 358.000 119.600 358.800 120.400 ;
        RECT 351.600 91.600 352.400 92.400 ;
        RECT 351.600 1.600 352.400 2.400 ;
        RECT 351.700 -2.300 352.300 1.600 ;
      LAYER metal3 ;
        RECT 353.200 120.300 354.000 120.400 ;
        RECT 358.000 120.300 358.800 120.400 ;
        RECT 353.200 119.700 358.800 120.300 ;
        RECT 353.200 119.600 354.000 119.700 ;
        RECT 358.000 119.600 358.800 119.700 ;
        RECT 350.000 92.300 350.800 92.400 ;
        RECT 351.600 92.300 352.400 92.400 ;
        RECT 353.200 92.300 354.000 92.400 ;
        RECT 350.000 91.700 354.000 92.300 ;
        RECT 350.000 91.600 350.800 91.700 ;
        RECT 351.600 91.600 352.400 91.700 ;
        RECT 353.200 91.600 354.000 91.700 ;
        RECT 350.000 2.300 350.800 2.400 ;
        RECT 351.600 2.300 352.400 2.400 ;
        RECT 350.000 1.700 352.400 2.300 ;
        RECT 350.000 1.600 350.800 1.700 ;
        RECT 351.600 1.600 352.400 1.700 ;
      LAYER metal4 ;
        RECT 349.800 1.400 351.000 92.600 ;
        RECT 353.000 91.400 354.200 120.600 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[0]
    PORT
      LAYER metal1 ;
        RECT 359.600 148.800 360.400 150.400 ;
        RECT 398.000 104.800 398.800 106.400 ;
        RECT 318.000 68.800 318.800 70.400 ;
      LAYER via1 ;
        RECT 359.600 149.600 360.400 150.400 ;
        RECT 398.000 105.600 398.800 106.400 ;
        RECT 318.000 69.600 318.800 70.400 ;
      LAYER metal2 ;
        RECT 359.600 149.600 360.400 150.400 ;
        RECT 359.700 130.400 360.300 149.600 ;
        RECT 335.600 129.600 336.400 130.400 ;
        RECT 359.600 129.600 360.400 130.400 ;
        RECT 398.000 129.600 398.800 130.400 ;
        RECT 335.700 70.400 336.300 129.600 ;
        RECT 398.100 106.400 398.700 129.600 ;
        RECT 398.000 105.600 398.800 106.400 ;
        RECT 318.000 69.600 318.800 70.400 ;
        RECT 322.800 69.600 323.600 70.400 ;
        RECT 335.600 69.600 336.400 70.400 ;
        RECT 322.900 -1.700 323.500 69.600 ;
        RECT 321.300 -2.300 323.500 -1.700 ;
      LAYER metal3 ;
        RECT 335.600 130.300 336.400 130.400 ;
        RECT 359.600 130.300 360.400 130.400 ;
        RECT 398.000 130.300 398.800 130.400 ;
        RECT 335.600 129.700 398.800 130.300 ;
        RECT 335.600 129.600 336.400 129.700 ;
        RECT 359.600 129.600 360.400 129.700 ;
        RECT 398.000 129.600 398.800 129.700 ;
        RECT 318.000 70.300 318.800 70.400 ;
        RECT 322.800 70.300 323.600 70.400 ;
        RECT 335.600 70.300 336.400 70.400 ;
        RECT 318.000 69.700 336.400 70.300 ;
        RECT 318.000 69.600 318.800 69.700 ;
        RECT 322.800 69.600 323.600 69.700 ;
        RECT 335.600 69.600 336.400 69.700 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_o[7]
    PORT
      LAYER metal1 ;
        RECT 342.000 311.800 342.800 319.800 ;
        RECT 342.000 309.600 342.600 311.800 ;
        RECT 342.000 302.200 342.800 309.600 ;
      LAYER via1 ;
        RECT 342.000 317.600 342.800 318.400 ;
      LAYER metal2 ;
        RECT 340.500 382.400 341.100 386.300 ;
        RECT 340.400 381.600 341.200 382.400 ;
        RECT 348.400 381.600 349.200 382.400 ;
        RECT 348.500 338.400 349.100 381.600 ;
        RECT 342.000 337.600 342.800 338.400 ;
        RECT 348.400 337.600 349.200 338.400 ;
        RECT 342.100 318.400 342.700 337.600 ;
        RECT 342.000 317.600 342.800 318.400 ;
      LAYER metal3 ;
        RECT 340.400 382.300 341.200 382.400 ;
        RECT 348.400 382.300 349.200 382.400 ;
        RECT 340.400 381.700 349.200 382.300 ;
        RECT 340.400 381.600 341.200 381.700 ;
        RECT 348.400 381.600 349.200 381.700 ;
        RECT 342.000 338.300 342.800 338.400 ;
        RECT 348.400 338.300 349.200 338.400 ;
        RECT 342.000 337.700 349.200 338.300 ;
        RECT 342.000 337.600 342.800 337.700 ;
        RECT 348.400 337.600 349.200 337.700 ;
    END
  END wb_dat_o[7]
  PIN wb_dat_o[6]
    PORT
      LAYER metal1 ;
        RECT 548.400 12.400 549.200 19.800 ;
        RECT 548.600 10.200 549.200 12.400 ;
        RECT 548.400 8.300 549.200 10.200 ;
        RECT 551.600 8.300 552.400 8.400 ;
        RECT 548.400 7.700 552.400 8.300 ;
        RECT 548.400 2.200 549.200 7.700 ;
        RECT 551.600 7.600 552.400 7.700 ;
      LAYER metal2 ;
        RECT 551.600 9.600 552.400 10.400 ;
        RECT 551.700 8.400 552.300 9.600 ;
        RECT 551.600 7.600 552.400 8.400 ;
      LAYER metal3 ;
        RECT 551.600 10.300 552.400 10.400 ;
        RECT 551.600 9.700 555.500 10.300 ;
        RECT 551.600 9.600 552.400 9.700 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[5]
    PORT
      LAYER metal1 ;
        RECT 548.400 271.800 549.200 279.800 ;
        RECT 548.600 269.600 549.200 271.800 ;
        RECT 548.400 268.300 549.200 269.600 ;
        RECT 551.600 268.300 552.400 268.400 ;
        RECT 548.400 267.700 552.400 268.300 ;
        RECT 548.400 262.200 549.200 267.700 ;
        RECT 551.600 267.600 552.400 267.700 ;
      LAYER metal2 ;
        RECT 551.600 269.600 552.400 270.400 ;
        RECT 551.700 268.400 552.300 269.600 ;
        RECT 551.600 267.600 552.400 268.400 ;
      LAYER metal3 ;
        RECT 551.600 270.300 552.400 270.400 ;
        RECT 551.600 269.700 555.500 270.300 ;
        RECT 551.600 269.600 552.400 269.700 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[4]
    PORT
      LAYER metal1 ;
        RECT 545.200 332.400 546.000 339.800 ;
        RECT 545.200 330.200 545.800 332.400 ;
        RECT 545.200 322.200 546.000 330.200 ;
      LAYER via1 ;
        RECT 545.200 327.600 546.000 328.400 ;
      LAYER metal2 ;
        RECT 545.200 329.600 546.000 330.400 ;
        RECT 545.300 328.400 545.900 329.600 ;
        RECT 545.200 327.600 546.000 328.400 ;
      LAYER metal3 ;
        RECT 545.200 330.300 546.000 330.400 ;
        RECT 545.200 329.700 555.500 330.300 ;
        RECT 545.200 329.600 546.000 329.700 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[3]
    PORT
      LAYER metal1 ;
        RECT 460.400 12.400 461.200 19.800 ;
        RECT 460.600 10.200 461.200 12.400 ;
        RECT 460.400 2.200 461.200 10.200 ;
      LAYER via1 ;
        RECT 460.400 3.600 461.200 4.400 ;
      LAYER metal2 ;
        RECT 460.400 3.600 461.200 4.400 ;
        RECT 460.500 -1.700 461.100 3.600 ;
        RECT 458.900 -2.300 461.100 -1.700 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[2]
    PORT
      LAYER metal1 ;
        RECT 548.400 151.800 549.200 159.800 ;
        RECT 548.600 149.600 549.200 151.800 ;
        RECT 548.400 148.300 549.200 149.600 ;
        RECT 551.600 148.300 552.400 148.400 ;
        RECT 548.400 147.700 552.400 148.300 ;
        RECT 548.400 142.200 549.200 147.700 ;
        RECT 551.600 147.600 552.400 147.700 ;
      LAYER metal2 ;
        RECT 551.600 149.600 552.400 150.400 ;
        RECT 551.700 148.400 552.300 149.600 ;
        RECT 551.600 147.600 552.400 148.400 ;
      LAYER metal3 ;
        RECT 551.600 150.300 552.400 150.400 ;
        RECT 551.600 149.700 555.500 150.300 ;
        RECT 551.600 149.600 552.400 149.700 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[1]
    PORT
      LAYER metal1 ;
        RECT 465.200 12.400 466.000 19.800 ;
        RECT 465.400 10.200 466.000 12.400 ;
        RECT 465.200 2.200 466.000 10.200 ;
      LAYER via1 ;
        RECT 465.200 3.600 466.000 4.400 ;
      LAYER metal2 ;
        RECT 465.200 3.600 466.000 4.400 ;
        RECT 465.300 -1.700 465.900 3.600 ;
        RECT 463.700 -2.300 465.900 -1.700 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[0]
    PORT
      LAYER metal1 ;
        RECT 372.400 12.400 373.200 19.800 ;
        RECT 372.400 10.200 373.000 12.400 ;
        RECT 372.400 2.200 373.200 10.200 ;
      LAYER via1 ;
        RECT 372.400 3.600 373.200 4.400 ;
      LAYER metal2 ;
        RECT 372.400 3.600 373.200 4.400 ;
        RECT 372.500 -1.700 373.100 3.600 ;
        RECT 372.500 -2.300 374.700 -1.700 ;
    END
  END wb_dat_o[0]
  PIN wb_inta_o
    PORT
      LAYER metal1 ;
        RECT 543.600 12.400 544.400 19.800 ;
        RECT 543.800 10.200 544.400 12.400 ;
        RECT 543.600 2.200 544.400 10.200 ;
      LAYER via1 ;
        RECT 543.600 3.600 544.400 4.400 ;
      LAYER metal2 ;
        RECT 543.600 3.600 544.400 4.400 ;
        RECT 543.700 -1.700 544.300 3.600 ;
        RECT 542.100 -2.300 544.300 -1.700 ;
    END
  END wb_inta_o
  PIN wb_rst_i
    PORT
      LAYER metal1 ;
        RECT 348.400 230.300 349.200 230.400 ;
        RECT 350.000 230.300 350.800 230.400 ;
        RECT 348.400 229.700 350.800 230.300 ;
        RECT 348.400 228.800 349.200 229.700 ;
        RECT 350.000 228.800 350.800 229.700 ;
        RECT 350.000 171.600 350.800 173.200 ;
        RECT 246.000 68.800 246.800 70.400 ;
        RECT 321.200 68.800 322.000 70.400 ;
        RECT 270.000 51.600 270.800 53.200 ;
      LAYER via1 ;
        RECT 348.400 229.600 349.200 230.400 ;
        RECT 246.000 69.600 246.800 70.400 ;
        RECT 321.200 69.600 322.000 70.400 ;
      LAYER metal2 ;
        RECT 348.400 229.600 349.200 230.400 ;
        RECT 348.500 204.300 349.100 229.600 ;
        RECT 348.500 203.700 350.700 204.300 ;
        RECT 350.100 172.400 350.700 203.700 ;
        RECT 350.000 171.600 350.800 172.400 ;
        RECT 350.100 168.400 350.700 171.600 ;
        RECT 350.000 167.600 350.800 168.400 ;
        RECT 321.200 77.600 322.000 78.400 ;
        RECT 321.300 70.400 321.900 77.600 ;
        RECT 246.000 69.600 246.800 70.400 ;
        RECT 321.200 69.600 322.000 70.400 ;
        RECT 246.100 68.400 246.700 69.600 ;
        RECT 321.300 68.400 321.900 69.600 ;
        RECT 246.000 67.600 246.800 68.400 ;
        RECT 270.000 67.600 270.800 68.400 ;
        RECT 282.800 67.600 283.600 68.400 ;
        RECT 321.200 67.600 322.000 68.400 ;
        RECT 270.100 52.400 270.700 67.600 ;
        RECT 270.000 51.600 270.800 52.400 ;
        RECT 282.900 -1.700 283.500 67.600 ;
        RECT 281.300 -2.300 283.500 -1.700 ;
      LAYER metal3 ;
        RECT 327.600 168.300 328.400 168.400 ;
        RECT 350.000 168.300 350.800 168.400 ;
        RECT 327.600 167.700 350.800 168.300 ;
        RECT 327.600 167.600 328.400 167.700 ;
        RECT 350.000 167.600 350.800 167.700 ;
        RECT 321.200 78.300 322.000 78.400 ;
        RECT 327.600 78.300 328.400 78.400 ;
        RECT 321.200 77.700 328.400 78.300 ;
        RECT 321.200 77.600 322.000 77.700 ;
        RECT 327.600 77.600 328.400 77.700 ;
        RECT 246.000 68.300 246.800 68.400 ;
        RECT 270.000 68.300 270.800 68.400 ;
        RECT 282.800 68.300 283.600 68.400 ;
        RECT 321.200 68.300 322.000 68.400 ;
        RECT 246.000 67.700 322.000 68.300 ;
        RECT 246.000 67.600 246.800 67.700 ;
        RECT 270.000 67.600 270.800 67.700 ;
        RECT 282.800 67.600 283.600 67.700 ;
        RECT 321.200 67.600 322.000 67.700 ;
      LAYER metal4 ;
        RECT 327.400 77.400 328.600 168.600 ;
    END
  END wb_rst_i
  PIN wb_stb_i
    PORT
      LAYER metal1 ;
        RECT 545.200 308.300 546.000 308.400 ;
        RECT 551.600 308.300 552.400 308.400 ;
        RECT 545.200 307.700 552.400 308.300 ;
        RECT 545.200 306.800 546.000 307.700 ;
        RECT 551.600 307.600 552.400 307.700 ;
      LAYER metal2 ;
        RECT 551.600 307.600 552.400 308.400 ;
      LAYER metal3 ;
        RECT 551.600 308.300 552.400 308.400 ;
        RECT 551.600 307.700 555.500 308.300 ;
        RECT 551.600 307.600 552.400 307.700 ;
    END
  END wb_stb_i
  PIN wb_we_i
    PORT
      LAYER metal1 ;
        RECT 534.800 230.400 535.600 230.800 ;
        RECT 534.800 229.800 536.400 230.400 ;
        RECT 535.600 229.600 536.400 229.800 ;
        RECT 540.400 226.800 541.200 228.400 ;
      LAYER via1 ;
        RECT 540.400 227.600 541.200 228.400 ;
      LAYER metal2 ;
        RECT 535.600 231.600 536.400 232.400 ;
        RECT 540.400 231.600 541.200 232.400 ;
        RECT 535.700 230.400 536.300 231.600 ;
        RECT 535.600 229.600 536.400 230.400 ;
        RECT 540.500 228.400 541.100 231.600 ;
        RECT 540.400 227.600 541.200 228.400 ;
      LAYER metal3 ;
        RECT 535.600 232.300 536.400 232.400 ;
        RECT 540.400 232.300 541.200 232.400 ;
        RECT 535.600 231.700 555.500 232.300 ;
        RECT 535.600 231.600 536.400 231.700 ;
        RECT 540.400 231.600 541.200 231.700 ;
    END
  END wb_we_i
  OBS
      LAYER metal1 ;
        RECT 2.800 376.000 3.600 379.800 ;
        RECT 2.600 375.200 3.600 376.000 ;
        RECT 2.600 370.800 3.400 375.200 ;
        RECT 4.400 374.600 5.200 379.800 ;
        RECT 10.800 376.600 11.600 379.800 ;
        RECT 12.400 377.000 13.200 379.800 ;
        RECT 14.000 377.000 14.800 379.800 ;
        RECT 15.600 377.000 16.400 379.800 ;
        RECT 17.200 377.000 18.000 379.800 ;
        RECT 20.400 377.000 21.200 379.800 ;
        RECT 23.600 377.000 24.400 379.800 ;
        RECT 25.200 377.000 26.000 379.800 ;
        RECT 26.800 377.000 27.600 379.800 ;
        RECT 9.200 375.800 11.600 376.600 ;
        RECT 28.400 376.600 29.200 379.800 ;
        RECT 9.200 375.200 10.000 375.800 ;
        RECT 4.000 374.000 5.200 374.600 ;
        RECT 8.200 374.600 10.000 375.200 ;
        RECT 14.000 375.600 15.000 376.400 ;
        RECT 18.000 375.600 19.600 376.400 ;
        RECT 20.400 375.800 25.000 376.400 ;
        RECT 28.400 375.800 31.000 376.600 ;
        RECT 20.400 375.600 21.200 375.800 ;
        RECT 4.000 372.000 4.600 374.000 ;
        RECT 8.200 373.400 9.000 374.600 ;
        RECT 5.200 372.600 9.000 373.400 ;
        RECT 14.000 372.800 14.800 375.600 ;
        RECT 20.400 374.800 21.200 375.000 ;
        RECT 16.800 374.200 21.200 374.800 ;
        RECT 16.800 374.000 17.600 374.200 ;
        RECT 22.000 373.600 22.800 375.200 ;
        RECT 24.200 373.400 25.000 375.800 ;
        RECT 30.200 375.200 31.000 375.800 ;
        RECT 30.200 374.400 33.200 375.200 ;
        RECT 34.800 373.800 35.600 379.800 ;
        RECT 17.200 372.600 20.400 373.400 ;
        RECT 24.200 372.600 26.200 373.400 ;
        RECT 26.800 373.000 35.600 373.800 ;
        RECT 10.800 372.000 11.600 372.600 ;
        RECT 28.400 372.000 29.200 372.400 ;
        RECT 31.600 372.000 32.400 372.400 ;
        RECT 33.400 372.000 34.200 372.200 ;
        RECT 4.000 371.400 4.800 372.000 ;
        RECT 10.800 371.400 34.200 372.000 ;
        RECT 2.600 370.000 3.600 370.800 ;
        RECT 1.200 368.300 2.000 368.400 ;
        RECT 2.800 368.300 3.600 370.000 ;
        RECT 1.200 367.700 3.600 368.300 ;
        RECT 1.200 367.600 2.000 367.700 ;
        RECT 2.800 362.200 3.600 367.700 ;
        RECT 4.200 369.600 4.800 371.400 ;
        RECT 4.200 369.000 13.200 369.600 ;
        RECT 4.200 367.400 4.800 369.000 ;
        RECT 12.400 368.800 13.200 369.000 ;
        RECT 15.600 369.000 24.200 369.600 ;
        RECT 15.600 368.800 16.400 369.000 ;
        RECT 7.400 367.600 10.000 368.400 ;
        RECT 4.200 366.800 6.800 367.400 ;
        RECT 6.000 362.200 6.800 366.800 ;
        RECT 9.200 362.200 10.000 367.600 ;
        RECT 10.600 366.800 14.800 367.600 ;
        RECT 12.400 362.200 13.200 365.000 ;
        RECT 14.000 362.200 14.800 365.000 ;
        RECT 15.600 362.200 16.400 365.000 ;
        RECT 17.200 362.200 18.000 368.400 ;
        RECT 20.400 367.600 23.000 368.400 ;
        RECT 23.600 368.200 24.200 369.000 ;
        RECT 25.200 369.400 26.000 369.600 ;
        RECT 25.200 369.000 30.600 369.400 ;
        RECT 25.200 368.800 31.400 369.000 ;
        RECT 30.000 368.200 31.400 368.800 ;
        RECT 23.600 367.600 29.400 368.200 ;
        RECT 32.400 368.000 34.000 368.800 ;
        RECT 32.400 367.600 33.000 368.000 ;
        RECT 20.400 362.200 21.200 367.000 ;
        RECT 23.600 362.200 24.400 367.000 ;
        RECT 28.800 366.800 33.000 367.600 ;
        RECT 34.800 367.400 35.600 373.000 ;
        RECT 33.600 366.800 35.600 367.400 ;
        RECT 36.400 373.800 37.200 379.800 ;
        RECT 42.800 376.600 43.600 379.800 ;
        RECT 44.400 377.000 45.200 379.800 ;
        RECT 46.000 377.000 46.800 379.800 ;
        RECT 47.600 377.000 48.400 379.800 ;
        RECT 50.800 377.000 51.600 379.800 ;
        RECT 54.000 377.000 54.800 379.800 ;
        RECT 55.600 377.000 56.400 379.800 ;
        RECT 57.200 377.000 58.000 379.800 ;
        RECT 58.800 377.000 59.600 379.800 ;
        RECT 41.000 375.800 43.600 376.600 ;
        RECT 60.400 376.600 61.200 379.800 ;
        RECT 47.000 375.800 51.600 376.400 ;
        RECT 41.000 375.200 41.800 375.800 ;
        RECT 38.800 374.400 41.800 375.200 ;
        RECT 36.400 373.000 45.200 373.800 ;
        RECT 47.000 373.400 47.800 375.800 ;
        RECT 50.800 375.600 51.600 375.800 ;
        RECT 52.400 375.600 54.000 376.400 ;
        RECT 57.000 375.600 58.000 376.400 ;
        RECT 60.400 375.800 62.800 376.600 ;
        RECT 49.200 373.600 50.000 375.200 ;
        RECT 50.800 374.800 51.600 375.000 ;
        RECT 50.800 374.200 55.200 374.800 ;
        RECT 54.400 374.000 55.200 374.200 ;
        RECT 36.400 367.400 37.200 373.000 ;
        RECT 45.800 372.600 47.800 373.400 ;
        RECT 51.600 372.600 54.800 373.400 ;
        RECT 57.200 372.800 58.000 375.600 ;
        RECT 62.000 375.200 62.800 375.800 ;
        RECT 62.000 374.600 63.800 375.200 ;
        RECT 63.000 373.400 63.800 374.600 ;
        RECT 66.800 374.600 67.600 379.800 ;
        RECT 68.400 376.000 69.200 379.800 ;
        RECT 73.200 376.000 74.000 379.800 ;
        RECT 68.400 375.200 69.400 376.000 ;
        RECT 66.800 374.000 68.000 374.600 ;
        RECT 63.000 372.600 66.800 373.400 ;
        RECT 38.000 372.200 38.800 372.400 ;
        RECT 37.800 372.000 38.800 372.200 ;
        RECT 42.800 372.000 43.600 372.400 ;
        RECT 60.400 372.000 61.200 372.600 ;
        RECT 67.400 372.000 68.000 374.000 ;
        RECT 37.800 371.400 61.200 372.000 ;
        RECT 67.200 371.400 68.000 372.000 ;
        RECT 67.200 369.600 67.800 371.400 ;
        RECT 68.600 370.800 69.400 375.200 ;
        RECT 46.000 369.400 46.800 369.600 ;
        RECT 41.400 369.000 46.800 369.400 ;
        RECT 40.600 368.800 46.800 369.000 ;
        RECT 47.800 369.000 56.400 369.600 ;
        RECT 38.000 368.000 39.600 368.800 ;
        RECT 40.600 368.200 42.000 368.800 ;
        RECT 47.800 368.200 48.400 369.000 ;
        RECT 55.600 368.800 56.400 369.000 ;
        RECT 58.800 369.000 67.800 369.600 ;
        RECT 58.800 368.800 59.600 369.000 ;
        RECT 39.000 367.600 39.600 368.000 ;
        RECT 42.600 367.600 48.400 368.200 ;
        RECT 49.000 367.600 51.600 368.400 ;
        RECT 36.400 366.800 38.400 367.400 ;
        RECT 39.000 366.800 43.200 367.600 ;
        RECT 25.200 362.200 26.000 365.000 ;
        RECT 26.800 362.200 27.600 365.000 ;
        RECT 30.000 362.200 30.800 366.800 ;
        RECT 33.600 366.200 34.200 366.800 ;
        RECT 33.200 365.600 34.200 366.200 ;
        RECT 37.800 366.200 38.400 366.800 ;
        RECT 37.800 365.600 38.800 366.200 ;
        RECT 33.200 362.200 34.000 365.600 ;
        RECT 38.000 362.200 38.800 365.600 ;
        RECT 41.200 362.200 42.000 366.800 ;
        RECT 44.400 362.200 45.200 365.000 ;
        RECT 46.000 362.200 46.800 365.000 ;
        RECT 47.600 362.200 48.400 367.000 ;
        RECT 50.800 362.200 51.600 367.000 ;
        RECT 54.000 362.200 54.800 368.400 ;
        RECT 62.000 367.600 64.600 368.400 ;
        RECT 57.200 366.800 61.400 367.600 ;
        RECT 55.600 362.200 56.400 365.000 ;
        RECT 57.200 362.200 58.000 365.000 ;
        RECT 58.800 362.200 59.600 365.000 ;
        RECT 62.000 362.200 62.800 367.600 ;
        RECT 67.200 367.400 67.800 369.000 ;
        RECT 65.200 366.800 67.800 367.400 ;
        RECT 68.400 370.000 69.400 370.800 ;
        RECT 73.000 375.200 74.000 376.000 ;
        RECT 73.000 370.800 73.800 375.200 ;
        RECT 74.800 374.600 75.600 379.800 ;
        RECT 81.200 376.600 82.000 379.800 ;
        RECT 82.800 377.000 83.600 379.800 ;
        RECT 84.400 377.000 85.200 379.800 ;
        RECT 86.000 377.000 86.800 379.800 ;
        RECT 87.600 377.000 88.400 379.800 ;
        RECT 90.800 377.000 91.600 379.800 ;
        RECT 94.000 377.000 94.800 379.800 ;
        RECT 95.600 377.000 96.400 379.800 ;
        RECT 97.200 377.000 98.000 379.800 ;
        RECT 79.600 375.800 82.000 376.600 ;
        RECT 98.800 376.600 99.600 379.800 ;
        RECT 79.600 375.200 80.400 375.800 ;
        RECT 74.400 374.000 75.600 374.600 ;
        RECT 78.600 374.600 80.400 375.200 ;
        RECT 84.400 375.600 85.400 376.400 ;
        RECT 88.400 375.600 90.000 376.400 ;
        RECT 90.800 375.800 95.400 376.400 ;
        RECT 98.800 375.800 101.400 376.600 ;
        RECT 90.800 375.600 91.600 375.800 ;
        RECT 74.400 372.000 75.000 374.000 ;
        RECT 78.600 373.400 79.400 374.600 ;
        RECT 75.600 372.600 79.400 373.400 ;
        RECT 84.400 372.800 85.200 375.600 ;
        RECT 90.800 374.800 91.600 375.000 ;
        RECT 87.200 374.200 91.600 374.800 ;
        RECT 87.200 374.000 88.000 374.200 ;
        RECT 92.400 373.600 93.200 375.200 ;
        RECT 94.600 373.400 95.400 375.800 ;
        RECT 100.600 375.200 101.400 375.800 ;
        RECT 100.600 374.400 103.600 375.200 ;
        RECT 105.200 373.800 106.000 379.800 ;
        RECT 114.800 376.000 115.600 379.800 ;
        RECT 87.600 372.600 90.800 373.400 ;
        RECT 94.600 372.600 96.600 373.400 ;
        RECT 97.200 373.000 106.000 373.800 ;
        RECT 81.200 372.000 82.000 372.600 ;
        RECT 98.800 372.000 99.600 372.400 ;
        RECT 100.400 372.000 101.200 372.400 ;
        RECT 103.800 372.000 104.600 372.200 ;
        RECT 74.400 371.400 75.200 372.000 ;
        RECT 81.200 371.400 104.600 372.000 ;
        RECT 73.000 370.000 74.000 370.800 ;
        RECT 65.200 362.200 66.000 366.800 ;
        RECT 68.400 362.200 69.200 370.000 ;
        RECT 73.200 362.200 74.000 370.000 ;
        RECT 74.600 369.600 75.200 371.400 ;
        RECT 74.600 369.000 83.600 369.600 ;
        RECT 74.600 367.400 75.200 369.000 ;
        RECT 82.800 368.800 83.600 369.000 ;
        RECT 86.000 369.000 94.600 369.600 ;
        RECT 86.000 368.800 86.800 369.000 ;
        RECT 77.800 367.600 80.400 368.400 ;
        RECT 74.600 366.800 77.200 367.400 ;
        RECT 76.400 362.200 77.200 366.800 ;
        RECT 79.600 362.200 80.400 367.600 ;
        RECT 81.000 366.800 85.200 367.600 ;
        RECT 82.800 362.200 83.600 365.000 ;
        RECT 84.400 362.200 85.200 365.000 ;
        RECT 86.000 362.200 86.800 365.000 ;
        RECT 87.600 362.200 88.400 368.400 ;
        RECT 90.800 367.600 93.400 368.400 ;
        RECT 94.000 368.200 94.600 369.000 ;
        RECT 95.600 369.400 96.400 369.600 ;
        RECT 95.600 369.000 101.000 369.400 ;
        RECT 95.600 368.800 101.800 369.000 ;
        RECT 100.400 368.200 101.800 368.800 ;
        RECT 94.000 367.600 99.800 368.200 ;
        RECT 102.800 368.000 104.400 368.800 ;
        RECT 102.800 367.600 103.400 368.000 ;
        RECT 90.800 362.200 91.600 367.000 ;
        RECT 94.000 362.200 94.800 367.000 ;
        RECT 99.200 366.800 103.400 367.600 ;
        RECT 105.200 367.400 106.000 373.000 ;
        RECT 114.600 375.200 115.600 376.000 ;
        RECT 114.600 370.800 115.400 375.200 ;
        RECT 116.400 374.600 117.200 379.800 ;
        RECT 122.800 376.600 123.600 379.800 ;
        RECT 124.400 377.000 125.200 379.800 ;
        RECT 126.000 377.000 126.800 379.800 ;
        RECT 127.600 377.000 128.400 379.800 ;
        RECT 129.200 377.000 130.000 379.800 ;
        RECT 132.400 377.000 133.200 379.800 ;
        RECT 135.600 377.000 136.400 379.800 ;
        RECT 137.200 377.000 138.000 379.800 ;
        RECT 138.800 377.000 139.600 379.800 ;
        RECT 121.200 375.800 123.600 376.600 ;
        RECT 140.400 376.600 141.200 379.800 ;
        RECT 121.200 375.200 122.000 375.800 ;
        RECT 116.000 374.000 117.200 374.600 ;
        RECT 120.200 374.600 122.000 375.200 ;
        RECT 126.000 375.600 127.000 376.400 ;
        RECT 130.000 375.600 131.600 376.400 ;
        RECT 132.400 375.800 137.000 376.400 ;
        RECT 140.400 375.800 143.000 376.600 ;
        RECT 132.400 375.600 133.200 375.800 ;
        RECT 116.000 372.000 116.600 374.000 ;
        RECT 120.200 373.400 121.000 374.600 ;
        RECT 117.200 372.600 121.000 373.400 ;
        RECT 126.000 372.800 126.800 375.600 ;
        RECT 132.400 374.800 133.200 375.000 ;
        RECT 128.800 374.200 133.200 374.800 ;
        RECT 128.800 374.000 129.600 374.200 ;
        RECT 134.000 373.600 134.800 375.200 ;
        RECT 136.200 373.400 137.000 375.800 ;
        RECT 142.200 375.200 143.000 375.800 ;
        RECT 142.200 374.400 145.200 375.200 ;
        RECT 146.800 373.800 147.600 379.800 ;
        RECT 129.200 372.600 132.400 373.400 ;
        RECT 136.200 372.600 138.200 373.400 ;
        RECT 138.800 373.000 147.600 373.800 ;
        RECT 122.800 372.000 123.600 372.600 ;
        RECT 140.400 372.000 141.200 372.400 ;
        RECT 145.400 372.000 146.200 372.200 ;
        RECT 116.000 371.400 116.800 372.000 ;
        RECT 122.800 371.400 146.200 372.000 ;
        RECT 114.600 370.000 115.600 370.800 ;
        RECT 104.000 366.800 106.000 367.400 ;
        RECT 95.600 362.200 96.400 365.000 ;
        RECT 97.200 362.200 98.000 365.000 ;
        RECT 100.400 362.200 101.200 366.800 ;
        RECT 104.000 366.200 104.600 366.800 ;
        RECT 103.600 365.600 104.600 366.200 ;
        RECT 103.600 362.200 104.400 365.600 ;
        RECT 114.800 362.200 115.600 370.000 ;
        RECT 116.200 369.600 116.800 371.400 ;
        RECT 116.200 369.000 125.200 369.600 ;
        RECT 116.200 367.400 116.800 369.000 ;
        RECT 124.400 368.800 125.200 369.000 ;
        RECT 127.600 369.000 136.200 369.600 ;
        RECT 127.600 368.800 128.400 369.000 ;
        RECT 119.400 367.600 122.000 368.400 ;
        RECT 116.200 366.800 118.800 367.400 ;
        RECT 118.000 362.200 118.800 366.800 ;
        RECT 121.200 362.200 122.000 367.600 ;
        RECT 122.600 366.800 126.800 367.600 ;
        RECT 124.400 362.200 125.200 365.000 ;
        RECT 126.000 362.200 126.800 365.000 ;
        RECT 127.600 362.200 128.400 365.000 ;
        RECT 129.200 362.200 130.000 368.400 ;
        RECT 132.400 367.600 135.000 368.400 ;
        RECT 135.600 368.200 136.200 369.000 ;
        RECT 137.200 369.400 138.000 369.600 ;
        RECT 137.200 369.000 142.600 369.400 ;
        RECT 137.200 368.800 143.400 369.000 ;
        RECT 142.000 368.200 143.400 368.800 ;
        RECT 135.600 367.600 141.400 368.200 ;
        RECT 144.400 368.000 146.000 368.800 ;
        RECT 144.400 367.600 145.000 368.000 ;
        RECT 132.400 362.200 133.200 367.000 ;
        RECT 135.600 362.200 136.400 367.000 ;
        RECT 140.800 366.800 145.000 367.600 ;
        RECT 146.800 367.400 147.600 373.000 ;
        RECT 145.600 366.800 147.600 367.400 ;
        RECT 148.400 373.800 149.200 379.800 ;
        RECT 154.800 376.600 155.600 379.800 ;
        RECT 156.400 377.000 157.200 379.800 ;
        RECT 158.000 377.000 158.800 379.800 ;
        RECT 159.600 377.000 160.400 379.800 ;
        RECT 162.800 377.000 163.600 379.800 ;
        RECT 166.000 377.000 166.800 379.800 ;
        RECT 167.600 377.000 168.400 379.800 ;
        RECT 169.200 377.000 170.000 379.800 ;
        RECT 170.800 377.000 171.600 379.800 ;
        RECT 153.000 375.800 155.600 376.600 ;
        RECT 172.400 376.600 173.200 379.800 ;
        RECT 159.000 375.800 163.600 376.400 ;
        RECT 153.000 375.200 153.800 375.800 ;
        RECT 150.800 374.400 153.800 375.200 ;
        RECT 148.400 373.000 157.200 373.800 ;
        RECT 159.000 373.400 159.800 375.800 ;
        RECT 162.800 375.600 163.600 375.800 ;
        RECT 164.400 375.600 166.000 376.400 ;
        RECT 169.000 375.600 170.000 376.400 ;
        RECT 172.400 375.800 174.800 376.600 ;
        RECT 161.200 373.600 162.000 375.200 ;
        RECT 162.800 374.800 163.600 375.000 ;
        RECT 162.800 374.200 167.200 374.800 ;
        RECT 166.400 374.000 167.200 374.200 ;
        RECT 148.400 367.400 149.200 373.000 ;
        RECT 157.800 372.600 159.800 373.400 ;
        RECT 163.600 372.600 166.800 373.400 ;
        RECT 169.200 372.800 170.000 375.600 ;
        RECT 174.000 375.200 174.800 375.800 ;
        RECT 174.000 374.600 175.800 375.200 ;
        RECT 175.000 373.400 175.800 374.600 ;
        RECT 178.800 374.600 179.600 379.800 ;
        RECT 180.400 376.000 181.200 379.800 ;
        RECT 180.400 375.200 181.400 376.000 ;
        RECT 178.800 374.000 180.000 374.600 ;
        RECT 175.000 372.600 178.800 373.400 ;
        RECT 149.800 372.000 150.600 372.200 ;
        RECT 153.200 372.000 154.000 372.400 ;
        RECT 154.800 372.000 155.600 372.400 ;
        RECT 172.400 372.000 173.200 372.600 ;
        RECT 179.400 372.000 180.000 374.000 ;
        RECT 149.800 371.400 173.200 372.000 ;
        RECT 179.200 371.400 180.000 372.000 ;
        RECT 179.200 369.600 179.800 371.400 ;
        RECT 180.600 370.800 181.400 375.200 ;
        RECT 158.000 369.400 158.800 369.600 ;
        RECT 153.400 369.000 158.800 369.400 ;
        RECT 152.600 368.800 158.800 369.000 ;
        RECT 159.800 369.000 168.400 369.600 ;
        RECT 150.000 368.000 151.600 368.800 ;
        RECT 152.600 368.200 154.000 368.800 ;
        RECT 159.800 368.200 160.400 369.000 ;
        RECT 167.600 368.800 168.400 369.000 ;
        RECT 170.800 369.000 179.800 369.600 ;
        RECT 170.800 368.800 171.600 369.000 ;
        RECT 151.000 367.600 151.600 368.000 ;
        RECT 154.600 367.600 160.400 368.200 ;
        RECT 161.000 367.600 163.600 368.400 ;
        RECT 148.400 366.800 150.400 367.400 ;
        RECT 151.000 366.800 155.200 367.600 ;
        RECT 137.200 362.200 138.000 365.000 ;
        RECT 138.800 362.200 139.600 365.000 ;
        RECT 142.000 362.200 142.800 366.800 ;
        RECT 145.600 366.200 146.200 366.800 ;
        RECT 145.200 365.600 146.200 366.200 ;
        RECT 149.800 366.200 150.400 366.800 ;
        RECT 149.800 365.600 150.800 366.200 ;
        RECT 145.200 362.200 146.000 365.600 ;
        RECT 150.000 362.200 150.800 365.600 ;
        RECT 153.200 362.200 154.000 366.800 ;
        RECT 156.400 362.200 157.200 365.000 ;
        RECT 158.000 362.200 158.800 365.000 ;
        RECT 159.600 362.200 160.400 367.000 ;
        RECT 162.800 362.200 163.600 367.000 ;
        RECT 166.000 362.200 166.800 368.400 ;
        RECT 174.000 367.600 176.600 368.400 ;
        RECT 169.200 366.800 173.400 367.600 ;
        RECT 167.600 362.200 168.400 365.000 ;
        RECT 169.200 362.200 170.000 365.000 ;
        RECT 170.800 362.200 171.600 365.000 ;
        RECT 174.000 362.200 174.800 367.600 ;
        RECT 179.200 367.400 179.800 369.000 ;
        RECT 177.200 366.800 179.800 367.400 ;
        RECT 180.400 370.000 181.400 370.800 ;
        RECT 183.600 373.800 184.400 379.800 ;
        RECT 190.000 376.600 190.800 379.800 ;
        RECT 191.600 377.000 192.400 379.800 ;
        RECT 193.200 377.000 194.000 379.800 ;
        RECT 194.800 377.000 195.600 379.800 ;
        RECT 198.000 377.000 198.800 379.800 ;
        RECT 201.200 377.000 202.000 379.800 ;
        RECT 202.800 377.000 203.600 379.800 ;
        RECT 204.400 377.000 205.200 379.800 ;
        RECT 206.000 377.000 206.800 379.800 ;
        RECT 188.200 375.800 190.800 376.600 ;
        RECT 207.600 376.600 208.400 379.800 ;
        RECT 194.200 375.800 198.800 376.400 ;
        RECT 188.200 375.200 189.000 375.800 ;
        RECT 186.000 374.400 189.000 375.200 ;
        RECT 183.600 373.000 192.400 373.800 ;
        RECT 194.200 373.400 195.000 375.800 ;
        RECT 198.000 375.600 198.800 375.800 ;
        RECT 199.600 375.600 201.200 376.400 ;
        RECT 204.200 375.600 205.200 376.400 ;
        RECT 207.600 375.800 210.000 376.600 ;
        RECT 196.400 373.600 197.200 375.200 ;
        RECT 198.000 374.800 198.800 375.000 ;
        RECT 198.000 374.200 202.400 374.800 ;
        RECT 201.600 374.000 202.400 374.200 ;
        RECT 180.400 368.300 181.200 370.000 ;
        RECT 182.000 368.300 182.800 368.400 ;
        RECT 180.400 367.700 182.800 368.300 ;
        RECT 177.200 362.200 178.000 366.800 ;
        RECT 180.400 362.200 181.200 367.700 ;
        RECT 182.000 367.600 182.800 367.700 ;
        RECT 183.600 367.400 184.400 373.000 ;
        RECT 193.000 372.600 195.000 373.400 ;
        RECT 198.800 372.600 202.000 373.400 ;
        RECT 204.400 372.800 205.200 375.600 ;
        RECT 209.200 375.200 210.000 375.800 ;
        RECT 209.200 374.600 211.000 375.200 ;
        RECT 210.200 373.400 211.000 374.600 ;
        RECT 214.000 374.600 214.800 379.800 ;
        RECT 215.600 376.000 216.400 379.800 ;
        RECT 219.400 378.400 220.200 379.800 ;
        RECT 218.800 377.600 220.200 378.400 ;
        RECT 219.400 376.400 220.200 377.600 ;
        RECT 215.600 375.200 216.600 376.000 ;
        RECT 219.400 375.800 221.200 376.400 ;
        RECT 223.600 375.800 224.400 379.800 ;
        RECT 225.200 376.000 226.000 379.800 ;
        RECT 228.400 376.000 229.200 379.800 ;
        RECT 225.200 375.800 229.200 376.000 ;
        RECT 230.000 375.800 230.800 379.800 ;
        RECT 231.600 376.000 232.400 379.800 ;
        RECT 234.800 376.000 235.600 379.800 ;
        RECT 231.600 375.800 235.600 376.000 ;
        RECT 237.000 376.400 237.800 379.800 ;
        RECT 237.000 375.800 238.800 376.400 ;
        RECT 241.200 375.800 242.000 379.800 ;
        RECT 242.800 376.000 243.600 379.800 ;
        RECT 246.000 376.000 246.800 379.800 ;
        RECT 250.200 376.400 251.000 379.800 ;
        RECT 242.800 375.800 246.800 376.000 ;
        RECT 249.200 375.800 251.000 376.400 ;
        RECT 254.000 376.000 254.800 379.800 ;
        RECT 214.000 374.000 215.200 374.600 ;
        RECT 210.200 372.600 214.000 373.400 ;
        RECT 185.000 372.000 185.800 372.200 ;
        RECT 186.800 372.000 187.600 372.400 ;
        RECT 190.000 372.000 190.800 372.400 ;
        RECT 207.600 372.000 208.400 372.600 ;
        RECT 214.600 372.000 215.200 374.000 ;
        RECT 185.000 371.400 208.400 372.000 ;
        RECT 214.400 371.400 215.200 372.000 ;
        RECT 214.400 369.600 215.000 371.400 ;
        RECT 215.800 370.800 216.600 375.200 ;
        RECT 193.200 369.400 194.000 369.600 ;
        RECT 188.600 369.000 194.000 369.400 ;
        RECT 187.800 368.800 194.000 369.000 ;
        RECT 195.000 369.000 203.600 369.600 ;
        RECT 185.200 368.000 186.800 368.800 ;
        RECT 187.800 368.200 189.200 368.800 ;
        RECT 195.000 368.200 195.600 369.000 ;
        RECT 202.800 368.800 203.600 369.000 ;
        RECT 206.000 369.000 215.000 369.600 ;
        RECT 206.000 368.800 206.800 369.000 ;
        RECT 186.200 367.600 186.800 368.000 ;
        RECT 189.800 367.600 195.600 368.200 ;
        RECT 196.200 367.600 198.800 368.400 ;
        RECT 183.600 366.800 185.600 367.400 ;
        RECT 186.200 366.800 190.400 367.600 ;
        RECT 185.000 366.200 185.600 366.800 ;
        RECT 185.000 365.600 186.000 366.200 ;
        RECT 185.200 362.200 186.000 365.600 ;
        RECT 188.400 362.200 189.200 366.800 ;
        RECT 191.600 362.200 192.400 365.000 ;
        RECT 193.200 362.200 194.000 365.000 ;
        RECT 194.800 362.200 195.600 367.000 ;
        RECT 198.000 362.200 198.800 367.000 ;
        RECT 201.200 362.200 202.000 368.400 ;
        RECT 209.200 367.600 211.800 368.400 ;
        RECT 204.400 366.800 208.600 367.600 ;
        RECT 202.800 362.200 203.600 365.000 ;
        RECT 204.400 362.200 205.200 365.000 ;
        RECT 206.000 362.200 206.800 365.000 ;
        RECT 209.200 362.200 210.000 367.600 ;
        RECT 214.400 367.400 215.000 369.000 ;
        RECT 212.400 366.800 215.000 367.400 ;
        RECT 215.600 370.000 216.600 370.800 ;
        RECT 212.400 362.200 213.200 366.800 ;
        RECT 215.600 362.200 216.400 370.000 ;
        RECT 218.800 368.800 219.600 370.400 ;
        RECT 220.400 362.200 221.200 375.800 ;
        RECT 222.000 374.300 222.800 375.200 ;
        RECT 223.800 374.400 224.400 375.800 ;
        RECT 225.400 375.400 229.000 375.800 ;
        RECT 227.600 374.400 228.400 374.800 ;
        RECT 230.200 374.400 230.800 375.800 ;
        RECT 231.800 375.400 235.400 375.800 ;
        RECT 234.000 374.400 234.800 374.800 ;
        RECT 223.600 374.300 226.200 374.400 ;
        RECT 222.000 373.700 226.200 374.300 ;
        RECT 227.600 373.800 229.200 374.400 ;
        RECT 222.000 373.600 222.800 373.700 ;
        RECT 223.600 373.600 226.200 373.700 ;
        RECT 228.400 373.600 229.200 373.800 ;
        RECT 230.000 373.600 232.600 374.400 ;
        RECT 234.000 373.800 235.600 374.400 ;
        RECT 234.800 373.600 235.600 373.800 ;
        RECT 236.400 374.300 237.200 374.400 ;
        RECT 238.000 374.300 238.800 375.800 ;
        RECT 236.400 373.700 238.800 374.300 ;
        RECT 236.400 373.600 237.200 373.700 ;
        RECT 222.000 370.300 222.800 370.400 ;
        RECT 223.600 370.300 224.400 370.400 ;
        RECT 222.000 370.200 224.400 370.300 ;
        RECT 225.600 370.200 226.200 373.600 ;
        RECT 226.800 371.600 227.600 373.200 ;
        RECT 230.000 370.200 230.800 370.400 ;
        RECT 232.000 370.200 232.600 373.600 ;
        RECT 233.200 371.600 234.000 373.200 ;
        RECT 222.000 369.700 225.000 370.200 ;
        RECT 222.000 369.600 222.800 369.700 ;
        RECT 223.600 369.600 225.000 369.700 ;
        RECT 225.600 369.600 226.600 370.200 ;
        RECT 230.000 369.600 231.400 370.200 ;
        RECT 232.000 369.600 233.000 370.200 ;
        RECT 224.400 368.400 225.000 369.600 ;
        RECT 224.400 367.600 225.200 368.400 ;
        RECT 225.800 362.200 226.600 369.600 ;
        RECT 230.800 368.400 231.400 369.600 ;
        RECT 232.200 368.400 233.000 369.600 ;
        RECT 236.400 368.800 237.200 370.400 ;
        RECT 230.000 367.600 231.600 368.400 ;
        RECT 232.200 367.600 234.000 368.400 ;
        RECT 232.200 362.200 233.000 367.600 ;
        RECT 238.000 362.200 238.800 373.700 ;
        RECT 239.600 373.600 240.400 375.200 ;
        RECT 241.400 374.400 242.000 375.800 ;
        RECT 243.000 375.400 246.600 375.800 ;
        RECT 245.200 374.400 246.000 374.800 ;
        RECT 241.200 373.600 243.800 374.400 ;
        RECT 245.200 373.800 246.800 374.400 ;
        RECT 246.000 373.600 246.800 373.800 ;
        RECT 247.600 373.600 248.400 375.200 ;
        RECT 241.200 370.200 242.000 370.400 ;
        RECT 243.200 370.200 243.800 373.600 ;
        RECT 244.400 371.600 245.200 373.200 ;
        RECT 241.200 369.600 242.600 370.200 ;
        RECT 243.200 369.600 244.200 370.200 ;
        RECT 242.000 368.400 242.600 369.600 ;
        RECT 239.600 368.300 240.400 368.400 ;
        RECT 242.000 368.300 242.800 368.400 ;
        RECT 239.600 367.700 242.800 368.300 ;
        RECT 239.600 367.600 240.400 367.700 ;
        RECT 242.000 367.600 242.800 367.700 ;
        RECT 243.400 362.200 244.200 369.600 ;
        RECT 249.200 362.200 250.000 375.800 ;
        RECT 253.800 375.200 254.800 376.000 ;
        RECT 253.800 370.800 254.600 375.200 ;
        RECT 255.600 374.600 256.400 379.800 ;
        RECT 262.000 376.600 262.800 379.800 ;
        RECT 263.600 377.000 264.400 379.800 ;
        RECT 265.200 377.000 266.000 379.800 ;
        RECT 266.800 377.000 267.600 379.800 ;
        RECT 268.400 377.000 269.200 379.800 ;
        RECT 271.600 377.000 272.400 379.800 ;
        RECT 274.800 377.000 275.600 379.800 ;
        RECT 276.400 377.000 277.200 379.800 ;
        RECT 278.000 377.000 278.800 379.800 ;
        RECT 260.400 375.800 262.800 376.600 ;
        RECT 279.600 376.600 280.400 379.800 ;
        RECT 260.400 375.200 261.200 375.800 ;
        RECT 255.200 374.000 256.400 374.600 ;
        RECT 259.400 374.600 261.200 375.200 ;
        RECT 265.200 375.600 266.200 376.400 ;
        RECT 269.200 375.600 270.800 376.400 ;
        RECT 271.600 375.800 276.200 376.400 ;
        RECT 279.600 375.800 282.200 376.600 ;
        RECT 271.600 375.600 272.400 375.800 ;
        RECT 255.200 372.000 255.800 374.000 ;
        RECT 259.400 373.400 260.200 374.600 ;
        RECT 256.400 372.600 260.200 373.400 ;
        RECT 265.200 372.800 266.000 375.600 ;
        RECT 271.600 374.800 272.400 375.000 ;
        RECT 268.000 374.200 272.400 374.800 ;
        RECT 268.000 374.000 268.800 374.200 ;
        RECT 273.200 373.600 274.000 375.200 ;
        RECT 275.400 373.400 276.200 375.800 ;
        RECT 281.400 375.200 282.200 375.800 ;
        RECT 281.400 374.400 284.400 375.200 ;
        RECT 286.000 373.800 286.800 379.800 ;
        RECT 294.000 375.800 294.800 379.800 ;
        RECT 295.600 376.000 296.400 379.800 ;
        RECT 298.800 376.000 299.600 379.800 ;
        RECT 303.000 376.400 303.800 379.800 ;
        RECT 295.600 375.800 299.600 376.000 ;
        RECT 302.000 375.800 303.800 376.400 ;
        RECT 294.200 374.400 294.800 375.800 ;
        RECT 295.800 375.400 299.400 375.800 ;
        RECT 298.000 374.400 298.800 374.800 ;
        RECT 268.400 372.600 271.600 373.400 ;
        RECT 275.400 372.600 277.400 373.400 ;
        RECT 278.000 373.000 286.800 373.800 ;
        RECT 294.000 373.600 296.600 374.400 ;
        RECT 298.000 373.800 299.600 374.400 ;
        RECT 298.800 373.600 299.600 373.800 ;
        RECT 300.400 373.600 301.200 375.200 ;
        RECT 262.000 372.000 262.800 372.600 ;
        RECT 279.600 372.000 280.400 372.400 ;
        RECT 281.200 372.000 282.000 372.400 ;
        RECT 284.600 372.000 285.400 372.200 ;
        RECT 255.200 371.400 256.000 372.000 ;
        RECT 262.000 371.400 285.400 372.000 ;
        RECT 250.800 368.800 251.600 370.400 ;
        RECT 253.800 370.000 254.800 370.800 ;
        RECT 254.000 362.200 254.800 370.000 ;
        RECT 255.400 369.600 256.000 371.400 ;
        RECT 255.400 369.000 264.400 369.600 ;
        RECT 255.400 367.400 256.000 369.000 ;
        RECT 263.600 368.800 264.400 369.000 ;
        RECT 266.800 369.000 275.400 369.600 ;
        RECT 266.800 368.800 267.600 369.000 ;
        RECT 258.600 367.600 261.200 368.400 ;
        RECT 255.400 366.800 258.000 367.400 ;
        RECT 257.200 362.200 258.000 366.800 ;
        RECT 260.400 362.200 261.200 367.600 ;
        RECT 261.800 366.800 266.000 367.600 ;
        RECT 263.600 362.200 264.400 365.000 ;
        RECT 265.200 362.200 266.000 365.000 ;
        RECT 266.800 362.200 267.600 365.000 ;
        RECT 268.400 362.200 269.200 368.400 ;
        RECT 271.600 367.600 274.200 368.400 ;
        RECT 274.800 368.200 275.400 369.000 ;
        RECT 276.400 369.400 277.200 369.600 ;
        RECT 276.400 369.000 281.800 369.400 ;
        RECT 276.400 368.800 282.600 369.000 ;
        RECT 281.200 368.200 282.600 368.800 ;
        RECT 274.800 367.600 280.600 368.200 ;
        RECT 283.600 368.000 285.200 368.800 ;
        RECT 283.600 367.600 284.200 368.000 ;
        RECT 271.600 362.200 272.400 367.000 ;
        RECT 274.800 362.200 275.600 367.000 ;
        RECT 280.000 366.800 284.200 367.600 ;
        RECT 286.000 367.400 286.800 373.000 ;
        RECT 294.000 370.200 294.800 370.400 ;
        RECT 296.000 370.200 296.600 373.600 ;
        RECT 297.200 371.600 298.000 373.200 ;
        RECT 294.000 369.600 295.400 370.200 ;
        RECT 296.000 369.600 297.000 370.200 ;
        RECT 294.800 368.400 295.400 369.600 ;
        RECT 292.400 368.300 293.200 368.400 ;
        RECT 294.800 368.300 295.600 368.400 ;
        RECT 292.400 367.700 295.600 368.300 ;
        RECT 292.400 367.600 293.200 367.700 ;
        RECT 294.800 367.600 295.600 367.700 ;
        RECT 284.800 366.800 286.800 367.400 ;
        RECT 276.400 362.200 277.200 365.000 ;
        RECT 278.000 362.200 278.800 365.000 ;
        RECT 281.200 362.200 282.000 366.800 ;
        RECT 284.800 366.200 285.400 366.800 ;
        RECT 284.400 365.600 285.400 366.200 ;
        RECT 284.400 362.200 285.200 365.600 ;
        RECT 296.200 362.200 297.000 369.600 ;
        RECT 302.000 362.200 302.800 375.800 ;
        RECT 303.600 368.800 304.400 370.400 ;
        RECT 305.200 362.200 306.000 379.800 ;
        RECT 306.800 373.600 307.600 375.200 ;
        RECT 312.000 374.200 312.800 379.800 ;
        RECT 316.400 377.800 317.200 379.800 ;
        RECT 314.800 375.600 315.600 377.200 ;
        RECT 316.600 374.400 317.200 377.800 ;
        RECT 319.600 376.000 320.400 379.800 ;
        RECT 322.800 376.000 323.600 379.800 ;
        RECT 319.600 375.800 323.600 376.000 ;
        RECT 324.400 375.800 325.200 379.800 ;
        RECT 319.800 375.400 323.400 375.800 ;
        RECT 320.400 374.400 321.200 374.800 ;
        RECT 324.400 374.400 325.000 375.800 ;
        RECT 312.000 373.800 313.800 374.200 ;
        RECT 312.200 373.600 313.800 373.800 ;
        RECT 316.400 373.600 317.200 374.400 ;
        RECT 319.600 373.800 321.200 374.400 ;
        RECT 319.600 373.600 320.400 373.800 ;
        RECT 322.600 373.600 325.200 374.400 ;
        RECT 329.600 374.200 330.400 379.800 ;
        RECT 333.000 376.400 333.800 379.800 ;
        RECT 337.800 376.400 338.600 379.800 ;
        RECT 342.600 378.400 343.400 379.800 ;
        RECT 342.000 377.600 343.400 378.400 ;
        RECT 342.600 376.800 343.400 377.600 ;
        RECT 333.000 375.800 334.800 376.400 ;
        RECT 337.800 375.800 339.600 376.400 ;
        RECT 329.600 373.800 331.400 374.200 ;
        RECT 329.800 373.600 331.400 373.800 ;
        RECT 310.000 371.600 311.600 372.400 ;
        RECT 308.400 369.600 309.200 371.200 ;
        RECT 313.200 370.400 313.800 373.600 ;
        RECT 314.800 372.300 315.600 372.400 ;
        RECT 316.600 372.300 317.200 373.600 ;
        RECT 314.800 371.700 317.200 372.300 ;
        RECT 314.800 371.600 315.600 371.700 ;
        RECT 313.200 369.600 314.000 370.400 ;
        RECT 316.600 370.200 317.200 371.700 ;
        RECT 318.000 370.800 318.800 372.400 ;
        RECT 319.600 372.300 320.400 372.400 ;
        RECT 321.200 372.300 322.000 373.200 ;
        RECT 319.600 371.700 322.000 372.300 ;
        RECT 319.600 371.600 320.400 371.700 ;
        RECT 321.200 371.600 322.000 371.700 ;
        RECT 322.600 372.400 323.200 373.600 ;
        RECT 322.600 371.600 323.600 372.400 ;
        RECT 327.600 371.600 329.200 372.400 ;
        RECT 322.600 370.200 323.200 371.600 ;
        RECT 324.400 370.300 325.200 370.400 ;
        RECT 326.000 370.300 326.800 371.200 ;
        RECT 324.400 370.200 326.800 370.300 ;
        RECT 310.000 368.300 310.800 368.400 ;
        RECT 311.600 368.300 312.400 369.200 ;
        RECT 310.000 367.700 312.400 368.300 ;
        RECT 310.000 367.600 310.800 367.700 ;
        RECT 311.600 367.600 312.400 367.700 ;
        RECT 313.200 368.400 313.800 369.600 ;
        RECT 316.400 369.400 318.200 370.200 ;
        RECT 313.200 367.600 314.000 368.400 ;
        RECT 313.200 367.000 313.800 367.600 ;
        RECT 310.200 366.400 313.800 367.000 ;
        RECT 310.200 366.200 310.800 366.400 ;
        RECT 310.000 362.200 310.800 366.200 ;
        RECT 313.200 366.200 313.800 366.400 ;
        RECT 313.200 362.200 314.000 366.200 ;
        RECT 317.400 362.200 318.200 369.400 ;
        RECT 322.200 369.600 323.200 370.200 ;
        RECT 323.800 369.700 326.800 370.200 ;
        RECT 323.800 369.600 325.200 369.700 ;
        RECT 326.000 369.600 326.800 369.700 ;
        RECT 330.800 370.400 331.400 373.600 ;
        RECT 330.800 369.600 331.600 370.400 ;
        RECT 322.200 362.200 323.000 369.600 ;
        RECT 323.800 368.400 324.400 369.600 ;
        RECT 323.600 367.600 324.400 368.400 ;
        RECT 329.200 367.600 330.000 369.200 ;
        RECT 330.800 367.000 331.400 369.600 ;
        RECT 332.400 368.800 333.200 370.400 ;
        RECT 327.800 366.400 331.400 367.000 ;
        RECT 327.600 362.200 328.400 366.400 ;
        RECT 330.800 366.200 331.400 366.400 ;
        RECT 330.800 362.200 331.600 366.200 ;
        RECT 334.000 362.200 334.800 375.800 ;
        RECT 335.600 373.600 336.400 375.200 ;
        RECT 337.200 374.300 338.000 374.400 ;
        RECT 338.800 374.300 339.600 375.800 ;
        RECT 342.000 375.800 343.400 376.800 ;
        RECT 346.800 375.800 347.600 379.800 ;
        RECT 337.200 373.700 339.600 374.300 ;
        RECT 337.200 373.600 338.000 373.700 ;
        RECT 337.200 368.800 338.000 370.400 ;
        RECT 338.800 362.200 339.600 373.700 ;
        RECT 340.400 373.600 341.200 375.200 ;
        RECT 342.000 372.400 342.600 375.800 ;
        RECT 346.800 375.600 347.400 375.800 ;
        RECT 345.600 375.200 347.400 375.600 ;
        RECT 343.200 375.000 347.400 375.200 ;
        RECT 343.200 374.600 346.200 375.000 ;
        RECT 343.200 374.400 344.000 374.600 ;
        RECT 342.000 371.600 342.800 372.400 ;
        RECT 342.000 370.200 342.600 371.600 ;
        RECT 343.400 371.000 344.000 374.400 ;
        RECT 344.800 373.800 345.600 374.000 ;
        RECT 344.800 373.200 345.800 373.800 ;
        RECT 345.200 372.400 345.800 373.200 ;
        RECT 346.800 372.800 347.600 374.400 ;
        RECT 348.400 373.800 349.200 379.800 ;
        RECT 354.800 376.600 355.600 379.800 ;
        RECT 356.400 377.000 357.200 379.800 ;
        RECT 358.000 377.000 358.800 379.800 ;
        RECT 359.600 377.000 360.400 379.800 ;
        RECT 362.800 377.000 363.600 379.800 ;
        RECT 366.000 377.000 366.800 379.800 ;
        RECT 367.600 377.000 368.400 379.800 ;
        RECT 369.200 377.000 370.000 379.800 ;
        RECT 370.800 377.000 371.600 379.800 ;
        RECT 353.000 375.800 355.600 376.600 ;
        RECT 372.400 376.600 373.200 379.800 ;
        RECT 359.000 375.800 363.600 376.400 ;
        RECT 353.000 375.200 353.800 375.800 ;
        RECT 350.800 374.400 353.800 375.200 ;
        RECT 348.400 373.000 357.200 373.800 ;
        RECT 359.000 373.400 359.800 375.800 ;
        RECT 362.800 375.600 363.600 375.800 ;
        RECT 364.400 375.600 366.000 376.400 ;
        RECT 369.000 375.600 370.000 376.400 ;
        RECT 372.400 375.800 374.800 376.600 ;
        RECT 361.200 373.600 362.000 375.200 ;
        RECT 362.800 374.800 363.600 375.000 ;
        RECT 362.800 374.200 367.200 374.800 ;
        RECT 366.400 374.000 367.200 374.200 ;
        RECT 345.200 371.600 346.000 372.400 ;
        RECT 343.400 370.400 345.800 371.000 ;
        RECT 342.000 362.200 342.800 370.200 ;
        RECT 345.200 366.200 345.800 370.400 ;
        RECT 348.400 367.400 349.200 373.000 ;
        RECT 357.800 372.600 359.800 373.400 ;
        RECT 363.600 372.600 366.800 373.400 ;
        RECT 369.200 372.800 370.000 375.600 ;
        RECT 374.000 375.200 374.800 375.800 ;
        RECT 374.000 374.600 375.800 375.200 ;
        RECT 375.000 373.400 375.800 374.600 ;
        RECT 378.800 374.600 379.600 379.800 ;
        RECT 380.400 376.300 381.200 379.800 ;
        RECT 385.200 377.800 386.000 379.800 ;
        RECT 383.600 376.300 384.400 377.200 ;
        RECT 380.400 375.700 384.400 376.300 ;
        RECT 380.400 375.200 381.400 375.700 ;
        RECT 383.600 375.600 384.400 375.700 ;
        RECT 378.800 374.000 380.000 374.600 ;
        RECT 375.000 372.600 378.800 373.400 ;
        RECT 379.400 372.000 380.000 374.000 ;
        RECT 379.200 371.400 380.000 372.000 ;
        RECT 377.800 370.800 378.600 371.000 ;
        RECT 351.600 370.200 378.600 370.800 ;
        RECT 351.600 369.600 352.400 370.200 ;
        RECT 355.000 370.000 355.800 370.200 ;
        RECT 379.200 369.600 379.800 371.400 ;
        RECT 380.600 370.800 381.400 375.200 ;
        RECT 385.400 374.400 386.000 377.800 ;
        RECT 388.400 375.800 389.200 379.800 ;
        RECT 390.000 376.000 390.800 379.800 ;
        RECT 393.200 376.000 394.000 379.800 ;
        RECT 390.000 375.800 394.000 376.000 ;
        RECT 388.600 374.400 389.200 375.800 ;
        RECT 390.200 375.400 393.800 375.800 ;
        RECT 392.400 374.400 393.200 374.800 ;
        RECT 385.200 373.600 386.000 374.400 ;
        RECT 388.400 373.600 391.000 374.400 ;
        RECT 392.400 373.800 394.000 374.400 ;
        RECT 393.200 373.600 394.000 373.800 ;
        RECT 394.800 373.800 395.600 379.800 ;
        RECT 401.200 376.600 402.000 379.800 ;
        RECT 402.800 377.000 403.600 379.800 ;
        RECT 404.400 377.000 405.200 379.800 ;
        RECT 406.000 377.000 406.800 379.800 ;
        RECT 409.200 377.000 410.000 379.800 ;
        RECT 412.400 377.000 413.200 379.800 ;
        RECT 414.000 377.000 414.800 379.800 ;
        RECT 415.600 377.000 416.400 379.800 ;
        RECT 417.200 377.000 418.000 379.800 ;
        RECT 399.400 375.800 402.000 376.600 ;
        RECT 418.800 376.600 419.600 379.800 ;
        RECT 405.400 375.800 410.000 376.400 ;
        RECT 399.400 375.200 400.200 375.800 ;
        RECT 397.200 374.400 400.200 375.200 ;
        RECT 382.000 372.300 382.800 372.400 ;
        RECT 385.400 372.300 386.000 373.600 ;
        RECT 382.000 371.700 386.000 372.300 ;
        RECT 382.000 371.600 382.800 371.700 ;
        RECT 358.000 369.400 358.800 369.600 ;
        RECT 353.400 369.000 358.800 369.400 ;
        RECT 352.600 368.800 358.800 369.000 ;
        RECT 359.800 369.000 368.400 369.600 ;
        RECT 350.000 368.000 351.600 368.800 ;
        RECT 352.600 368.200 354.000 368.800 ;
        RECT 359.800 368.200 360.400 369.000 ;
        RECT 367.600 368.800 368.400 369.000 ;
        RECT 370.800 369.000 379.800 369.600 ;
        RECT 370.800 368.800 371.600 369.000 ;
        RECT 351.000 367.600 351.600 368.000 ;
        RECT 354.600 367.600 360.400 368.200 ;
        RECT 361.000 367.600 363.600 368.400 ;
        RECT 348.400 366.800 350.400 367.400 ;
        RECT 351.000 366.800 355.200 367.600 ;
        RECT 349.800 366.200 350.400 366.800 ;
        RECT 345.200 362.200 346.000 366.200 ;
        RECT 349.800 365.600 350.800 366.200 ;
        RECT 350.000 362.200 350.800 365.600 ;
        RECT 353.200 362.200 354.000 366.800 ;
        RECT 356.400 362.200 357.200 365.000 ;
        RECT 358.000 362.200 358.800 365.000 ;
        RECT 359.600 362.200 360.400 367.000 ;
        RECT 362.800 362.200 363.600 367.000 ;
        RECT 366.000 362.200 366.800 368.400 ;
        RECT 374.000 367.600 376.600 368.400 ;
        RECT 369.200 366.800 373.400 367.600 ;
        RECT 367.600 362.200 368.400 365.000 ;
        RECT 369.200 362.200 370.000 365.000 ;
        RECT 370.800 362.200 371.600 365.000 ;
        RECT 374.000 362.200 374.800 367.600 ;
        RECT 379.200 367.400 379.800 369.000 ;
        RECT 377.200 366.800 379.800 367.400 ;
        RECT 380.400 370.000 381.400 370.800 ;
        RECT 385.400 370.200 386.000 371.700 ;
        RECT 386.800 370.800 387.600 372.400 ;
        RECT 388.400 370.200 389.200 370.400 ;
        RECT 390.400 370.200 391.000 373.600 ;
        RECT 391.600 371.600 392.400 373.200 ;
        RECT 394.800 373.000 403.600 373.800 ;
        RECT 405.400 373.400 406.200 375.800 ;
        RECT 409.200 375.600 410.000 375.800 ;
        RECT 410.800 375.600 412.400 376.400 ;
        RECT 415.400 375.600 416.400 376.400 ;
        RECT 418.800 375.800 421.200 376.600 ;
        RECT 407.600 373.600 408.400 375.200 ;
        RECT 409.200 374.800 410.000 375.000 ;
        RECT 409.200 374.200 413.600 374.800 ;
        RECT 412.800 374.000 413.600 374.200 ;
        RECT 377.200 362.200 378.000 366.800 ;
        RECT 380.400 362.200 381.200 370.000 ;
        RECT 385.200 369.400 387.000 370.200 ;
        RECT 388.400 369.600 389.800 370.200 ;
        RECT 390.400 369.600 391.400 370.200 ;
        RECT 386.200 362.200 387.000 369.400 ;
        RECT 389.200 368.400 389.800 369.600 ;
        RECT 389.200 367.600 390.000 368.400 ;
        RECT 390.600 362.200 391.400 369.600 ;
        RECT 394.800 367.400 395.600 373.000 ;
        RECT 404.200 372.600 406.200 373.400 ;
        RECT 410.000 372.600 413.200 373.400 ;
        RECT 415.600 372.800 416.400 375.600 ;
        RECT 420.400 375.200 421.200 375.800 ;
        RECT 420.400 374.600 422.200 375.200 ;
        RECT 421.400 373.400 422.200 374.600 ;
        RECT 425.200 374.600 426.000 379.800 ;
        RECT 426.800 376.000 427.600 379.800 ;
        RECT 438.000 376.000 438.800 379.800 ;
        RECT 426.800 375.200 427.800 376.000 ;
        RECT 425.200 374.000 426.400 374.600 ;
        RECT 421.400 372.600 425.200 373.400 ;
        RECT 396.200 372.000 397.000 372.200 ;
        RECT 399.600 372.000 400.400 372.400 ;
        RECT 401.200 372.000 402.000 372.400 ;
        RECT 418.800 372.000 419.600 372.600 ;
        RECT 425.800 372.000 426.400 374.000 ;
        RECT 396.200 371.400 419.600 372.000 ;
        RECT 425.600 371.400 426.400 372.000 ;
        RECT 425.600 369.600 426.200 371.400 ;
        RECT 427.000 370.800 427.800 375.200 ;
        RECT 404.400 369.400 405.200 369.600 ;
        RECT 399.800 369.000 405.200 369.400 ;
        RECT 399.000 368.800 405.200 369.000 ;
        RECT 406.200 369.000 414.800 369.600 ;
        RECT 396.400 368.000 398.000 368.800 ;
        RECT 399.000 368.200 400.400 368.800 ;
        RECT 406.200 368.200 406.800 369.000 ;
        RECT 414.000 368.800 414.800 369.000 ;
        RECT 417.200 369.000 426.200 369.600 ;
        RECT 417.200 368.800 418.000 369.000 ;
        RECT 397.400 367.600 398.000 368.000 ;
        RECT 401.000 367.600 406.800 368.200 ;
        RECT 407.400 367.600 410.000 368.400 ;
        RECT 394.800 366.800 396.800 367.400 ;
        RECT 397.400 366.800 401.600 367.600 ;
        RECT 396.200 366.200 396.800 366.800 ;
        RECT 396.200 365.600 397.200 366.200 ;
        RECT 396.400 362.200 397.200 365.600 ;
        RECT 399.600 362.200 400.400 366.800 ;
        RECT 402.800 362.200 403.600 365.000 ;
        RECT 404.400 362.200 405.200 365.000 ;
        RECT 406.000 362.200 406.800 367.000 ;
        RECT 409.200 362.200 410.000 367.000 ;
        RECT 412.400 362.200 413.200 368.400 ;
        RECT 420.400 367.600 423.000 368.400 ;
        RECT 415.600 366.800 419.800 367.600 ;
        RECT 414.000 362.200 414.800 365.000 ;
        RECT 415.600 362.200 416.400 365.000 ;
        RECT 417.200 362.200 418.000 365.000 ;
        RECT 420.400 362.200 421.200 367.600 ;
        RECT 425.600 367.400 426.200 369.000 ;
        RECT 423.600 366.800 426.200 367.400 ;
        RECT 426.800 370.000 427.800 370.800 ;
        RECT 437.800 375.200 438.800 376.000 ;
        RECT 437.800 370.800 438.600 375.200 ;
        RECT 439.600 374.600 440.400 379.800 ;
        RECT 446.000 376.600 446.800 379.800 ;
        RECT 447.600 377.000 448.400 379.800 ;
        RECT 449.200 377.000 450.000 379.800 ;
        RECT 450.800 377.000 451.600 379.800 ;
        RECT 452.400 377.000 453.200 379.800 ;
        RECT 455.600 377.000 456.400 379.800 ;
        RECT 458.800 377.000 459.600 379.800 ;
        RECT 460.400 377.000 461.200 379.800 ;
        RECT 462.000 377.000 462.800 379.800 ;
        RECT 444.400 375.800 446.800 376.600 ;
        RECT 463.600 376.600 464.400 379.800 ;
        RECT 444.400 375.200 445.200 375.800 ;
        RECT 439.200 374.000 440.400 374.600 ;
        RECT 443.400 374.600 445.200 375.200 ;
        RECT 449.200 375.600 450.200 376.400 ;
        RECT 453.200 375.600 454.800 376.400 ;
        RECT 455.600 375.800 460.200 376.400 ;
        RECT 463.600 375.800 466.200 376.600 ;
        RECT 455.600 375.600 456.400 375.800 ;
        RECT 439.200 372.000 439.800 374.000 ;
        RECT 443.400 373.400 444.200 374.600 ;
        RECT 440.400 372.600 444.200 373.400 ;
        RECT 449.200 372.800 450.000 375.600 ;
        RECT 455.600 374.800 456.400 375.000 ;
        RECT 452.000 374.200 456.400 374.800 ;
        RECT 452.000 374.000 452.800 374.200 ;
        RECT 457.200 373.600 458.000 375.200 ;
        RECT 459.400 373.400 460.200 375.800 ;
        RECT 465.400 375.200 466.200 375.800 ;
        RECT 465.400 374.400 468.400 375.200 ;
        RECT 470.000 373.800 470.800 379.800 ;
        RECT 452.400 372.600 455.600 373.400 ;
        RECT 459.400 372.600 461.400 373.400 ;
        RECT 462.000 373.000 470.800 373.800 ;
        RECT 446.000 372.000 446.800 372.600 ;
        RECT 463.600 372.000 464.400 372.400 ;
        RECT 468.600 372.000 469.400 372.200 ;
        RECT 439.200 371.400 440.000 372.000 ;
        RECT 446.000 371.400 469.400 372.000 ;
        RECT 437.800 370.000 438.800 370.800 ;
        RECT 423.600 362.200 424.400 366.800 ;
        RECT 426.800 362.200 427.600 370.000 ;
        RECT 438.000 362.200 438.800 370.000 ;
        RECT 439.400 369.600 440.000 371.400 ;
        RECT 439.400 369.000 448.400 369.600 ;
        RECT 439.400 367.400 440.000 369.000 ;
        RECT 447.600 368.800 448.400 369.000 ;
        RECT 450.800 369.000 459.400 369.600 ;
        RECT 450.800 368.800 451.600 369.000 ;
        RECT 442.600 367.600 445.200 368.400 ;
        RECT 439.400 366.800 442.000 367.400 ;
        RECT 441.200 362.200 442.000 366.800 ;
        RECT 444.400 362.200 445.200 367.600 ;
        RECT 445.800 366.800 450.000 367.600 ;
        RECT 447.600 362.200 448.400 365.000 ;
        RECT 449.200 362.200 450.000 365.000 ;
        RECT 450.800 362.200 451.600 365.000 ;
        RECT 452.400 362.200 453.200 368.400 ;
        RECT 455.600 367.600 458.200 368.400 ;
        RECT 458.800 368.200 459.400 369.000 ;
        RECT 460.400 369.400 461.200 369.600 ;
        RECT 460.400 369.000 465.800 369.400 ;
        RECT 460.400 368.800 466.600 369.000 ;
        RECT 465.200 368.200 466.600 368.800 ;
        RECT 458.800 367.600 464.600 368.200 ;
        RECT 467.600 368.000 469.200 368.800 ;
        RECT 467.600 367.600 468.200 368.000 ;
        RECT 455.600 362.200 456.400 367.000 ;
        RECT 458.800 362.200 459.600 367.000 ;
        RECT 464.000 366.800 468.200 367.600 ;
        RECT 470.000 367.400 470.800 373.000 ;
        RECT 468.800 366.800 470.800 367.400 ;
        RECT 471.600 373.800 472.400 379.800 ;
        RECT 478.000 376.600 478.800 379.800 ;
        RECT 479.600 377.000 480.400 379.800 ;
        RECT 481.200 377.000 482.000 379.800 ;
        RECT 482.800 377.000 483.600 379.800 ;
        RECT 486.000 377.000 486.800 379.800 ;
        RECT 489.200 377.000 490.000 379.800 ;
        RECT 490.800 377.000 491.600 379.800 ;
        RECT 492.400 377.000 493.200 379.800 ;
        RECT 494.000 377.000 494.800 379.800 ;
        RECT 476.200 375.800 478.800 376.600 ;
        RECT 495.600 376.600 496.400 379.800 ;
        RECT 482.200 375.800 486.800 376.400 ;
        RECT 476.200 375.200 477.000 375.800 ;
        RECT 474.000 374.400 477.000 375.200 ;
        RECT 471.600 373.000 480.400 373.800 ;
        RECT 482.200 373.400 483.000 375.800 ;
        RECT 486.000 375.600 486.800 375.800 ;
        RECT 487.600 375.600 489.200 376.400 ;
        RECT 492.200 375.600 493.200 376.400 ;
        RECT 495.600 375.800 498.000 376.600 ;
        RECT 484.400 373.600 485.200 375.200 ;
        RECT 486.000 374.800 486.800 375.000 ;
        RECT 486.000 374.200 490.400 374.800 ;
        RECT 489.600 374.000 490.400 374.200 ;
        RECT 471.600 367.400 472.400 373.000 ;
        RECT 481.000 372.600 483.000 373.400 ;
        RECT 486.800 372.600 490.000 373.400 ;
        RECT 492.400 372.800 493.200 375.600 ;
        RECT 497.200 375.200 498.000 375.800 ;
        RECT 497.200 374.600 499.000 375.200 ;
        RECT 498.200 373.400 499.000 374.600 ;
        RECT 502.000 374.600 502.800 379.800 ;
        RECT 503.600 376.000 504.400 379.800 ;
        RECT 509.400 376.400 510.200 379.800 ;
        RECT 503.600 375.200 504.600 376.000 ;
        RECT 508.400 375.800 510.200 376.400 ;
        RECT 513.200 376.000 514.000 379.800 ;
        RECT 502.000 374.000 503.200 374.600 ;
        RECT 498.200 372.600 502.000 373.400 ;
        RECT 473.000 372.000 473.800 372.200 ;
        RECT 474.800 372.000 475.600 372.400 ;
        RECT 478.000 372.000 478.800 372.400 ;
        RECT 495.600 372.000 496.400 372.600 ;
        RECT 502.600 372.000 503.200 374.000 ;
        RECT 473.000 371.400 496.400 372.000 ;
        RECT 502.400 371.400 503.200 372.000 ;
        RECT 502.400 369.600 503.000 371.400 ;
        RECT 503.800 370.800 504.600 375.200 ;
        RECT 506.800 373.600 507.600 375.200 ;
        RECT 481.200 369.400 482.000 369.600 ;
        RECT 476.600 369.000 482.000 369.400 ;
        RECT 475.800 368.800 482.000 369.000 ;
        RECT 483.000 369.000 491.600 369.600 ;
        RECT 473.200 368.000 474.800 368.800 ;
        RECT 475.800 368.200 477.200 368.800 ;
        RECT 483.000 368.200 483.600 369.000 ;
        RECT 490.800 368.800 491.600 369.000 ;
        RECT 494.000 369.000 503.000 369.600 ;
        RECT 494.000 368.800 494.800 369.000 ;
        RECT 474.200 367.600 474.800 368.000 ;
        RECT 477.800 367.600 483.600 368.200 ;
        RECT 484.200 367.600 486.800 368.400 ;
        RECT 471.600 366.800 473.600 367.400 ;
        RECT 474.200 366.800 478.400 367.600 ;
        RECT 460.400 362.200 461.200 365.000 ;
        RECT 462.000 362.200 462.800 365.000 ;
        RECT 465.200 362.200 466.000 366.800 ;
        RECT 468.800 366.200 469.400 366.800 ;
        RECT 468.400 365.600 469.400 366.200 ;
        RECT 473.000 366.200 473.600 366.800 ;
        RECT 473.000 365.600 474.000 366.200 ;
        RECT 468.400 362.200 469.200 365.600 ;
        RECT 473.200 362.200 474.000 365.600 ;
        RECT 476.400 362.200 477.200 366.800 ;
        RECT 479.600 362.200 480.400 365.000 ;
        RECT 481.200 362.200 482.000 365.000 ;
        RECT 482.800 362.200 483.600 367.000 ;
        RECT 486.000 362.200 486.800 367.000 ;
        RECT 489.200 362.200 490.000 368.400 ;
        RECT 497.200 367.600 499.800 368.400 ;
        RECT 492.400 366.800 496.600 367.600 ;
        RECT 490.800 362.200 491.600 365.000 ;
        RECT 492.400 362.200 493.200 365.000 ;
        RECT 494.000 362.200 494.800 365.000 ;
        RECT 497.200 362.200 498.000 367.600 ;
        RECT 502.400 367.400 503.000 369.000 ;
        RECT 500.400 366.800 503.000 367.400 ;
        RECT 503.600 370.000 504.600 370.800 ;
        RECT 500.400 362.200 501.200 366.800 ;
        RECT 503.600 362.200 504.400 370.000 ;
        RECT 506.800 368.300 507.600 368.400 ;
        RECT 508.400 368.300 509.200 375.800 ;
        RECT 513.000 375.200 514.000 376.000 ;
        RECT 513.000 370.800 513.800 375.200 ;
        RECT 514.800 374.600 515.600 379.800 ;
        RECT 521.200 376.600 522.000 379.800 ;
        RECT 522.800 377.000 523.600 379.800 ;
        RECT 524.400 377.000 525.200 379.800 ;
        RECT 526.000 377.000 526.800 379.800 ;
        RECT 527.600 377.000 528.400 379.800 ;
        RECT 530.800 377.000 531.600 379.800 ;
        RECT 534.000 377.000 534.800 379.800 ;
        RECT 535.600 377.000 536.400 379.800 ;
        RECT 537.200 377.000 538.000 379.800 ;
        RECT 519.600 375.800 522.000 376.600 ;
        RECT 538.800 376.600 539.600 379.800 ;
        RECT 519.600 375.200 520.400 375.800 ;
        RECT 514.400 374.000 515.600 374.600 ;
        RECT 518.600 374.600 520.400 375.200 ;
        RECT 524.400 375.600 525.400 376.400 ;
        RECT 528.400 375.600 530.000 376.400 ;
        RECT 530.800 375.800 535.400 376.400 ;
        RECT 538.800 375.800 541.400 376.600 ;
        RECT 530.800 375.600 531.600 375.800 ;
        RECT 514.400 372.000 515.000 374.000 ;
        RECT 518.600 373.400 519.400 374.600 ;
        RECT 515.600 372.600 519.400 373.400 ;
        RECT 524.400 372.800 525.200 375.600 ;
        RECT 530.800 374.800 531.600 375.000 ;
        RECT 527.200 374.200 531.600 374.800 ;
        RECT 527.200 374.000 528.000 374.200 ;
        RECT 532.400 373.600 533.200 375.200 ;
        RECT 534.600 373.400 535.400 375.800 ;
        RECT 540.600 375.200 541.400 375.800 ;
        RECT 540.600 374.400 543.600 375.200 ;
        RECT 545.200 373.800 546.000 379.800 ;
        RECT 527.600 372.600 530.800 373.400 ;
        RECT 534.600 372.600 536.600 373.400 ;
        RECT 537.200 373.000 546.000 373.800 ;
        RECT 521.200 372.000 522.000 372.600 ;
        RECT 538.800 372.000 539.600 372.400 ;
        RECT 542.000 372.000 542.800 372.400 ;
        RECT 543.800 372.000 544.600 372.200 ;
        RECT 514.400 371.400 515.200 372.000 ;
        RECT 521.200 371.400 544.600 372.000 ;
        RECT 510.000 368.800 510.800 370.400 ;
        RECT 513.000 370.000 514.000 370.800 ;
        RECT 506.800 367.700 509.200 368.300 ;
        RECT 506.800 367.600 507.600 367.700 ;
        RECT 508.400 362.200 509.200 367.700 ;
        RECT 513.200 362.200 514.000 370.000 ;
        RECT 514.600 369.600 515.200 371.400 ;
        RECT 514.600 369.000 523.600 369.600 ;
        RECT 514.600 367.400 515.200 369.000 ;
        RECT 522.800 368.800 523.600 369.000 ;
        RECT 526.000 369.000 534.600 369.600 ;
        RECT 526.000 368.800 526.800 369.000 ;
        RECT 517.800 367.600 520.400 368.400 ;
        RECT 514.600 366.800 517.200 367.400 ;
        RECT 516.400 362.200 517.200 366.800 ;
        RECT 519.600 362.200 520.400 367.600 ;
        RECT 521.000 366.800 525.200 367.600 ;
        RECT 522.800 362.200 523.600 365.000 ;
        RECT 524.400 362.200 525.200 365.000 ;
        RECT 526.000 362.200 526.800 365.000 ;
        RECT 527.600 362.200 528.400 368.400 ;
        RECT 530.800 367.600 533.400 368.400 ;
        RECT 534.000 368.200 534.600 369.000 ;
        RECT 535.600 369.400 536.400 369.600 ;
        RECT 535.600 369.000 541.000 369.400 ;
        RECT 535.600 368.800 541.800 369.000 ;
        RECT 540.400 368.200 541.800 368.800 ;
        RECT 534.000 367.600 539.800 368.200 ;
        RECT 542.800 368.000 544.400 368.800 ;
        RECT 542.800 367.600 543.400 368.000 ;
        RECT 530.800 362.200 531.600 367.000 ;
        RECT 534.000 362.200 534.800 367.000 ;
        RECT 539.200 366.800 543.400 367.600 ;
        RECT 545.200 367.400 546.000 373.000 ;
        RECT 544.000 366.800 546.000 367.400 ;
        RECT 535.600 362.200 536.400 365.000 ;
        RECT 537.200 362.200 538.000 365.000 ;
        RECT 540.400 362.200 541.200 366.800 ;
        RECT 544.000 366.200 544.600 366.800 ;
        RECT 543.600 365.600 544.600 366.200 ;
        RECT 543.600 362.200 544.400 365.600 ;
        RECT 546.800 362.200 547.600 379.800 ;
        RECT 548.400 375.600 549.200 377.200 ;
        RECT 2.800 352.000 3.600 359.800 ;
        RECT 6.000 355.200 6.800 359.800 ;
        RECT 2.600 351.200 3.600 352.000 ;
        RECT 4.200 354.600 6.800 355.200 ;
        RECT 4.200 353.000 4.800 354.600 ;
        RECT 9.200 354.400 10.000 359.800 ;
        RECT 12.400 357.000 13.200 359.800 ;
        RECT 14.000 357.000 14.800 359.800 ;
        RECT 15.600 357.000 16.400 359.800 ;
        RECT 10.600 354.400 14.800 355.200 ;
        RECT 7.400 353.600 10.000 354.400 ;
        RECT 17.200 353.600 18.000 359.800 ;
        RECT 20.400 355.000 21.200 359.800 ;
        RECT 23.600 355.000 24.400 359.800 ;
        RECT 25.200 357.000 26.000 359.800 ;
        RECT 26.800 357.000 27.600 359.800 ;
        RECT 30.000 355.200 30.800 359.800 ;
        RECT 33.200 356.400 34.000 359.800 ;
        RECT 33.200 355.800 34.200 356.400 ;
        RECT 33.600 355.200 34.200 355.800 ;
        RECT 28.800 354.400 33.000 355.200 ;
        RECT 33.600 354.600 35.600 355.200 ;
        RECT 20.400 353.600 23.000 354.400 ;
        RECT 23.600 353.800 29.400 354.400 ;
        RECT 32.400 354.000 33.000 354.400 ;
        RECT 12.400 353.000 13.200 353.200 ;
        RECT 4.200 352.400 13.200 353.000 ;
        RECT 15.600 353.000 16.400 353.200 ;
        RECT 23.600 353.000 24.200 353.800 ;
        RECT 30.000 353.200 31.400 353.800 ;
        RECT 32.400 353.200 34.000 354.000 ;
        RECT 15.600 352.400 24.200 353.000 ;
        RECT 25.200 353.000 31.400 353.200 ;
        RECT 25.200 352.600 30.600 353.000 ;
        RECT 25.200 352.400 26.000 352.600 ;
        RECT 2.600 346.800 3.400 351.200 ;
        RECT 4.200 350.600 4.800 352.400 ;
        RECT 4.000 350.000 4.800 350.600 ;
        RECT 10.800 350.000 34.200 350.600 ;
        RECT 4.000 348.000 4.600 350.000 ;
        RECT 10.800 349.400 11.600 350.000 ;
        RECT 28.400 349.600 29.200 350.000 ;
        RECT 31.600 349.600 32.400 350.000 ;
        RECT 33.400 349.800 34.200 350.000 ;
        RECT 5.200 348.600 9.000 349.400 ;
        RECT 4.000 347.400 5.200 348.000 ;
        RECT 2.600 346.000 3.600 346.800 ;
        RECT 2.800 342.200 3.600 346.000 ;
        RECT 4.400 342.200 5.200 347.400 ;
        RECT 8.200 347.400 9.000 348.600 ;
        RECT 8.200 346.800 10.000 347.400 ;
        RECT 9.200 346.200 10.000 346.800 ;
        RECT 14.000 346.400 14.800 349.200 ;
        RECT 17.200 348.600 20.400 349.400 ;
        RECT 24.200 348.600 26.200 349.400 ;
        RECT 34.800 349.000 35.600 354.600 ;
        RECT 16.800 347.800 17.600 348.000 ;
        RECT 16.800 347.200 21.200 347.800 ;
        RECT 20.400 347.000 21.200 347.200 ;
        RECT 22.000 346.800 22.800 348.400 ;
        RECT 9.200 345.400 11.600 346.200 ;
        RECT 14.000 345.600 15.000 346.400 ;
        RECT 18.000 345.600 19.600 346.400 ;
        RECT 20.400 346.200 21.200 346.400 ;
        RECT 24.200 346.200 25.000 348.600 ;
        RECT 26.800 348.200 35.600 349.000 ;
        RECT 30.200 346.800 33.200 347.600 ;
        RECT 30.200 346.200 31.000 346.800 ;
        RECT 20.400 345.600 25.000 346.200 ;
        RECT 10.800 342.200 11.600 345.400 ;
        RECT 28.400 345.400 31.000 346.200 ;
        RECT 12.400 342.200 13.200 345.000 ;
        RECT 14.000 342.200 14.800 345.000 ;
        RECT 15.600 342.200 16.400 345.000 ;
        RECT 17.200 342.200 18.000 345.000 ;
        RECT 20.400 342.200 21.200 345.000 ;
        RECT 23.600 342.200 24.400 345.000 ;
        RECT 25.200 342.200 26.000 345.000 ;
        RECT 26.800 342.200 27.600 345.000 ;
        RECT 28.400 342.200 29.200 345.400 ;
        RECT 34.800 342.200 35.600 348.200 ;
        RECT 36.400 350.300 37.200 359.800 ;
        RECT 40.200 352.600 41.000 359.800 ;
        RECT 45.000 352.600 45.800 359.800 ;
        RECT 51.800 352.600 52.600 359.800 ;
        RECT 40.200 351.800 42.000 352.600 ;
        RECT 45.000 351.800 46.800 352.600 ;
        RECT 50.800 351.800 52.600 352.600 ;
        RECT 39.600 350.300 40.400 351.200 ;
        RECT 36.400 349.700 40.400 350.300 ;
        RECT 36.400 342.200 37.200 349.700 ;
        RECT 39.600 349.600 40.400 349.700 ;
        RECT 41.200 348.400 41.800 351.800 ;
        RECT 44.400 349.600 45.200 351.200 ;
        RECT 46.000 348.400 46.600 351.800 ;
        RECT 51.000 348.400 51.600 351.800 ;
        RECT 52.400 350.300 53.200 351.200 ;
        RECT 55.600 350.300 56.400 359.800 ;
        RECT 60.400 356.400 61.200 359.800 ;
        RECT 60.200 355.800 61.200 356.400 ;
        RECT 60.200 355.200 60.800 355.800 ;
        RECT 63.600 355.200 64.400 359.800 ;
        RECT 66.800 357.000 67.600 359.800 ;
        RECT 68.400 357.000 69.200 359.800 ;
        RECT 58.800 354.600 60.800 355.200 ;
        RECT 57.200 351.600 58.000 353.200 ;
        RECT 52.400 349.700 56.400 350.300 ;
        RECT 52.400 349.600 53.200 349.700 ;
        RECT 41.200 347.600 42.000 348.400 ;
        RECT 46.000 347.600 46.800 348.400 ;
        RECT 50.800 347.600 51.600 348.400 ;
        RECT 38.000 344.800 38.800 346.400 ;
        RECT 41.200 344.400 41.800 347.600 ;
        RECT 42.800 344.800 43.600 346.400 ;
        RECT 46.000 344.400 46.600 347.600 ;
        RECT 47.600 344.800 48.400 346.400 ;
        RECT 49.200 344.800 50.000 346.400 ;
        RECT 51.000 346.300 51.600 347.600 ;
        RECT 54.000 346.800 54.800 348.400 ;
        RECT 52.400 346.300 53.200 346.400 ;
        RECT 50.900 345.700 53.200 346.300 ;
        RECT 41.200 342.200 42.000 344.400 ;
        RECT 46.000 342.200 46.800 344.400 ;
        RECT 51.000 344.200 51.600 345.700 ;
        RECT 52.400 345.600 53.200 345.700 ;
        RECT 55.600 346.200 56.400 349.700 ;
        RECT 58.800 349.000 59.600 354.600 ;
        RECT 61.400 354.400 65.600 355.200 ;
        RECT 70.000 355.000 70.800 359.800 ;
        RECT 73.200 355.000 74.000 359.800 ;
        RECT 61.400 354.000 62.000 354.400 ;
        RECT 60.400 353.200 62.000 354.000 ;
        RECT 65.000 353.800 70.800 354.400 ;
        RECT 63.000 353.200 64.400 353.800 ;
        RECT 63.000 353.000 69.200 353.200 ;
        RECT 63.800 352.600 69.200 353.000 ;
        RECT 68.400 352.400 69.200 352.600 ;
        RECT 70.200 353.000 70.800 353.800 ;
        RECT 71.400 353.600 74.000 354.400 ;
        RECT 76.400 353.600 77.200 359.800 ;
        RECT 78.000 357.000 78.800 359.800 ;
        RECT 79.600 357.000 80.400 359.800 ;
        RECT 81.200 357.000 82.000 359.800 ;
        RECT 79.600 354.400 83.800 355.200 ;
        RECT 84.400 354.400 85.200 359.800 ;
        RECT 87.600 355.200 88.400 359.800 ;
        RECT 87.600 354.600 90.200 355.200 ;
        RECT 84.400 353.600 87.000 354.400 ;
        RECT 78.000 353.000 78.800 353.200 ;
        RECT 70.200 352.400 78.800 353.000 ;
        RECT 81.200 353.000 82.000 353.200 ;
        RECT 89.600 353.000 90.200 354.600 ;
        RECT 81.200 352.400 90.200 353.000 ;
        RECT 89.600 350.600 90.200 352.400 ;
        RECT 90.800 352.000 91.600 359.800 ;
        RECT 94.600 352.600 95.400 359.800 ;
        RECT 100.400 356.400 101.200 359.800 ;
        RECT 100.200 355.800 101.200 356.400 ;
        RECT 100.200 355.200 100.800 355.800 ;
        RECT 103.600 355.200 104.400 359.800 ;
        RECT 106.800 357.000 107.600 359.800 ;
        RECT 108.400 357.000 109.200 359.800 ;
        RECT 98.800 354.600 100.800 355.200 ;
        RECT 90.800 351.200 91.800 352.000 ;
        RECT 94.600 351.800 96.400 352.600 ;
        RECT 60.200 350.000 83.600 350.600 ;
        RECT 89.600 350.000 90.400 350.600 ;
        RECT 60.200 349.800 61.200 350.000 ;
        RECT 60.400 349.600 61.200 349.800 ;
        RECT 65.200 349.600 66.000 350.000 ;
        RECT 82.800 349.400 83.600 350.000 ;
        RECT 58.800 348.200 67.600 349.000 ;
        RECT 68.200 348.600 70.200 349.400 ;
        RECT 74.000 348.600 77.200 349.400 ;
        RECT 55.600 345.600 57.400 346.200 ;
        RECT 50.800 342.200 51.600 344.200 ;
        RECT 56.600 342.200 57.400 345.600 ;
        RECT 58.800 342.200 59.600 348.200 ;
        RECT 61.200 346.800 64.200 347.600 ;
        RECT 63.400 346.200 64.200 346.800 ;
        RECT 69.400 346.200 70.200 348.600 ;
        RECT 71.600 346.800 72.400 348.400 ;
        RECT 76.800 347.800 77.600 348.000 ;
        RECT 73.200 347.200 77.600 347.800 ;
        RECT 73.200 347.000 74.000 347.200 ;
        RECT 79.600 346.400 80.400 349.200 ;
        RECT 85.400 348.600 89.200 349.400 ;
        RECT 85.400 347.400 86.200 348.600 ;
        RECT 89.800 348.000 90.400 350.000 ;
        RECT 73.200 346.200 74.000 346.400 ;
        RECT 63.400 345.400 66.000 346.200 ;
        RECT 69.400 345.600 74.000 346.200 ;
        RECT 74.800 345.600 76.400 346.400 ;
        RECT 79.400 345.600 80.400 346.400 ;
        RECT 84.400 346.800 86.200 347.400 ;
        RECT 89.200 347.400 90.400 348.000 ;
        RECT 84.400 346.200 85.200 346.800 ;
        RECT 65.200 342.200 66.000 345.400 ;
        RECT 82.800 345.400 85.200 346.200 ;
        RECT 66.800 342.200 67.600 345.000 ;
        RECT 68.400 342.200 69.200 345.000 ;
        RECT 70.000 342.200 70.800 345.000 ;
        RECT 73.200 342.200 74.000 345.000 ;
        RECT 76.400 342.200 77.200 345.000 ;
        RECT 78.000 342.200 78.800 345.000 ;
        RECT 79.600 342.200 80.400 345.000 ;
        RECT 81.200 342.200 82.000 345.000 ;
        RECT 82.800 342.200 83.600 345.400 ;
        RECT 89.200 342.200 90.000 347.400 ;
        RECT 91.000 346.800 91.800 351.200 ;
        RECT 92.400 350.300 93.200 350.400 ;
        RECT 94.000 350.300 94.800 351.200 ;
        RECT 92.400 349.700 94.800 350.300 ;
        RECT 92.400 349.600 93.200 349.700 ;
        RECT 94.000 349.600 94.800 349.700 ;
        RECT 90.800 346.300 91.800 346.800 ;
        RECT 95.600 348.400 96.200 351.800 ;
        RECT 98.800 349.000 99.600 354.600 ;
        RECT 101.400 354.400 105.600 355.200 ;
        RECT 110.000 355.000 110.800 359.800 ;
        RECT 113.200 355.000 114.000 359.800 ;
        RECT 101.400 354.000 102.000 354.400 ;
        RECT 100.400 353.200 102.000 354.000 ;
        RECT 105.000 353.800 110.800 354.400 ;
        RECT 103.000 353.200 104.400 353.800 ;
        RECT 103.000 353.000 109.200 353.200 ;
        RECT 103.800 352.600 109.200 353.000 ;
        RECT 108.400 352.400 109.200 352.600 ;
        RECT 110.200 353.000 110.800 353.800 ;
        RECT 111.400 353.600 114.000 354.400 ;
        RECT 116.400 353.600 117.200 359.800 ;
        RECT 118.000 357.000 118.800 359.800 ;
        RECT 119.600 357.000 120.400 359.800 ;
        RECT 121.200 357.000 122.000 359.800 ;
        RECT 119.600 354.400 123.800 355.200 ;
        RECT 124.400 354.400 125.200 359.800 ;
        RECT 127.600 355.200 128.400 359.800 ;
        RECT 127.600 354.600 130.200 355.200 ;
        RECT 124.400 353.600 127.000 354.400 ;
        RECT 118.000 353.000 118.800 353.200 ;
        RECT 110.200 352.400 118.800 353.000 ;
        RECT 121.200 353.000 122.000 353.200 ;
        RECT 129.600 353.000 130.200 354.600 ;
        RECT 121.200 352.400 130.200 353.000 ;
        RECT 129.600 350.600 130.200 352.400 ;
        RECT 130.800 352.000 131.600 359.800 ;
        RECT 142.000 356.400 142.800 359.800 ;
        RECT 141.800 355.800 142.800 356.400 ;
        RECT 141.800 355.200 142.400 355.800 ;
        RECT 145.200 355.200 146.000 359.800 ;
        RECT 148.400 357.000 149.200 359.800 ;
        RECT 150.000 357.000 150.800 359.800 ;
        RECT 140.400 354.600 142.400 355.200 ;
        RECT 130.800 351.200 131.800 352.000 ;
        RECT 100.200 350.000 123.600 350.600 ;
        RECT 129.600 350.000 130.400 350.600 ;
        RECT 100.200 349.800 101.200 350.000 ;
        RECT 100.400 349.600 101.200 349.800 ;
        RECT 105.200 349.600 106.000 350.000 ;
        RECT 122.800 349.400 123.600 350.000 ;
        RECT 95.600 347.600 96.400 348.400 ;
        RECT 98.800 348.200 107.600 349.000 ;
        RECT 108.200 348.600 110.200 349.400 ;
        RECT 114.000 348.600 117.200 349.400 ;
        RECT 94.000 346.300 94.800 346.400 ;
        RECT 90.800 345.700 94.800 346.300 ;
        RECT 90.800 342.200 91.600 345.700 ;
        RECT 94.000 345.600 94.800 345.700 ;
        RECT 95.600 344.400 96.200 347.600 ;
        RECT 97.200 344.800 98.000 346.400 ;
        RECT 95.600 342.200 96.400 344.400 ;
        RECT 98.800 342.200 99.600 348.200 ;
        RECT 101.200 346.800 104.200 347.600 ;
        RECT 103.400 346.200 104.200 346.800 ;
        RECT 109.400 346.200 110.200 348.600 ;
        RECT 111.600 346.800 112.400 348.400 ;
        RECT 116.800 347.800 117.600 348.000 ;
        RECT 113.200 347.200 117.600 347.800 ;
        RECT 113.200 347.000 114.000 347.200 ;
        RECT 119.600 346.400 120.400 349.200 ;
        RECT 125.400 348.600 129.200 349.400 ;
        RECT 125.400 347.400 126.200 348.600 ;
        RECT 129.800 348.000 130.400 350.000 ;
        RECT 113.200 346.200 114.000 346.400 ;
        RECT 103.400 345.400 106.000 346.200 ;
        RECT 109.400 345.600 114.000 346.200 ;
        RECT 114.800 345.600 116.400 346.400 ;
        RECT 119.400 345.600 120.400 346.400 ;
        RECT 124.400 346.800 126.200 347.400 ;
        RECT 129.200 347.400 130.400 348.000 ;
        RECT 124.400 346.200 125.200 346.800 ;
        RECT 105.200 342.200 106.000 345.400 ;
        RECT 122.800 345.400 125.200 346.200 ;
        RECT 106.800 342.200 107.600 345.000 ;
        RECT 108.400 342.200 109.200 345.000 ;
        RECT 110.000 342.200 110.800 345.000 ;
        RECT 113.200 342.200 114.000 345.000 ;
        RECT 116.400 342.200 117.200 345.000 ;
        RECT 118.000 342.200 118.800 345.000 ;
        RECT 119.600 342.200 120.400 345.000 ;
        RECT 121.200 342.200 122.000 345.000 ;
        RECT 122.800 342.200 123.600 345.400 ;
        RECT 129.200 342.200 130.000 347.400 ;
        RECT 131.000 346.800 131.800 351.200 ;
        RECT 130.800 346.000 131.800 346.800 ;
        RECT 140.400 349.000 141.200 354.600 ;
        RECT 143.000 354.400 147.200 355.200 ;
        RECT 151.600 355.000 152.400 359.800 ;
        RECT 154.800 355.000 155.600 359.800 ;
        RECT 143.000 354.000 143.600 354.400 ;
        RECT 142.000 353.200 143.600 354.000 ;
        RECT 146.600 353.800 152.400 354.400 ;
        RECT 144.600 353.200 146.000 353.800 ;
        RECT 144.600 353.000 150.800 353.200 ;
        RECT 145.400 352.600 150.800 353.000 ;
        RECT 150.000 352.400 150.800 352.600 ;
        RECT 151.800 353.000 152.400 353.800 ;
        RECT 153.000 353.600 155.600 354.400 ;
        RECT 158.000 353.600 158.800 359.800 ;
        RECT 159.600 357.000 160.400 359.800 ;
        RECT 161.200 357.000 162.000 359.800 ;
        RECT 162.800 357.000 163.600 359.800 ;
        RECT 161.200 354.400 165.400 355.200 ;
        RECT 166.000 354.400 166.800 359.800 ;
        RECT 169.200 355.200 170.000 359.800 ;
        RECT 169.200 354.600 171.800 355.200 ;
        RECT 166.000 353.600 168.600 354.400 ;
        RECT 159.600 353.000 160.400 353.200 ;
        RECT 151.800 352.400 160.400 353.000 ;
        RECT 162.800 353.000 163.600 353.200 ;
        RECT 171.200 353.000 171.800 354.600 ;
        RECT 162.800 352.400 171.800 353.000 ;
        RECT 171.200 350.600 171.800 352.400 ;
        RECT 172.400 352.000 173.200 359.800 ;
        RECT 177.200 352.000 178.000 359.800 ;
        RECT 180.400 355.200 181.200 359.800 ;
        RECT 172.400 351.200 173.400 352.000 ;
        RECT 141.800 350.000 165.200 350.600 ;
        RECT 171.200 350.000 172.000 350.600 ;
        RECT 141.800 349.800 142.600 350.000 ;
        RECT 143.600 349.600 144.400 350.000 ;
        RECT 146.800 349.600 147.600 350.000 ;
        RECT 153.200 349.600 154.000 350.000 ;
        RECT 164.400 349.400 165.200 350.000 ;
        RECT 140.400 348.200 149.200 349.000 ;
        RECT 149.800 348.600 151.800 349.400 ;
        RECT 155.600 348.600 158.800 349.400 ;
        RECT 130.800 342.200 131.600 346.000 ;
        RECT 140.400 342.200 141.200 348.200 ;
        RECT 142.800 346.800 145.800 347.600 ;
        RECT 145.000 346.200 145.800 346.800 ;
        RECT 151.000 346.200 151.800 348.600 ;
        RECT 153.200 346.800 154.000 348.400 ;
        RECT 158.400 347.800 159.200 348.000 ;
        RECT 154.800 347.200 159.200 347.800 ;
        RECT 154.800 347.000 155.600 347.200 ;
        RECT 161.200 346.400 162.000 349.200 ;
        RECT 167.000 348.600 170.800 349.400 ;
        RECT 167.000 347.400 167.800 348.600 ;
        RECT 171.400 348.000 172.000 350.000 ;
        RECT 154.800 346.200 155.600 346.400 ;
        RECT 145.000 345.400 147.600 346.200 ;
        RECT 151.000 345.600 155.600 346.200 ;
        RECT 156.400 345.600 158.000 346.400 ;
        RECT 161.000 345.600 162.000 346.400 ;
        RECT 166.000 346.800 167.800 347.400 ;
        RECT 170.800 347.400 172.000 348.000 ;
        RECT 166.000 346.200 166.800 346.800 ;
        RECT 146.800 342.200 147.600 345.400 ;
        RECT 164.400 345.400 166.800 346.200 ;
        RECT 148.400 342.200 149.200 345.000 ;
        RECT 150.000 342.200 150.800 345.000 ;
        RECT 151.600 342.200 152.400 345.000 ;
        RECT 154.800 342.200 155.600 345.000 ;
        RECT 158.000 342.200 158.800 345.000 ;
        RECT 159.600 342.200 160.400 345.000 ;
        RECT 161.200 342.200 162.000 345.000 ;
        RECT 162.800 342.200 163.600 345.000 ;
        RECT 164.400 342.200 165.200 345.400 ;
        RECT 170.800 342.200 171.600 347.400 ;
        RECT 172.600 346.800 173.400 351.200 ;
        RECT 172.400 346.000 173.400 346.800 ;
        RECT 177.000 351.200 178.000 352.000 ;
        RECT 178.600 354.600 181.200 355.200 ;
        RECT 178.600 353.000 179.200 354.600 ;
        RECT 183.600 354.400 184.400 359.800 ;
        RECT 186.800 357.000 187.600 359.800 ;
        RECT 188.400 357.000 189.200 359.800 ;
        RECT 190.000 357.000 190.800 359.800 ;
        RECT 185.000 354.400 189.200 355.200 ;
        RECT 181.800 353.600 184.400 354.400 ;
        RECT 191.600 353.600 192.400 359.800 ;
        RECT 194.800 355.000 195.600 359.800 ;
        RECT 198.000 355.000 198.800 359.800 ;
        RECT 199.600 357.000 200.400 359.800 ;
        RECT 201.200 357.000 202.000 359.800 ;
        RECT 204.400 355.200 205.200 359.800 ;
        RECT 207.600 356.400 208.400 359.800 ;
        RECT 207.600 355.800 208.600 356.400 ;
        RECT 208.000 355.200 208.600 355.800 ;
        RECT 203.200 354.400 207.400 355.200 ;
        RECT 208.000 354.600 210.000 355.200 ;
        RECT 194.800 353.600 197.400 354.400 ;
        RECT 198.000 353.800 203.800 354.400 ;
        RECT 206.800 354.000 207.400 354.400 ;
        RECT 186.800 353.000 187.600 353.200 ;
        RECT 178.600 352.400 187.600 353.000 ;
        RECT 190.000 353.000 190.800 353.200 ;
        RECT 198.000 353.000 198.600 353.800 ;
        RECT 204.400 353.200 205.800 353.800 ;
        RECT 206.800 353.200 208.400 354.000 ;
        RECT 190.000 352.400 198.600 353.000 ;
        RECT 199.600 353.000 205.800 353.200 ;
        RECT 199.600 352.600 205.000 353.000 ;
        RECT 199.600 352.400 200.400 352.600 ;
        RECT 177.000 346.800 177.800 351.200 ;
        RECT 178.600 350.600 179.200 352.400 ;
        RECT 178.400 350.000 179.200 350.600 ;
        RECT 185.200 350.000 208.600 350.600 ;
        RECT 178.400 348.000 179.000 350.000 ;
        RECT 185.200 349.400 186.000 350.000 ;
        RECT 202.800 349.600 203.600 350.000 ;
        RECT 206.000 349.600 206.800 350.000 ;
        RECT 207.800 349.800 208.600 350.000 ;
        RECT 179.600 348.600 183.400 349.400 ;
        RECT 178.400 347.400 179.600 348.000 ;
        RECT 177.000 346.000 178.000 346.800 ;
        RECT 172.400 342.200 173.200 346.000 ;
        RECT 177.200 342.200 178.000 346.000 ;
        RECT 178.800 342.200 179.600 347.400 ;
        RECT 182.600 347.400 183.400 348.600 ;
        RECT 182.600 346.800 184.400 347.400 ;
        RECT 183.600 346.200 184.400 346.800 ;
        RECT 188.400 346.400 189.200 349.200 ;
        RECT 191.600 348.600 194.800 349.400 ;
        RECT 198.600 348.600 200.600 349.400 ;
        RECT 209.200 349.000 210.000 354.600 ;
        RECT 212.400 352.000 213.200 359.800 ;
        RECT 215.600 355.200 216.400 359.800 ;
        RECT 191.200 347.800 192.000 348.000 ;
        RECT 191.200 347.200 195.600 347.800 ;
        RECT 194.800 347.000 195.600 347.200 ;
        RECT 196.400 346.800 197.200 348.400 ;
        RECT 183.600 345.400 186.000 346.200 ;
        RECT 188.400 345.600 189.400 346.400 ;
        RECT 192.400 345.600 194.000 346.400 ;
        RECT 194.800 346.200 195.600 346.400 ;
        RECT 198.600 346.200 199.400 348.600 ;
        RECT 201.200 348.200 210.000 349.000 ;
        RECT 204.600 346.800 207.600 347.600 ;
        RECT 204.600 346.200 205.400 346.800 ;
        RECT 194.800 345.600 199.400 346.200 ;
        RECT 185.200 342.200 186.000 345.400 ;
        RECT 202.800 345.400 205.400 346.200 ;
        RECT 186.800 342.200 187.600 345.000 ;
        RECT 188.400 342.200 189.200 345.000 ;
        RECT 190.000 342.200 190.800 345.000 ;
        RECT 191.600 342.200 192.400 345.000 ;
        RECT 194.800 342.200 195.600 345.000 ;
        RECT 198.000 342.200 198.800 345.000 ;
        RECT 199.600 342.200 200.400 345.000 ;
        RECT 201.200 342.200 202.000 345.000 ;
        RECT 202.800 342.200 203.600 345.400 ;
        RECT 209.200 342.200 210.000 348.200 ;
        RECT 212.200 351.200 213.200 352.000 ;
        RECT 213.800 354.600 216.400 355.200 ;
        RECT 213.800 353.000 214.400 354.600 ;
        RECT 218.800 354.400 219.600 359.800 ;
        RECT 222.000 357.000 222.800 359.800 ;
        RECT 223.600 357.000 224.400 359.800 ;
        RECT 225.200 357.000 226.000 359.800 ;
        RECT 220.200 354.400 224.400 355.200 ;
        RECT 217.000 353.600 219.600 354.400 ;
        RECT 226.800 353.600 227.600 359.800 ;
        RECT 230.000 355.000 230.800 359.800 ;
        RECT 233.200 355.000 234.000 359.800 ;
        RECT 234.800 357.000 235.600 359.800 ;
        RECT 236.400 357.000 237.200 359.800 ;
        RECT 239.600 355.200 240.400 359.800 ;
        RECT 242.800 356.400 243.600 359.800 ;
        RECT 242.800 355.800 243.800 356.400 ;
        RECT 246.000 355.800 246.800 359.800 ;
        RECT 243.200 355.200 243.800 355.800 ;
        RECT 246.200 355.600 246.800 355.800 ;
        RECT 249.200 355.800 250.000 359.800 ;
        RECT 252.400 355.800 253.200 359.800 ;
        RECT 249.200 355.600 249.800 355.800 ;
        RECT 238.400 354.400 242.600 355.200 ;
        RECT 243.200 354.600 245.200 355.200 ;
        RECT 230.000 353.600 232.600 354.400 ;
        RECT 233.200 353.800 239.000 354.400 ;
        RECT 242.000 354.000 242.600 354.400 ;
        RECT 222.000 353.000 222.800 353.200 ;
        RECT 213.800 352.400 222.800 353.000 ;
        RECT 225.200 353.000 226.000 353.200 ;
        RECT 233.200 353.000 233.800 353.800 ;
        RECT 239.600 353.200 241.000 353.800 ;
        RECT 242.000 353.200 243.600 354.000 ;
        RECT 225.200 352.400 233.800 353.000 ;
        RECT 234.800 353.000 241.000 353.200 ;
        RECT 234.800 352.600 240.200 353.000 ;
        RECT 234.800 352.400 235.600 352.600 ;
        RECT 212.200 346.800 213.000 351.200 ;
        RECT 213.800 350.600 214.400 352.400 ;
        RECT 213.600 350.000 214.400 350.600 ;
        RECT 220.400 350.000 243.800 350.600 ;
        RECT 213.600 348.000 214.200 350.000 ;
        RECT 220.400 349.400 221.200 350.000 ;
        RECT 238.000 349.600 238.800 350.000 ;
        RECT 242.800 349.800 243.800 350.000 ;
        RECT 242.800 349.600 243.600 349.800 ;
        RECT 214.800 348.600 218.600 349.400 ;
        RECT 213.600 347.400 214.800 348.000 ;
        RECT 212.200 346.000 213.200 346.800 ;
        RECT 212.400 342.200 213.200 346.000 ;
        RECT 214.000 342.200 214.800 347.400 ;
        RECT 217.800 347.400 218.600 348.600 ;
        RECT 217.800 346.800 219.600 347.400 ;
        RECT 218.800 346.200 219.600 346.800 ;
        RECT 223.600 346.400 224.400 349.200 ;
        RECT 226.800 348.600 230.000 349.400 ;
        RECT 233.800 348.600 235.800 349.400 ;
        RECT 244.400 349.000 245.200 354.600 ;
        RECT 246.200 355.000 249.800 355.600 ;
        RECT 252.600 355.600 253.200 355.800 ;
        RECT 255.600 355.800 256.400 359.800 ;
        RECT 266.800 356.400 267.600 359.800 ;
        RECT 266.600 355.800 267.600 356.400 ;
        RECT 255.600 355.600 256.200 355.800 ;
        RECT 252.600 355.000 256.200 355.600 ;
        RECT 266.600 355.200 267.200 355.800 ;
        RECT 270.000 355.200 270.800 359.800 ;
        RECT 273.200 357.000 274.000 359.800 ;
        RECT 274.800 357.000 275.600 359.800 ;
        RECT 246.200 352.400 246.800 355.000 ;
        RECT 247.600 352.800 248.400 354.400 ;
        RECT 252.600 352.400 253.200 355.000 ;
        RECT 265.200 354.600 267.200 355.200 ;
        RECT 254.000 352.800 254.800 354.400 ;
        RECT 246.000 351.600 246.800 352.400 ;
        RECT 226.400 347.800 227.200 348.000 ;
        RECT 226.400 347.200 230.800 347.800 ;
        RECT 230.000 347.000 230.800 347.200 ;
        RECT 231.600 346.800 232.400 348.400 ;
        RECT 218.800 345.400 221.200 346.200 ;
        RECT 223.600 345.600 224.600 346.400 ;
        RECT 227.600 345.600 229.200 346.400 ;
        RECT 230.000 346.200 230.800 346.400 ;
        RECT 233.800 346.200 234.600 348.600 ;
        RECT 236.400 348.200 245.200 349.000 ;
        RECT 239.800 346.800 242.800 347.600 ;
        RECT 239.800 346.200 240.600 346.800 ;
        RECT 230.000 345.600 234.600 346.200 ;
        RECT 220.400 342.200 221.200 345.400 ;
        RECT 238.000 345.400 240.600 346.200 ;
        RECT 222.000 342.200 222.800 345.000 ;
        RECT 223.600 342.200 224.400 345.000 ;
        RECT 225.200 342.200 226.000 345.000 ;
        RECT 226.800 342.200 227.600 345.000 ;
        RECT 230.000 342.200 230.800 345.000 ;
        RECT 233.200 342.200 234.000 345.000 ;
        RECT 234.800 342.200 235.600 345.000 ;
        RECT 236.400 342.200 237.200 345.000 ;
        RECT 238.000 342.200 238.800 345.400 ;
        RECT 244.400 342.200 245.200 348.200 ;
        RECT 246.200 348.400 246.800 351.600 ;
        RECT 250.800 350.800 251.600 352.400 ;
        RECT 252.400 351.600 253.200 352.400 ;
        RECT 248.400 349.600 250.000 350.400 ;
        RECT 252.600 348.400 253.200 351.600 ;
        RECT 257.200 350.800 258.000 352.400 ;
        RECT 254.800 349.600 256.400 350.400 ;
        RECT 265.200 349.000 266.000 354.600 ;
        RECT 267.800 354.400 272.000 355.200 ;
        RECT 276.400 355.000 277.200 359.800 ;
        RECT 279.600 355.000 280.400 359.800 ;
        RECT 267.800 354.000 268.400 354.400 ;
        RECT 266.800 353.200 268.400 354.000 ;
        RECT 271.400 353.800 277.200 354.400 ;
        RECT 269.400 353.200 270.800 353.800 ;
        RECT 269.400 353.000 275.600 353.200 ;
        RECT 270.200 352.600 275.600 353.000 ;
        RECT 274.800 352.400 275.600 352.600 ;
        RECT 276.600 353.000 277.200 353.800 ;
        RECT 277.800 353.600 280.400 354.400 ;
        RECT 282.800 353.600 283.600 359.800 ;
        RECT 284.400 357.000 285.200 359.800 ;
        RECT 286.000 357.000 286.800 359.800 ;
        RECT 287.600 357.000 288.400 359.800 ;
        RECT 286.000 354.400 290.200 355.200 ;
        RECT 290.800 354.400 291.600 359.800 ;
        RECT 294.000 355.200 294.800 359.800 ;
        RECT 294.000 354.600 296.600 355.200 ;
        RECT 290.800 353.600 293.400 354.400 ;
        RECT 284.400 353.000 285.200 353.200 ;
        RECT 276.600 352.400 285.200 353.000 ;
        RECT 287.600 353.000 288.400 353.200 ;
        RECT 296.000 353.000 296.600 354.600 ;
        RECT 287.600 352.400 296.600 353.000 ;
        RECT 296.000 350.600 296.600 352.400 ;
        RECT 297.200 352.000 298.000 359.800 ;
        RECT 300.400 355.800 301.200 359.800 ;
        RECT 300.600 355.600 301.200 355.800 ;
        RECT 303.600 355.800 304.400 359.800 ;
        RECT 303.600 355.600 304.200 355.800 ;
        RECT 300.600 355.000 304.200 355.600 ;
        RECT 300.600 352.400 301.200 355.000 ;
        RECT 302.000 352.800 302.800 354.400 ;
        RECT 307.400 352.600 308.200 359.800 ;
        RECT 297.200 351.200 298.200 352.000 ;
        RECT 300.400 351.600 301.200 352.400 ;
        RECT 266.600 350.000 290.000 350.600 ;
        RECT 296.000 350.000 296.800 350.600 ;
        RECT 266.600 349.800 267.400 350.000 ;
        RECT 268.400 349.600 269.200 350.000 ;
        RECT 270.000 349.600 270.800 350.000 ;
        RECT 271.600 349.600 272.400 350.000 ;
        RECT 289.200 349.400 290.000 350.000 ;
        RECT 246.200 348.200 247.800 348.400 ;
        RECT 252.600 348.200 254.200 348.400 ;
        RECT 265.200 348.200 274.000 349.000 ;
        RECT 274.600 348.600 276.600 349.400 ;
        RECT 280.400 348.600 283.600 349.400 ;
        RECT 246.200 347.800 248.000 348.200 ;
        RECT 252.600 347.800 254.400 348.200 ;
        RECT 247.200 342.200 248.000 347.800 ;
        RECT 253.600 342.200 254.400 347.800 ;
        RECT 265.200 342.200 266.000 348.200 ;
        RECT 267.600 346.800 270.600 347.600 ;
        RECT 269.800 346.200 270.600 346.800 ;
        RECT 275.800 346.200 276.600 348.600 ;
        RECT 278.000 346.800 278.800 348.400 ;
        RECT 283.200 347.800 284.000 348.000 ;
        RECT 279.600 347.200 284.000 347.800 ;
        RECT 279.600 347.000 280.400 347.200 ;
        RECT 286.000 346.400 286.800 349.200 ;
        RECT 291.800 348.600 295.600 349.400 ;
        RECT 291.800 347.400 292.600 348.600 ;
        RECT 296.200 348.000 296.800 350.000 ;
        RECT 279.600 346.200 280.400 346.400 ;
        RECT 269.800 345.400 272.400 346.200 ;
        RECT 275.800 345.600 280.400 346.200 ;
        RECT 281.200 345.600 282.800 346.400 ;
        RECT 285.800 345.600 286.800 346.400 ;
        RECT 290.800 346.800 292.600 347.400 ;
        RECT 295.600 347.400 296.800 348.000 ;
        RECT 290.800 346.200 291.600 346.800 ;
        RECT 271.600 342.200 272.400 345.400 ;
        RECT 289.200 345.400 291.600 346.200 ;
        RECT 273.200 342.200 274.000 345.000 ;
        RECT 274.800 342.200 275.600 345.000 ;
        RECT 276.400 342.200 277.200 345.000 ;
        RECT 279.600 342.200 280.400 345.000 ;
        RECT 282.800 342.200 283.600 345.000 ;
        RECT 284.400 342.200 285.200 345.000 ;
        RECT 286.000 342.200 286.800 345.000 ;
        RECT 287.600 342.200 288.400 345.000 ;
        RECT 289.200 342.200 290.000 345.400 ;
        RECT 295.600 342.200 296.400 347.400 ;
        RECT 297.400 346.800 298.200 351.200 ;
        RECT 300.600 348.400 301.200 351.600 ;
        RECT 305.200 350.800 306.000 352.400 ;
        RECT 307.400 351.800 309.200 352.600 ;
        RECT 311.600 351.800 312.400 359.800 ;
        RECT 314.800 355.800 315.600 359.800 ;
        RECT 302.800 349.600 304.400 350.400 ;
        RECT 306.800 349.600 307.600 351.200 ;
        RECT 308.400 350.300 309.000 351.800 ;
        RECT 311.600 350.400 312.200 351.800 ;
        RECT 314.800 351.600 315.400 355.800 ;
        RECT 313.000 351.000 315.400 351.600 ;
        RECT 310.000 350.300 310.800 350.400 ;
        RECT 308.400 349.700 310.800 350.300 ;
        RECT 308.400 348.400 309.000 349.700 ;
        RECT 310.000 349.600 310.800 349.700 ;
        RECT 311.600 349.600 312.400 350.400 ;
        RECT 300.600 348.200 302.200 348.400 ;
        RECT 300.600 347.800 302.400 348.200 ;
        RECT 297.200 346.000 298.200 346.800 ;
        RECT 297.200 342.200 298.000 346.000 ;
        RECT 301.600 342.200 302.400 347.800 ;
        RECT 308.400 347.600 309.200 348.400 ;
        RECT 308.400 344.200 309.000 347.600 ;
        RECT 310.000 344.800 310.800 346.400 ;
        RECT 311.600 346.200 312.200 349.600 ;
        RECT 313.000 347.600 313.600 351.000 ;
        RECT 314.800 349.600 315.600 350.400 ;
        RECT 314.800 348.800 315.400 349.600 ;
        RECT 314.400 348.200 315.400 348.800 ;
        RECT 316.400 348.300 317.200 349.200 ;
        RECT 318.000 348.300 318.800 348.400 ;
        RECT 314.400 348.000 315.200 348.200 ;
        RECT 316.400 347.700 318.800 348.300 ;
        RECT 316.400 347.600 317.200 347.700 ;
        RECT 312.800 347.400 313.600 347.600 ;
        RECT 312.800 347.000 315.800 347.400 ;
        RECT 312.800 346.800 317.000 347.000 ;
        RECT 318.000 346.800 318.800 347.700 ;
        RECT 315.200 346.400 317.000 346.800 ;
        RECT 316.400 346.200 317.000 346.400 ;
        RECT 319.600 346.200 320.400 359.800 ;
        RECT 322.800 355.800 323.600 359.800 ;
        RECT 323.000 355.600 323.600 355.800 ;
        RECT 326.000 355.800 326.800 359.800 ;
        RECT 326.000 355.600 326.600 355.800 ;
        RECT 323.000 355.000 326.600 355.600 ;
        RECT 321.200 351.600 322.000 353.200 ;
        RECT 323.000 352.400 323.600 355.000 ;
        RECT 324.400 352.800 325.200 354.400 ;
        RECT 322.800 351.600 323.600 352.400 ;
        RECT 323.000 348.400 323.600 351.600 ;
        RECT 327.600 350.800 328.400 352.400 ;
        RECT 329.200 351.800 330.000 359.800 ;
        RECT 330.800 352.400 331.600 359.800 ;
        RECT 334.000 352.400 334.800 359.800 ;
        RECT 335.600 355.800 336.400 359.800 ;
        RECT 335.800 355.600 336.400 355.800 ;
        RECT 338.800 355.800 339.600 359.800 ;
        RECT 338.800 355.600 339.400 355.800 ;
        RECT 335.800 355.000 339.400 355.600 ;
        RECT 335.800 352.400 336.400 355.000 ;
        RECT 337.200 352.800 338.000 354.400 ;
        RECT 338.800 354.300 339.600 354.400 ;
        RECT 342.600 354.300 343.400 359.800 ;
        RECT 338.800 353.700 343.400 354.300 ;
        RECT 338.800 353.600 339.600 353.700 ;
        RECT 342.600 352.600 343.400 353.700 ;
        RECT 347.400 352.600 348.200 359.800 ;
        RECT 330.800 351.800 334.800 352.400 ;
        RECT 329.400 350.400 330.000 351.800 ;
        RECT 335.600 351.600 336.400 352.400 ;
        RECT 333.200 350.400 334.000 350.800 ;
        RECT 325.200 349.600 326.800 350.400 ;
        RECT 329.200 349.800 331.600 350.400 ;
        RECT 333.200 349.800 334.800 350.400 ;
        RECT 329.200 349.600 330.000 349.800 ;
        RECT 330.800 349.600 331.600 349.800 ;
        RECT 334.000 349.600 334.800 349.800 ;
        RECT 323.000 348.200 324.600 348.400 ;
        RECT 323.000 347.800 324.800 348.200 ;
        RECT 311.600 345.200 313.000 346.200 ;
        RECT 308.400 342.200 309.200 344.200 ;
        RECT 312.200 342.200 313.000 345.200 ;
        RECT 316.400 342.200 317.200 346.200 ;
        RECT 319.600 345.600 321.400 346.200 ;
        RECT 320.600 342.200 321.400 345.600 ;
        RECT 324.000 342.200 324.800 347.800 ;
        RECT 329.200 345.600 330.000 346.400 ;
        RECT 331.000 346.200 331.600 349.600 ;
        RECT 332.400 347.600 333.200 349.200 ;
        RECT 335.800 348.400 336.400 351.600 ;
        RECT 340.400 350.800 341.200 352.400 ;
        RECT 342.600 351.800 344.400 352.600 ;
        RECT 347.400 351.800 349.200 352.600 ;
        RECT 354.200 352.400 355.000 359.800 ;
        RECT 360.200 358.400 361.000 359.800 ;
        RECT 367.000 358.400 369.000 359.800 ;
        RECT 360.200 357.600 362.000 358.400 ;
        RECT 367.000 357.600 370.000 358.400 ;
        RECT 355.600 353.600 356.400 354.400 ;
        RECT 355.800 352.400 356.400 353.600 ;
        RECT 358.800 353.600 359.600 354.400 ;
        RECT 358.800 352.400 359.400 353.600 ;
        RECT 360.200 352.400 361.000 357.600 ;
        RECT 354.200 351.800 355.200 352.400 ;
        RECT 355.800 351.800 357.200 352.400 ;
        RECT 338.000 349.600 339.600 350.400 ;
        RECT 342.000 349.600 342.800 351.200 ;
        RECT 343.600 348.400 344.200 351.800 ;
        RECT 346.800 349.600 347.600 351.200 ;
        RECT 348.400 348.400 349.000 351.800 ;
        RECT 353.200 348.800 354.000 350.400 ;
        RECT 354.600 350.300 355.200 351.800 ;
        RECT 356.400 351.600 357.200 351.800 ;
        RECT 358.000 351.800 359.400 352.400 ;
        RECT 360.000 351.800 361.000 352.400 ;
        RECT 367.000 351.800 369.000 357.600 ;
        RECT 374.600 354.400 375.400 359.800 ;
        RECT 373.200 353.600 374.000 354.400 ;
        RECT 374.600 353.600 376.400 354.400 ;
        RECT 373.200 352.400 373.800 353.600 ;
        RECT 374.600 352.400 375.400 353.600 ;
        RECT 372.400 351.800 373.800 352.400 ;
        RECT 374.400 351.800 375.400 352.400 ;
        RECT 378.800 351.800 379.600 359.800 ;
        RECT 380.400 352.400 381.200 359.800 ;
        RECT 383.600 352.400 384.400 359.800 ;
        RECT 380.400 351.800 384.400 352.400 ;
        RECT 358.000 351.600 358.800 351.800 ;
        RECT 358.100 350.300 358.700 351.600 ;
        RECT 354.600 349.700 358.700 350.300 ;
        RECT 354.600 348.400 355.200 349.700 ;
        RECT 360.000 348.400 360.600 351.800 ;
        RECT 361.200 348.800 362.000 350.400 ;
        RECT 366.000 348.800 366.800 350.400 ;
        RECT 367.600 348.400 368.200 351.800 ;
        RECT 372.400 351.600 373.200 351.800 ;
        RECT 369.200 348.800 370.000 350.400 ;
        RECT 335.800 347.800 338.000 348.400 ;
        RECT 336.800 347.600 338.000 347.800 ;
        RECT 343.600 347.600 344.400 348.400 ;
        RECT 345.200 348.300 346.000 348.400 ;
        RECT 348.400 348.300 349.200 348.400 ;
        RECT 351.600 348.300 352.400 348.400 ;
        RECT 345.200 347.700 349.200 348.300 ;
        RECT 345.200 347.600 346.000 347.700 ;
        RECT 348.400 347.600 349.200 347.700 ;
        RECT 350.100 348.200 352.400 348.300 ;
        RECT 350.100 347.700 353.200 348.200 ;
        RECT 329.400 344.800 330.200 345.600 ;
        RECT 330.800 342.200 331.600 346.200 ;
        RECT 336.800 342.200 337.600 347.600 ;
        RECT 343.600 344.200 344.200 347.600 ;
        RECT 345.200 344.800 346.000 346.400 ;
        RECT 348.400 344.200 349.000 347.600 ;
        RECT 350.100 346.400 350.700 347.700 ;
        RECT 351.600 347.600 353.200 347.700 ;
        RECT 354.600 347.600 357.200 348.400 ;
        RECT 358.000 347.600 360.600 348.400 ;
        RECT 362.800 348.200 363.600 348.400 ;
        RECT 362.000 347.600 363.600 348.200 ;
        RECT 364.400 348.200 365.200 348.400 ;
        RECT 367.600 348.200 368.400 348.400 ;
        RECT 364.400 347.600 366.000 348.200 ;
        RECT 367.600 347.600 370.000 348.200 ;
        RECT 370.800 347.600 371.600 349.200 ;
        RECT 374.400 348.400 375.000 351.800 ;
        RECT 379.000 350.400 379.600 351.800 ;
        RECT 382.800 350.400 383.600 350.800 ;
        RECT 375.600 348.800 376.400 350.400 ;
        RECT 378.800 349.800 381.200 350.400 ;
        RECT 382.800 349.800 384.400 350.400 ;
        RECT 378.800 349.600 379.600 349.800 ;
        RECT 372.400 347.600 375.000 348.400 ;
        RECT 377.200 348.200 378.000 348.400 ;
        RECT 376.400 347.600 378.000 348.200 ;
        RECT 352.400 347.200 353.200 347.600 ;
        RECT 350.000 344.800 350.800 346.400 ;
        RECT 351.800 346.200 355.400 346.600 ;
        RECT 356.400 346.200 357.000 347.600 ;
        RECT 358.200 346.200 358.800 347.600 ;
        RECT 362.000 347.200 362.800 347.600 ;
        RECT 365.200 347.200 366.000 347.600 ;
        RECT 359.800 346.200 363.400 346.600 ;
        RECT 364.600 346.200 368.200 346.600 ;
        RECT 369.400 346.200 370.000 347.600 ;
        RECT 372.600 346.200 373.200 347.600 ;
        RECT 376.400 347.200 377.200 347.600 ;
        RECT 374.200 346.200 377.800 346.600 ;
        RECT 351.600 346.000 355.600 346.200 ;
        RECT 343.600 342.200 344.400 344.200 ;
        RECT 348.400 342.200 349.200 344.200 ;
        RECT 351.600 342.200 352.400 346.000 ;
        RECT 354.800 342.200 355.600 346.000 ;
        RECT 356.400 342.200 357.200 346.200 ;
        RECT 358.000 342.200 358.800 346.200 ;
        RECT 359.600 346.000 363.600 346.200 ;
        RECT 359.600 342.200 360.400 346.000 ;
        RECT 362.800 342.200 363.600 346.000 ;
        RECT 364.400 346.000 368.400 346.200 ;
        RECT 364.400 342.200 365.200 346.000 ;
        RECT 367.600 342.800 368.400 346.000 ;
        RECT 369.200 343.400 370.000 346.200 ;
        RECT 370.800 342.800 371.600 346.200 ;
        RECT 367.600 342.200 371.600 342.800 ;
        RECT 372.400 342.200 373.200 346.200 ;
        RECT 374.000 346.000 378.000 346.200 ;
        RECT 374.000 342.200 374.800 346.000 ;
        RECT 377.200 342.200 378.000 346.000 ;
        RECT 378.800 345.600 379.600 346.400 ;
        RECT 380.600 346.200 381.200 349.800 ;
        RECT 383.600 349.600 384.400 349.800 ;
        RECT 382.000 347.600 382.800 349.200 ;
        RECT 379.000 344.800 379.800 345.600 ;
        RECT 380.400 342.200 381.200 346.200 ;
        RECT 385.200 342.200 386.000 359.800 ;
        RECT 388.400 351.800 389.200 359.800 ;
        RECT 390.000 352.400 390.800 359.800 ;
        RECT 393.200 352.400 394.000 359.800 ;
        RECT 390.000 351.800 394.000 352.400 ;
        RECT 394.800 352.400 395.600 359.800 ;
        RECT 398.000 352.400 398.800 359.800 ;
        RECT 394.800 351.800 398.800 352.400 ;
        RECT 399.600 351.800 400.400 359.800 ;
        RECT 401.200 352.400 402.000 359.800 ;
        RECT 404.400 352.400 405.200 359.800 ;
        RECT 401.200 351.800 405.200 352.400 ;
        RECT 406.000 351.800 406.800 359.800 ;
        RECT 407.600 353.800 408.400 359.800 ;
        RECT 407.800 353.200 408.400 353.800 ;
        RECT 410.800 359.200 414.800 359.800 ;
        RECT 410.800 353.800 411.600 359.200 ;
        RECT 412.400 353.800 413.200 358.600 ;
        RECT 414.000 354.000 414.800 359.200 ;
        RECT 415.800 359.200 419.400 359.800 ;
        RECT 415.800 359.000 416.400 359.200 ;
        RECT 410.800 353.200 411.400 353.800 ;
        RECT 407.800 352.600 411.400 353.200 ;
        RECT 412.600 353.400 413.200 353.800 ;
        RECT 415.600 353.400 416.400 359.000 ;
        RECT 418.800 359.000 419.400 359.200 ;
        RECT 412.600 353.000 416.400 353.400 ;
        RECT 417.200 353.000 418.000 358.600 ;
        RECT 418.800 353.000 419.600 359.000 ;
        RECT 421.000 354.400 421.800 359.800 ;
        RECT 420.400 353.600 421.800 354.400 ;
        RECT 412.600 352.800 416.200 353.000 ;
        RECT 417.200 352.400 417.800 353.000 ;
        RECT 421.000 352.600 421.800 353.600 ;
        RECT 417.200 352.200 418.000 352.400 ;
        RECT 388.600 350.400 389.200 351.800 ;
        RECT 392.400 350.400 393.200 350.800 ;
        RECT 395.600 350.400 396.400 350.800 ;
        RECT 399.600 350.400 400.200 351.800 ;
        RECT 402.000 350.400 402.800 350.800 ;
        RECT 406.000 350.400 406.600 351.800 ;
        RECT 414.600 351.600 418.000 352.200 ;
        RECT 421.000 351.800 422.800 352.600 ;
        RECT 388.400 349.800 390.800 350.400 ;
        RECT 392.400 349.800 394.000 350.400 ;
        RECT 388.400 349.600 389.200 349.800 ;
        RECT 386.800 346.800 387.600 348.400 ;
        RECT 388.400 345.600 389.200 346.400 ;
        RECT 390.200 346.200 390.800 349.800 ;
        RECT 393.200 349.600 394.000 349.800 ;
        RECT 394.800 349.800 396.400 350.400 ;
        RECT 398.000 349.800 400.400 350.400 ;
        RECT 394.800 349.600 395.600 349.800 ;
        RECT 398.000 349.600 398.800 349.800 ;
        RECT 399.600 349.600 400.400 349.800 ;
        RECT 401.200 349.800 402.800 350.400 ;
        RECT 404.400 349.800 406.800 350.400 ;
        RECT 401.200 349.600 402.000 349.800 ;
        RECT 391.600 347.600 392.400 349.200 ;
        RECT 396.400 347.600 397.200 349.200 ;
        RECT 388.600 344.800 389.400 345.600 ;
        RECT 390.000 342.200 390.800 346.200 ;
        RECT 398.000 346.200 398.600 349.600 ;
        RECT 402.800 347.600 403.600 349.200 ;
        RECT 398.000 342.200 398.800 346.200 ;
        RECT 399.600 345.600 400.400 346.400 ;
        RECT 404.400 346.200 405.000 349.800 ;
        RECT 406.000 349.600 406.800 349.800 ;
        RECT 412.400 349.600 414.000 350.400 ;
        RECT 410.800 347.600 412.400 348.400 ;
        RECT 406.000 346.300 406.800 346.400 ;
        RECT 407.600 346.300 408.400 346.400 ;
        RECT 399.400 344.800 400.200 345.600 ;
        RECT 404.400 342.200 405.200 346.200 ;
        RECT 406.000 345.700 408.400 346.300 ;
        RECT 406.000 345.600 406.800 345.700 ;
        RECT 407.600 345.600 408.400 345.700 ;
        RECT 409.200 345.600 411.000 346.400 ;
        RECT 405.800 344.800 406.600 345.600 ;
        RECT 414.600 345.000 415.200 351.600 ;
        RECT 420.400 349.600 421.200 351.200 ;
        RECT 411.200 344.400 415.200 345.000 ;
        RECT 410.800 343.600 411.800 344.400 ;
        RECT 414.000 344.200 415.200 344.400 ;
        RECT 422.000 348.400 422.600 351.800 ;
        RECT 433.200 350.300 434.000 359.800 ;
        RECT 434.800 351.600 435.600 353.200 ;
        RECT 436.400 350.300 437.200 350.400 ;
        RECT 433.200 349.700 437.200 350.300 ;
        RECT 422.000 348.300 422.800 348.400 ;
        RECT 431.600 348.300 432.400 348.400 ;
        RECT 422.000 347.700 432.400 348.300 ;
        RECT 422.000 347.600 422.800 347.700 ;
        RECT 422.000 344.200 422.600 347.600 ;
        RECT 431.600 346.800 432.400 347.700 ;
        RECT 423.600 344.800 424.400 346.400 ;
        RECT 433.200 346.200 434.000 349.700 ;
        RECT 436.400 349.600 437.200 349.700 ;
        RECT 436.400 346.800 437.200 348.400 ;
        RECT 438.000 346.200 438.800 359.800 ;
        RECT 442.800 355.800 443.600 359.800 ;
        RECT 443.000 355.600 443.600 355.800 ;
        RECT 446.000 355.800 446.800 359.800 ;
        RECT 446.000 355.600 446.600 355.800 ;
        RECT 443.000 355.000 446.600 355.600 ;
        RECT 439.600 351.600 440.400 353.200 ;
        RECT 444.400 352.800 445.200 354.400 ;
        RECT 446.000 352.400 446.600 355.000 ;
        RECT 450.200 354.400 451.000 359.800 ;
        RECT 449.200 353.600 451.000 354.400 ;
        RECT 451.600 353.600 452.400 354.400 ;
        RECT 450.200 352.400 451.000 353.600 ;
        RECT 451.800 352.400 452.400 353.600 ;
        RECT 441.200 350.800 442.000 352.400 ;
        RECT 446.000 351.600 446.800 352.400 ;
        RECT 450.200 351.800 451.200 352.400 ;
        RECT 451.800 351.800 453.200 352.400 ;
        RECT 456.600 351.800 458.600 359.800 ;
        RECT 462.800 353.600 463.600 354.400 ;
        RECT 462.800 352.400 463.400 353.600 ;
        RECT 464.200 352.400 465.000 359.800 ;
        RECT 462.000 351.800 463.400 352.400 ;
        RECT 442.800 349.600 444.400 350.400 ;
        RECT 446.000 348.400 446.600 351.600 ;
        RECT 449.200 348.800 450.000 350.400 ;
        RECT 450.600 348.400 451.200 351.800 ;
        RECT 452.400 351.600 453.200 351.800 ;
        RECT 455.600 348.800 456.400 350.400 ;
        RECT 457.200 348.400 457.800 351.800 ;
        RECT 462.000 351.600 462.800 351.800 ;
        RECT 464.000 351.600 466.000 352.400 ;
        RECT 458.800 348.800 459.600 350.400 ;
        RECT 462.000 350.300 462.800 350.400 ;
        RECT 464.000 350.300 464.600 351.600 ;
        RECT 462.000 349.700 464.600 350.300 ;
        RECT 462.000 349.600 462.800 349.700 ;
        RECT 445.000 348.200 446.600 348.400 ;
        RECT 444.800 347.800 446.600 348.200 ;
        RECT 447.600 348.200 448.400 348.400 ;
        RECT 433.200 345.600 435.000 346.200 ;
        RECT 438.000 345.600 439.800 346.200 ;
        RECT 410.800 342.200 411.600 343.600 ;
        RECT 414.000 342.200 414.800 344.200 ;
        RECT 422.000 342.200 422.800 344.200 ;
        RECT 434.200 342.200 435.000 345.600 ;
        RECT 439.000 344.400 439.800 345.600 ;
        RECT 439.000 343.600 440.400 344.400 ;
        RECT 439.000 342.200 439.800 343.600 ;
        RECT 444.800 342.200 445.600 347.800 ;
        RECT 447.600 347.600 449.200 348.200 ;
        RECT 450.600 347.600 453.200 348.400 ;
        RECT 454.000 348.200 454.800 348.400 ;
        RECT 457.200 348.200 458.000 348.400 ;
        RECT 454.000 347.600 455.600 348.200 ;
        RECT 457.200 347.600 459.600 348.200 ;
        RECT 460.400 347.600 461.200 349.200 ;
        RECT 464.000 348.400 464.600 349.700 ;
        RECT 465.200 348.800 466.000 350.400 ;
        RECT 462.000 347.600 464.600 348.400 ;
        RECT 466.800 348.200 467.600 348.400 ;
        RECT 466.000 347.600 467.600 348.200 ;
        RECT 448.400 347.200 449.200 347.600 ;
        RECT 447.800 346.200 451.400 346.600 ;
        RECT 452.400 346.200 453.000 347.600 ;
        RECT 454.800 347.200 455.600 347.600 ;
        RECT 454.200 346.200 457.800 346.600 ;
        RECT 459.000 346.200 459.600 347.600 ;
        RECT 462.200 346.200 462.800 347.600 ;
        RECT 466.000 347.200 466.800 347.600 ;
        RECT 463.800 346.200 467.400 346.600 ;
        RECT 447.600 346.000 451.600 346.200 ;
        RECT 447.600 342.200 448.400 346.000 ;
        RECT 450.800 342.200 451.600 346.000 ;
        RECT 452.400 342.200 453.200 346.200 ;
        RECT 454.000 346.000 458.000 346.200 ;
        RECT 454.000 342.200 454.800 346.000 ;
        RECT 457.200 342.800 458.000 346.000 ;
        RECT 458.800 343.400 459.600 346.200 ;
        RECT 460.400 342.800 461.200 346.200 ;
        RECT 457.200 342.200 461.200 342.800 ;
        RECT 462.000 342.200 462.800 346.200 ;
        RECT 463.600 346.000 467.600 346.200 ;
        RECT 463.600 342.200 464.400 346.000 ;
        RECT 466.800 342.200 467.600 346.000 ;
        RECT 468.400 342.200 469.200 359.800 ;
        RECT 474.200 356.400 475.000 359.800 ;
        RECT 480.600 358.400 481.400 359.800 ;
        RECT 479.600 357.600 481.400 358.400 ;
        RECT 473.200 355.600 475.000 356.400 ;
        RECT 474.200 352.400 475.000 355.600 ;
        RECT 475.600 353.600 476.400 354.400 ;
        RECT 475.800 352.400 476.400 353.600 ;
        RECT 480.600 352.400 481.400 357.600 ;
        RECT 482.000 353.600 482.800 354.400 ;
        RECT 482.200 352.400 482.800 353.600 ;
        RECT 474.200 351.800 475.200 352.400 ;
        RECT 475.800 351.800 477.200 352.400 ;
        RECT 480.600 351.800 481.600 352.400 ;
        RECT 482.200 351.800 483.600 352.400 ;
        RECT 473.200 348.800 474.000 350.400 ;
        RECT 474.600 348.400 475.200 351.800 ;
        RECT 476.400 351.600 477.200 351.800 ;
        RECT 479.600 348.800 480.400 350.400 ;
        RECT 481.000 348.400 481.600 351.800 ;
        RECT 482.800 351.600 483.600 351.800 ;
        RECT 471.600 348.200 472.400 348.400 ;
        RECT 471.600 347.600 473.200 348.200 ;
        RECT 474.600 347.600 477.200 348.400 ;
        RECT 478.000 348.200 478.800 348.400 ;
        RECT 478.000 347.600 479.600 348.200 ;
        RECT 481.000 347.600 483.600 348.400 ;
        RECT 472.400 347.200 473.200 347.600 ;
        RECT 470.000 344.800 470.800 346.400 ;
        RECT 471.800 346.200 475.400 346.600 ;
        RECT 476.400 346.200 477.000 347.600 ;
        RECT 478.800 347.200 479.600 347.600 ;
        RECT 478.200 346.200 481.800 346.600 ;
        RECT 482.800 346.200 483.400 347.600 ;
        RECT 471.600 346.000 475.600 346.200 ;
        RECT 471.600 342.200 472.400 346.000 ;
        RECT 474.800 342.200 475.600 346.000 ;
        RECT 476.400 342.200 477.200 346.200 ;
        RECT 478.000 346.000 482.000 346.200 ;
        RECT 478.000 342.200 478.800 346.000 ;
        RECT 481.200 342.200 482.000 346.000 ;
        RECT 482.800 342.200 483.600 346.200 ;
        RECT 484.400 344.800 485.200 346.400 ;
        RECT 486.000 342.200 486.800 359.800 ;
        RECT 489.200 352.300 490.000 359.800 ;
        RECT 492.400 355.600 493.200 359.800 ;
        RECT 495.600 355.800 496.400 359.800 ;
        RECT 495.600 355.600 496.200 355.800 ;
        RECT 498.800 355.600 499.600 359.800 ;
        RECT 502.000 355.800 502.800 359.800 ;
        RECT 504.200 358.400 505.000 359.800 ;
        RECT 504.200 357.600 506.000 358.400 ;
        RECT 502.000 355.600 502.600 355.800 ;
        RECT 492.600 355.000 496.200 355.600 ;
        RECT 499.000 355.000 502.600 355.600 ;
        RECT 494.000 352.800 494.800 354.400 ;
        RECT 495.600 352.400 496.200 355.000 ;
        RECT 500.400 352.800 501.200 354.400 ;
        RECT 502.000 352.400 502.600 355.000 ;
        RECT 504.200 352.600 505.000 357.600 ;
        RECT 490.800 352.300 491.600 352.400 ;
        RECT 489.200 351.700 491.600 352.300 ;
        RECT 487.600 344.800 488.400 346.400 ;
        RECT 489.200 342.200 490.000 351.700 ;
        RECT 490.800 350.800 491.600 351.700 ;
        RECT 495.600 351.600 496.400 352.400 ;
        RECT 492.400 349.600 494.000 350.400 ;
        RECT 495.600 348.400 496.200 351.600 ;
        RECT 497.200 350.800 498.000 352.400 ;
        RECT 502.000 351.600 502.800 352.400 ;
        RECT 504.200 351.800 506.000 352.600 ;
        RECT 508.400 351.800 509.200 359.800 ;
        RECT 510.000 352.400 510.800 359.800 ;
        RECT 513.200 352.400 514.000 359.800 ;
        RECT 510.000 351.800 514.000 352.400 ;
        RECT 516.400 352.000 517.200 359.800 ;
        RECT 519.600 355.200 520.400 359.800 ;
        RECT 498.800 349.600 500.400 350.400 ;
        RECT 502.000 348.400 502.600 351.600 ;
        RECT 503.600 349.600 504.400 351.200 ;
        RECT 494.600 348.200 496.200 348.400 ;
        RECT 501.000 348.200 502.600 348.400 ;
        RECT 494.400 347.800 496.200 348.200 ;
        RECT 500.800 347.800 502.600 348.200 ;
        RECT 505.200 348.400 505.800 351.800 ;
        RECT 508.600 350.400 509.200 351.800 ;
        RECT 516.200 351.200 517.200 352.000 ;
        RECT 517.800 354.600 520.400 355.200 ;
        RECT 517.800 353.000 518.400 354.600 ;
        RECT 522.800 354.400 523.600 359.800 ;
        RECT 526.000 357.000 526.800 359.800 ;
        RECT 527.600 357.000 528.400 359.800 ;
        RECT 529.200 357.000 530.000 359.800 ;
        RECT 524.200 354.400 528.400 355.200 ;
        RECT 521.000 353.600 523.600 354.400 ;
        RECT 530.800 353.600 531.600 359.800 ;
        RECT 534.000 355.000 534.800 359.800 ;
        RECT 537.200 355.000 538.000 359.800 ;
        RECT 538.800 357.000 539.600 359.800 ;
        RECT 540.400 357.000 541.200 359.800 ;
        RECT 543.600 355.200 544.400 359.800 ;
        RECT 546.800 356.400 547.600 359.800 ;
        RECT 546.800 355.800 547.800 356.400 ;
        RECT 547.200 355.200 547.800 355.800 ;
        RECT 542.400 354.400 546.600 355.200 ;
        RECT 547.200 354.600 549.200 355.200 ;
        RECT 534.000 353.600 536.600 354.400 ;
        RECT 537.200 353.800 543.000 354.400 ;
        RECT 546.000 354.000 546.600 354.400 ;
        RECT 526.000 353.000 526.800 353.200 ;
        RECT 517.800 352.400 526.800 353.000 ;
        RECT 529.200 353.000 530.000 353.200 ;
        RECT 537.200 353.000 537.800 353.800 ;
        RECT 543.600 353.200 545.000 353.800 ;
        RECT 546.000 353.200 547.600 354.000 ;
        RECT 529.200 352.400 537.800 353.000 ;
        RECT 538.800 353.000 545.000 353.200 ;
        RECT 538.800 352.600 544.200 353.000 ;
        RECT 538.800 352.400 539.600 352.600 ;
        RECT 512.400 350.400 513.200 350.800 ;
        RECT 508.400 349.800 510.800 350.400 ;
        RECT 512.400 349.800 514.000 350.400 ;
        RECT 508.400 349.600 509.200 349.800 ;
        RECT 494.400 342.200 495.200 347.800 ;
        RECT 500.800 342.200 501.600 347.800 ;
        RECT 505.200 347.600 506.000 348.400 ;
        RECT 505.200 344.200 505.800 347.600 ;
        RECT 506.800 344.800 507.600 346.400 ;
        RECT 508.400 345.600 509.200 346.400 ;
        RECT 510.200 346.200 510.800 349.800 ;
        RECT 513.200 349.600 514.000 349.800 ;
        RECT 511.600 347.600 512.400 349.200 ;
        RECT 508.600 344.800 509.400 345.600 ;
        RECT 505.200 342.200 506.000 344.200 ;
        RECT 510.000 342.200 510.800 346.200 ;
        RECT 516.200 346.800 517.000 351.200 ;
        RECT 517.800 350.600 518.400 352.400 ;
        RECT 517.600 350.000 518.400 350.600 ;
        RECT 524.400 350.000 547.800 350.600 ;
        RECT 517.600 348.000 518.200 350.000 ;
        RECT 524.400 349.400 525.200 350.000 ;
        RECT 542.000 349.600 542.800 350.000 ;
        RECT 547.000 349.800 547.800 350.000 ;
        RECT 518.800 348.600 522.600 349.400 ;
        RECT 517.600 347.400 518.800 348.000 ;
        RECT 516.200 346.000 517.200 346.800 ;
        RECT 516.400 342.200 517.200 346.000 ;
        RECT 518.000 342.200 518.800 347.400 ;
        RECT 521.800 347.400 522.600 348.600 ;
        RECT 521.800 346.800 523.600 347.400 ;
        RECT 522.800 346.200 523.600 346.800 ;
        RECT 527.600 346.400 528.400 349.200 ;
        RECT 530.800 348.600 534.000 349.400 ;
        RECT 537.800 348.600 539.800 349.400 ;
        RECT 548.400 349.000 549.200 354.600 ;
        RECT 530.400 347.800 531.200 348.000 ;
        RECT 530.400 347.200 534.800 347.800 ;
        RECT 534.000 347.000 534.800 347.200 ;
        RECT 535.600 346.800 536.400 348.400 ;
        RECT 522.800 345.400 525.200 346.200 ;
        RECT 527.600 345.600 528.600 346.400 ;
        RECT 531.600 345.600 533.200 346.400 ;
        RECT 534.000 346.200 534.800 346.400 ;
        RECT 537.800 346.200 538.600 348.600 ;
        RECT 540.400 348.200 549.200 349.000 ;
        RECT 543.800 346.800 546.800 347.600 ;
        RECT 543.800 346.200 544.600 346.800 ;
        RECT 534.000 345.600 538.600 346.200 ;
        RECT 524.400 342.200 525.200 345.400 ;
        RECT 542.000 345.400 544.600 346.200 ;
        RECT 526.000 342.200 526.800 345.000 ;
        RECT 527.600 342.200 528.400 345.000 ;
        RECT 529.200 342.200 530.000 345.000 ;
        RECT 530.800 342.200 531.600 345.000 ;
        RECT 534.000 342.200 534.800 345.000 ;
        RECT 537.200 342.200 538.000 345.000 ;
        RECT 538.800 342.200 539.600 345.000 ;
        RECT 540.400 342.200 541.200 345.000 ;
        RECT 542.000 342.200 542.800 345.400 ;
        RECT 548.400 342.200 549.200 348.200 ;
        RECT 1.200 335.600 2.000 337.200 ;
        RECT 2.800 322.200 3.600 339.800 ;
        RECT 6.000 336.000 6.800 339.800 ;
        RECT 5.800 335.200 6.800 336.000 ;
        RECT 5.800 330.800 6.600 335.200 ;
        RECT 7.600 334.600 8.400 339.800 ;
        RECT 14.000 336.600 14.800 339.800 ;
        RECT 15.600 337.000 16.400 339.800 ;
        RECT 17.200 337.000 18.000 339.800 ;
        RECT 18.800 337.000 19.600 339.800 ;
        RECT 20.400 337.000 21.200 339.800 ;
        RECT 23.600 337.000 24.400 339.800 ;
        RECT 26.800 337.000 27.600 339.800 ;
        RECT 28.400 337.000 29.200 339.800 ;
        RECT 30.000 337.000 30.800 339.800 ;
        RECT 12.400 335.800 14.800 336.600 ;
        RECT 31.600 336.600 32.400 339.800 ;
        RECT 12.400 335.200 13.200 335.800 ;
        RECT 7.200 334.000 8.400 334.600 ;
        RECT 11.400 334.600 13.200 335.200 ;
        RECT 17.200 335.600 18.200 336.400 ;
        RECT 21.200 335.600 22.800 336.400 ;
        RECT 23.600 335.800 28.200 336.400 ;
        RECT 31.600 335.800 34.200 336.600 ;
        RECT 23.600 335.600 24.400 335.800 ;
        RECT 7.200 332.000 7.800 334.000 ;
        RECT 11.400 333.400 12.200 334.600 ;
        RECT 8.400 332.600 12.200 333.400 ;
        RECT 17.200 332.800 18.000 335.600 ;
        RECT 23.600 334.800 24.400 335.000 ;
        RECT 20.000 334.200 24.400 334.800 ;
        RECT 20.000 334.000 20.800 334.200 ;
        RECT 25.200 333.600 26.000 335.200 ;
        RECT 27.400 333.400 28.200 335.800 ;
        RECT 33.400 335.200 34.200 335.800 ;
        RECT 33.400 334.400 36.400 335.200 ;
        RECT 38.000 333.800 38.800 339.800 ;
        RECT 42.200 336.400 43.000 339.800 ;
        RECT 41.200 335.800 43.000 336.400 ;
        RECT 44.400 335.800 45.200 339.800 ;
        RECT 46.000 336.000 46.800 339.800 ;
        RECT 49.200 336.000 50.000 339.800 ;
        RECT 46.000 335.800 50.000 336.000 ;
        RECT 20.400 332.600 23.600 333.400 ;
        RECT 27.400 332.600 29.400 333.400 ;
        RECT 30.000 333.000 38.800 333.800 ;
        RECT 39.600 333.600 40.400 335.200 ;
        RECT 14.000 332.000 14.800 332.600 ;
        RECT 31.600 332.000 32.400 332.400 ;
        RECT 36.600 332.000 37.400 332.200 ;
        RECT 7.200 331.400 8.000 332.000 ;
        RECT 14.000 331.400 37.400 332.000 ;
        RECT 5.800 330.000 6.800 330.800 ;
        RECT 4.400 328.300 5.200 328.400 ;
        RECT 6.000 328.300 6.800 330.000 ;
        RECT 4.400 327.700 6.800 328.300 ;
        RECT 4.400 327.600 5.200 327.700 ;
        RECT 6.000 322.200 6.800 327.700 ;
        RECT 7.400 329.600 8.000 331.400 ;
        RECT 7.400 329.000 16.400 329.600 ;
        RECT 7.400 327.400 8.000 329.000 ;
        RECT 15.600 328.800 16.400 329.000 ;
        RECT 18.800 329.000 27.400 329.600 ;
        RECT 18.800 328.800 19.600 329.000 ;
        RECT 10.600 327.600 13.200 328.400 ;
        RECT 7.400 326.800 10.000 327.400 ;
        RECT 9.200 322.200 10.000 326.800 ;
        RECT 12.400 322.200 13.200 327.600 ;
        RECT 13.800 326.800 18.000 327.600 ;
        RECT 15.600 322.200 16.400 325.000 ;
        RECT 17.200 322.200 18.000 325.000 ;
        RECT 18.800 322.200 19.600 325.000 ;
        RECT 20.400 322.200 21.200 328.400 ;
        RECT 23.600 327.600 26.200 328.400 ;
        RECT 26.800 328.200 27.400 329.000 ;
        RECT 28.400 329.400 29.200 329.600 ;
        RECT 28.400 329.000 33.800 329.400 ;
        RECT 28.400 328.800 34.600 329.000 ;
        RECT 33.200 328.200 34.600 328.800 ;
        RECT 26.800 327.600 32.600 328.200 ;
        RECT 35.600 328.000 37.200 328.800 ;
        RECT 35.600 327.600 36.200 328.000 ;
        RECT 23.600 322.200 24.400 327.000 ;
        RECT 26.800 322.200 27.600 327.000 ;
        RECT 32.000 326.800 36.200 327.600 ;
        RECT 38.000 327.400 38.800 333.000 ;
        RECT 36.800 326.800 38.800 327.400 ;
        RECT 41.200 332.300 42.000 335.800 ;
        RECT 44.600 334.400 45.200 335.800 ;
        RECT 46.200 335.400 49.800 335.800 ;
        RECT 48.400 334.400 49.200 334.800 ;
        RECT 44.400 333.600 47.000 334.400 ;
        RECT 48.400 333.800 50.000 334.400 ;
        RECT 54.400 334.200 55.200 339.800 ;
        RECT 60.800 334.200 61.600 339.800 ;
        RECT 63.600 335.800 64.400 339.800 ;
        RECT 65.200 336.000 66.000 339.800 ;
        RECT 68.400 336.000 69.200 339.800 ;
        RECT 65.200 335.800 69.200 336.000 ;
        RECT 70.600 336.400 71.400 339.800 ;
        RECT 75.400 336.400 76.200 339.800 ;
        RECT 81.200 337.800 82.000 339.800 ;
        RECT 70.600 335.800 72.400 336.400 ;
        RECT 63.800 334.400 64.400 335.800 ;
        RECT 65.400 335.400 69.000 335.800 ;
        RECT 67.600 334.400 68.400 334.800 ;
        RECT 54.400 333.800 56.200 334.200 ;
        RECT 60.800 333.800 62.600 334.200 ;
        RECT 49.200 333.600 50.000 333.800 ;
        RECT 54.600 333.600 56.200 333.800 ;
        RECT 61.000 333.600 62.600 333.800 ;
        RECT 63.600 333.600 66.200 334.400 ;
        RECT 67.600 334.300 69.200 334.400 ;
        RECT 71.600 334.300 72.400 335.800 ;
        RECT 74.800 335.600 77.200 336.400 ;
        RECT 79.600 335.600 80.400 337.200 ;
        RECT 67.600 333.800 72.400 334.300 ;
        RECT 68.400 333.700 72.400 333.800 ;
        RECT 68.400 333.600 69.200 333.700 ;
        RECT 41.200 331.700 45.100 332.300 ;
        RECT 28.400 322.200 29.200 325.000 ;
        RECT 30.000 322.200 30.800 325.000 ;
        RECT 33.200 322.200 34.000 326.800 ;
        RECT 36.800 326.200 37.400 326.800 ;
        RECT 36.400 325.600 37.400 326.200 ;
        RECT 36.400 322.200 37.200 325.600 ;
        RECT 41.200 322.200 42.000 331.700 ;
        RECT 44.500 330.400 45.100 331.700 ;
        RECT 42.800 328.800 43.600 330.400 ;
        RECT 44.400 330.200 45.200 330.400 ;
        RECT 46.400 330.200 47.000 333.600 ;
        RECT 47.600 331.600 48.400 333.200 ;
        RECT 52.400 331.600 54.000 332.400 ;
        RECT 44.400 329.600 45.800 330.200 ;
        RECT 46.400 329.600 47.400 330.200 ;
        RECT 50.800 329.600 51.600 331.200 ;
        RECT 55.600 330.400 56.200 333.600 ;
        RECT 58.800 331.600 60.400 332.400 ;
        RECT 62.000 332.300 62.600 333.600 ;
        RECT 63.600 332.300 64.400 332.400 ;
        RECT 62.000 331.700 64.400 332.300 ;
        RECT 55.600 329.600 56.400 330.400 ;
        RECT 57.200 329.600 58.000 331.200 ;
        RECT 62.000 330.400 62.600 331.700 ;
        RECT 63.600 331.600 64.400 331.700 ;
        RECT 62.000 329.600 62.800 330.400 ;
        RECT 63.600 330.200 64.400 330.400 ;
        RECT 65.600 330.200 66.200 333.600 ;
        RECT 66.800 331.600 67.600 333.200 ;
        RECT 63.600 329.600 65.000 330.200 ;
        RECT 65.600 329.600 66.600 330.200 ;
        RECT 45.200 328.400 45.800 329.600 ;
        RECT 45.200 327.600 46.000 328.400 ;
        RECT 46.600 322.200 47.400 329.600 ;
        RECT 54.000 327.600 54.800 329.200 ;
        RECT 55.600 327.000 56.200 329.600 ;
        RECT 60.400 327.600 61.200 329.200 ;
        RECT 62.000 327.000 62.600 329.600 ;
        RECT 64.400 328.400 65.000 329.600 ;
        RECT 64.400 327.600 65.200 328.400 ;
        RECT 52.600 326.400 56.200 327.000 ;
        RECT 52.400 322.200 53.200 326.400 ;
        RECT 55.600 326.200 56.200 326.400 ;
        RECT 59.000 326.400 62.600 327.000 ;
        RECT 59.000 326.200 59.600 326.400 ;
        RECT 55.600 322.200 56.400 326.200 ;
        RECT 58.800 322.200 59.600 326.200 ;
        RECT 62.000 326.200 62.600 326.400 ;
        RECT 62.000 322.200 62.800 326.200 ;
        RECT 65.800 322.200 66.600 329.600 ;
        RECT 70.000 328.800 70.800 330.400 ;
        RECT 71.600 322.200 72.400 333.700 ;
        RECT 73.200 333.600 74.000 335.200 ;
        RECT 74.800 328.800 75.600 330.400 ;
        RECT 76.400 322.200 77.200 335.600 ;
        RECT 78.000 334.300 78.800 335.200 ;
        RECT 81.400 334.400 82.000 337.800 ;
        RECT 81.200 334.300 82.000 334.400 ;
        RECT 78.000 333.700 82.000 334.300 ;
        RECT 85.600 334.200 86.400 339.800 ;
        RECT 78.000 333.600 78.800 333.700 ;
        RECT 81.200 333.600 82.000 333.700 ;
        RECT 81.400 330.200 82.000 333.600 ;
        RECT 84.600 333.800 86.400 334.200 ;
        RECT 84.600 333.600 86.200 333.800 ;
        RECT 82.800 330.800 83.600 332.400 ;
        RECT 84.600 330.400 85.200 333.600 ;
        RECT 86.800 331.600 88.400 332.400 ;
        RECT 81.200 329.400 83.000 330.200 ;
        RECT 84.400 329.600 85.200 330.400 ;
        RECT 89.200 329.600 90.000 331.200 ;
        RECT 82.200 322.200 83.000 329.400 ;
        RECT 84.600 327.000 85.200 329.600 ;
        RECT 86.000 327.600 86.800 329.200 ;
        RECT 84.600 326.400 88.200 327.000 ;
        RECT 84.600 326.200 85.200 326.400 ;
        RECT 84.400 322.200 85.200 326.200 ;
        RECT 87.600 326.200 88.200 326.400 ;
        RECT 87.600 322.200 88.400 326.200 ;
        RECT 90.800 322.200 91.600 339.800 ;
        RECT 92.400 335.600 93.200 337.200 ;
        RECT 95.600 336.000 96.400 339.800 ;
        RECT 95.400 335.200 96.400 336.000 ;
        RECT 95.400 330.800 96.200 335.200 ;
        RECT 97.200 334.600 98.000 339.800 ;
        RECT 103.600 336.600 104.400 339.800 ;
        RECT 105.200 337.000 106.000 339.800 ;
        RECT 106.800 337.000 107.600 339.800 ;
        RECT 108.400 337.000 109.200 339.800 ;
        RECT 110.000 337.000 110.800 339.800 ;
        RECT 113.200 337.000 114.000 339.800 ;
        RECT 116.400 337.000 117.200 339.800 ;
        RECT 118.000 337.000 118.800 339.800 ;
        RECT 119.600 337.000 120.400 339.800 ;
        RECT 102.000 335.800 104.400 336.600 ;
        RECT 121.200 336.600 122.000 339.800 ;
        RECT 102.000 335.200 102.800 335.800 ;
        RECT 96.800 334.000 98.000 334.600 ;
        RECT 101.000 334.600 102.800 335.200 ;
        RECT 106.800 335.600 107.800 336.400 ;
        RECT 110.800 335.600 112.400 336.400 ;
        RECT 113.200 335.800 117.800 336.400 ;
        RECT 121.200 335.800 123.800 336.600 ;
        RECT 113.200 335.600 114.000 335.800 ;
        RECT 96.800 332.000 97.400 334.000 ;
        RECT 101.000 333.400 101.800 334.600 ;
        RECT 98.000 332.600 101.800 333.400 ;
        RECT 106.800 332.800 107.600 335.600 ;
        RECT 113.200 334.800 114.000 335.000 ;
        RECT 109.600 334.200 114.000 334.800 ;
        RECT 109.600 334.000 110.400 334.200 ;
        RECT 114.800 333.600 115.600 335.200 ;
        RECT 117.000 333.400 117.800 335.800 ;
        RECT 123.000 335.200 123.800 335.800 ;
        RECT 123.000 334.400 126.000 335.200 ;
        RECT 127.600 333.800 128.400 339.800 ;
        RECT 110.000 332.600 113.200 333.400 ;
        RECT 117.000 332.600 119.000 333.400 ;
        RECT 119.600 333.000 128.400 333.800 ;
        RECT 103.600 332.000 104.400 332.600 ;
        RECT 121.200 332.000 122.000 332.400 ;
        RECT 122.800 332.000 123.600 332.400 ;
        RECT 126.200 332.000 127.000 332.200 ;
        RECT 96.800 331.400 97.600 332.000 ;
        RECT 103.600 331.400 127.000 332.000 ;
        RECT 95.400 330.000 96.400 330.800 ;
        RECT 95.600 322.200 96.400 330.000 ;
        RECT 97.000 329.600 97.600 331.400 ;
        RECT 97.000 329.000 106.000 329.600 ;
        RECT 97.000 327.400 97.600 329.000 ;
        RECT 105.200 328.800 106.000 329.000 ;
        RECT 108.400 329.000 117.000 329.600 ;
        RECT 108.400 328.800 109.200 329.000 ;
        RECT 100.200 327.600 102.800 328.400 ;
        RECT 97.000 326.800 99.600 327.400 ;
        RECT 98.800 322.200 99.600 326.800 ;
        RECT 102.000 322.200 102.800 327.600 ;
        RECT 103.400 326.800 107.600 327.600 ;
        RECT 105.200 322.200 106.000 325.000 ;
        RECT 106.800 322.200 107.600 325.000 ;
        RECT 108.400 322.200 109.200 325.000 ;
        RECT 110.000 322.200 110.800 328.400 ;
        RECT 113.200 327.600 115.800 328.400 ;
        RECT 116.400 328.200 117.000 329.000 ;
        RECT 118.000 329.400 118.800 329.600 ;
        RECT 118.000 329.000 123.400 329.400 ;
        RECT 118.000 328.800 124.200 329.000 ;
        RECT 122.800 328.200 124.200 328.800 ;
        RECT 116.400 327.600 122.200 328.200 ;
        RECT 125.200 328.000 126.800 328.800 ;
        RECT 125.200 327.600 125.800 328.000 ;
        RECT 113.200 322.200 114.000 327.000 ;
        RECT 116.400 322.200 117.200 327.000 ;
        RECT 121.600 326.800 125.800 327.600 ;
        RECT 127.600 327.400 128.400 333.000 ;
        RECT 126.400 326.800 128.400 327.400 ;
        RECT 135.600 333.800 136.400 339.800 ;
        RECT 142.000 336.600 142.800 339.800 ;
        RECT 143.600 337.000 144.400 339.800 ;
        RECT 145.200 337.000 146.000 339.800 ;
        RECT 146.800 337.000 147.600 339.800 ;
        RECT 150.000 337.000 150.800 339.800 ;
        RECT 153.200 337.000 154.000 339.800 ;
        RECT 154.800 337.000 155.600 339.800 ;
        RECT 156.400 337.000 157.200 339.800 ;
        RECT 158.000 337.000 158.800 339.800 ;
        RECT 140.200 335.800 142.800 336.600 ;
        RECT 159.600 336.600 160.400 339.800 ;
        RECT 146.200 335.800 150.800 336.400 ;
        RECT 140.200 335.200 141.000 335.800 ;
        RECT 138.000 334.400 141.000 335.200 ;
        RECT 135.600 333.000 144.400 333.800 ;
        RECT 146.200 333.400 147.000 335.800 ;
        RECT 150.000 335.600 150.800 335.800 ;
        RECT 151.600 335.600 153.200 336.400 ;
        RECT 156.200 335.600 157.200 336.400 ;
        RECT 159.600 335.800 162.000 336.600 ;
        RECT 148.400 333.600 149.200 335.200 ;
        RECT 150.000 334.800 150.800 335.000 ;
        RECT 150.000 334.200 154.400 334.800 ;
        RECT 153.600 334.000 154.400 334.200 ;
        RECT 135.600 327.400 136.400 333.000 ;
        RECT 145.000 332.600 147.000 333.400 ;
        RECT 150.800 332.600 154.000 333.400 ;
        RECT 156.400 332.800 157.200 335.600 ;
        RECT 161.200 335.200 162.000 335.800 ;
        RECT 161.200 334.600 163.000 335.200 ;
        RECT 162.200 333.400 163.000 334.600 ;
        RECT 166.000 334.600 166.800 339.800 ;
        RECT 167.600 336.000 168.400 339.800 ;
        RECT 167.600 335.200 168.600 336.000 ;
        RECT 166.000 334.000 167.200 334.600 ;
        RECT 162.200 332.600 166.000 333.400 ;
        RECT 137.000 332.000 137.800 332.200 ;
        RECT 140.400 332.000 141.200 332.400 ;
        RECT 142.000 332.000 142.800 332.400 ;
        RECT 159.600 332.000 160.400 332.600 ;
        RECT 166.600 332.000 167.200 334.000 ;
        RECT 137.000 331.400 160.400 332.000 ;
        RECT 166.400 331.400 167.200 332.000 ;
        RECT 166.400 329.600 167.000 331.400 ;
        RECT 167.800 330.800 168.600 335.200 ;
        RECT 169.200 334.300 170.000 334.400 ;
        RECT 170.800 334.300 171.600 339.800 ;
        RECT 174.000 335.200 174.800 339.800 ;
        RECT 175.600 335.800 176.400 339.800 ;
        RECT 177.200 336.000 178.000 339.800 ;
        RECT 180.400 336.000 181.200 339.800 ;
        RECT 177.200 335.800 181.200 336.000 ;
        RECT 169.200 333.700 171.600 334.300 ;
        RECT 169.200 333.600 170.000 333.700 ;
        RECT 145.200 329.400 146.000 329.600 ;
        RECT 140.600 329.000 146.000 329.400 ;
        RECT 139.800 328.800 146.000 329.000 ;
        RECT 147.000 329.000 155.600 329.600 ;
        RECT 137.200 328.000 138.800 328.800 ;
        RECT 139.800 328.200 141.200 328.800 ;
        RECT 147.000 328.200 147.600 329.000 ;
        RECT 154.800 328.800 155.600 329.000 ;
        RECT 158.000 329.000 167.000 329.600 ;
        RECT 158.000 328.800 158.800 329.000 ;
        RECT 138.200 327.600 138.800 328.000 ;
        RECT 141.800 327.600 147.600 328.200 ;
        RECT 148.200 327.600 150.800 328.400 ;
        RECT 135.600 326.800 137.600 327.400 ;
        RECT 138.200 326.800 142.400 327.600 ;
        RECT 118.000 322.200 118.800 325.000 ;
        RECT 119.600 322.200 120.400 325.000 ;
        RECT 122.800 322.200 123.600 326.800 ;
        RECT 126.400 326.200 127.000 326.800 ;
        RECT 126.000 325.600 127.000 326.200 ;
        RECT 137.000 326.200 137.600 326.800 ;
        RECT 137.000 325.600 138.000 326.200 ;
        RECT 126.000 322.200 126.800 325.600 ;
        RECT 137.200 322.200 138.000 325.600 ;
        RECT 140.400 322.200 141.200 326.800 ;
        RECT 143.600 322.200 144.400 325.000 ;
        RECT 145.200 322.200 146.000 325.000 ;
        RECT 146.800 322.200 147.600 327.000 ;
        RECT 150.000 322.200 150.800 327.000 ;
        RECT 153.200 322.200 154.000 328.400 ;
        RECT 161.200 327.600 163.800 328.400 ;
        RECT 156.400 326.800 160.600 327.600 ;
        RECT 154.800 322.200 155.600 325.000 ;
        RECT 156.400 322.200 157.200 325.000 ;
        RECT 158.000 322.200 158.800 325.000 ;
        RECT 161.200 322.200 162.000 327.600 ;
        RECT 166.400 327.400 167.000 329.000 ;
        RECT 164.400 326.800 167.000 327.400 ;
        RECT 167.600 330.000 168.600 330.800 ;
        RECT 170.800 332.400 171.600 333.700 ;
        RECT 172.600 334.600 174.800 335.200 ;
        RECT 170.800 330.200 171.400 332.400 ;
        RECT 172.600 331.600 173.200 334.600 ;
        RECT 175.800 334.400 176.400 335.800 ;
        RECT 177.400 335.400 181.000 335.800 ;
        RECT 182.000 335.600 182.800 337.200 ;
        RECT 179.600 334.400 180.400 334.800 ;
        RECT 175.600 333.600 178.200 334.400 ;
        RECT 179.600 334.300 181.200 334.400 ;
        RECT 183.600 334.300 184.400 339.800 ;
        RECT 179.600 333.800 184.400 334.300 ;
        RECT 188.800 334.200 189.600 339.800 ;
        RECT 191.600 335.600 192.400 337.200 ;
        RECT 193.200 334.300 194.000 339.800 ;
        RECT 194.800 336.000 195.600 339.800 ;
        RECT 198.000 336.000 198.800 339.800 ;
        RECT 194.800 335.800 198.800 336.000 ;
        RECT 199.600 335.800 200.400 339.800 ;
        RECT 203.800 336.400 204.600 339.800 ;
        RECT 202.800 335.800 204.600 336.400 ;
        RECT 195.000 335.400 198.600 335.800 ;
        RECT 195.600 334.400 196.400 334.800 ;
        RECT 199.600 334.400 200.200 335.800 ;
        RECT 194.800 334.300 196.400 334.400 ;
        RECT 188.800 333.800 190.600 334.200 ;
        RECT 180.400 333.700 184.400 333.800 ;
        RECT 180.400 333.600 181.200 333.700 ;
        RECT 172.000 330.800 173.200 331.600 ;
        RECT 172.600 330.200 173.200 330.800 ;
        RECT 175.600 330.200 176.400 330.400 ;
        RECT 177.600 330.200 178.200 333.600 ;
        RECT 178.800 332.300 179.600 333.200 ;
        RECT 180.400 332.300 181.200 332.400 ;
        RECT 178.800 331.700 181.200 332.300 ;
        RECT 178.800 331.600 179.600 331.700 ;
        RECT 180.400 331.600 181.200 331.700 ;
        RECT 183.600 330.300 184.400 333.700 ;
        RECT 189.000 333.600 190.600 333.800 ;
        RECT 186.800 331.600 188.400 332.400 ;
        RECT 185.200 330.300 186.000 331.200 ;
        RECT 164.400 322.200 165.200 326.800 ;
        RECT 167.600 322.200 168.400 330.000 ;
        RECT 170.800 322.200 171.600 330.200 ;
        RECT 172.600 329.600 174.800 330.200 ;
        RECT 175.600 329.600 177.000 330.200 ;
        RECT 177.600 329.600 178.600 330.200 ;
        RECT 174.000 322.200 174.800 329.600 ;
        RECT 176.400 328.400 177.000 329.600 ;
        RECT 176.400 327.600 177.200 328.400 ;
        RECT 177.800 322.200 178.600 329.600 ;
        RECT 183.600 329.700 186.000 330.300 ;
        RECT 183.600 322.200 184.400 329.700 ;
        RECT 185.200 329.600 186.000 329.700 ;
        RECT 190.000 330.400 190.600 333.600 ;
        RECT 193.200 333.800 196.400 334.300 ;
        RECT 193.200 333.700 195.600 333.800 ;
        RECT 190.000 329.600 190.800 330.400 ;
        RECT 188.400 327.600 189.200 329.200 ;
        RECT 190.000 327.000 190.600 329.600 ;
        RECT 187.000 326.400 190.600 327.000 ;
        RECT 187.000 326.200 187.600 326.400 ;
        RECT 186.800 322.200 187.600 326.200 ;
        RECT 190.000 326.200 190.600 326.400 ;
        RECT 190.000 322.200 190.800 326.200 ;
        RECT 193.200 322.200 194.000 333.700 ;
        RECT 194.800 333.600 195.600 333.700 ;
        RECT 197.800 333.600 200.400 334.400 ;
        RECT 201.200 333.600 202.000 335.200 ;
        RECT 196.400 331.600 197.200 333.200 ;
        RECT 197.800 330.200 198.400 333.600 ;
        RECT 199.600 330.200 200.400 330.400 ;
        RECT 197.400 329.600 198.400 330.200 ;
        RECT 199.000 329.600 200.400 330.200 ;
        RECT 197.400 322.200 198.200 329.600 ;
        RECT 199.000 328.400 199.600 329.600 ;
        RECT 198.800 327.600 199.600 328.400 ;
        RECT 202.800 322.200 203.600 335.800 ;
        RECT 206.000 335.200 206.800 339.800 ;
        RECT 206.000 334.600 208.200 335.200 ;
        RECT 207.600 331.600 208.200 334.600 ;
        RECT 209.200 332.400 210.000 339.800 ;
        RECT 207.600 330.800 208.800 331.600 ;
        RECT 204.400 328.800 205.200 330.400 ;
        RECT 207.600 330.200 208.200 330.800 ;
        RECT 209.400 330.200 210.000 332.400 ;
        RECT 206.000 329.600 208.200 330.200 ;
        RECT 206.000 322.200 206.800 329.600 ;
        RECT 209.200 322.200 210.000 330.200 ;
        RECT 210.800 322.200 211.600 339.800 ;
        RECT 215.600 337.800 216.400 339.800 ;
        RECT 212.400 335.600 213.200 337.200 ;
        RECT 214.000 335.600 214.800 337.200 ;
        RECT 212.500 334.400 213.100 335.600 ;
        RECT 215.800 334.400 216.400 337.800 ;
        RECT 220.400 336.000 221.200 339.800 ;
        RECT 212.400 334.300 213.200 334.400 ;
        RECT 215.600 334.300 216.400 334.400 ;
        RECT 212.400 333.700 216.400 334.300 ;
        RECT 212.400 333.600 213.200 333.700 ;
        RECT 215.600 333.600 216.400 333.700 ;
        RECT 215.800 330.200 216.400 333.600 ;
        RECT 220.200 335.200 221.200 336.000 ;
        RECT 217.200 332.300 218.000 332.400 ;
        RECT 220.200 332.300 221.000 335.200 ;
        RECT 222.000 334.600 222.800 339.800 ;
        RECT 228.400 336.600 229.200 339.800 ;
        RECT 230.000 337.000 230.800 339.800 ;
        RECT 231.600 337.000 232.400 339.800 ;
        RECT 233.200 337.000 234.000 339.800 ;
        RECT 234.800 337.000 235.600 339.800 ;
        RECT 238.000 337.000 238.800 339.800 ;
        RECT 241.200 337.000 242.000 339.800 ;
        RECT 242.800 337.000 243.600 339.800 ;
        RECT 244.400 337.000 245.200 339.800 ;
        RECT 226.800 335.800 229.200 336.600 ;
        RECT 246.000 336.600 246.800 339.800 ;
        RECT 226.800 335.200 227.600 335.800 ;
        RECT 217.200 331.700 221.000 332.300 ;
        RECT 217.200 330.800 218.000 331.700 ;
        RECT 220.200 330.800 221.000 331.700 ;
        RECT 221.600 334.000 222.800 334.600 ;
        RECT 225.800 334.600 227.600 335.200 ;
        RECT 231.600 335.600 232.600 336.400 ;
        RECT 235.600 335.600 237.200 336.400 ;
        RECT 238.000 335.800 242.600 336.400 ;
        RECT 246.000 335.800 248.600 336.600 ;
        RECT 238.000 335.600 238.800 335.800 ;
        RECT 221.600 332.000 222.200 334.000 ;
        RECT 225.800 333.400 226.600 334.600 ;
        RECT 222.800 332.600 226.600 333.400 ;
        RECT 231.600 332.800 232.400 335.600 ;
        RECT 238.000 334.800 238.800 335.000 ;
        RECT 234.400 334.200 238.800 334.800 ;
        RECT 234.400 334.000 235.200 334.200 ;
        RECT 239.600 333.600 240.400 335.200 ;
        RECT 241.800 333.400 242.600 335.800 ;
        RECT 247.800 335.200 248.600 335.800 ;
        RECT 247.800 334.400 250.800 335.200 ;
        RECT 252.400 333.800 253.200 339.800 ;
        RECT 255.600 335.200 256.400 339.800 ;
        RECT 258.800 335.200 259.600 339.800 ;
        RECT 262.000 335.200 262.800 339.800 ;
        RECT 265.200 335.200 266.000 339.800 ;
        RECT 255.600 334.400 257.400 335.200 ;
        RECT 258.800 334.400 261.000 335.200 ;
        RECT 262.000 334.400 264.200 335.200 ;
        RECT 265.200 334.400 267.600 335.200 ;
        RECT 234.800 332.600 238.000 333.400 ;
        RECT 241.800 332.600 243.800 333.400 ;
        RECT 244.400 333.000 253.200 333.800 ;
        RECT 228.400 332.000 229.200 332.600 ;
        RECT 246.000 332.000 246.800 332.400 ;
        RECT 251.000 332.000 251.800 332.200 ;
        RECT 221.600 331.400 222.400 332.000 ;
        RECT 228.400 331.400 251.800 332.000 ;
        RECT 215.600 329.400 217.400 330.200 ;
        RECT 220.200 330.000 221.200 330.800 ;
        RECT 216.600 322.200 217.400 329.400 ;
        RECT 220.400 322.200 221.200 330.000 ;
        RECT 221.800 329.600 222.400 331.400 ;
        RECT 221.800 329.000 230.800 329.600 ;
        RECT 221.800 327.400 222.400 329.000 ;
        RECT 230.000 328.800 230.800 329.000 ;
        RECT 233.200 329.000 241.800 329.600 ;
        RECT 233.200 328.800 234.000 329.000 ;
        RECT 225.000 327.600 227.600 328.400 ;
        RECT 221.800 326.800 224.400 327.400 ;
        RECT 223.600 322.200 224.400 326.800 ;
        RECT 226.800 322.200 227.600 327.600 ;
        RECT 228.200 326.800 232.400 327.600 ;
        RECT 230.000 322.200 230.800 325.000 ;
        RECT 231.600 322.200 232.400 325.000 ;
        RECT 233.200 322.200 234.000 325.000 ;
        RECT 234.800 322.200 235.600 328.400 ;
        RECT 238.000 327.600 240.600 328.400 ;
        RECT 241.200 328.200 241.800 329.000 ;
        RECT 242.800 329.400 243.600 329.600 ;
        RECT 242.800 329.000 248.200 329.400 ;
        RECT 242.800 328.800 249.000 329.000 ;
        RECT 247.600 328.200 249.000 328.800 ;
        RECT 241.200 327.600 247.000 328.200 ;
        RECT 250.000 328.000 251.600 328.800 ;
        RECT 250.000 327.600 250.600 328.000 ;
        RECT 238.000 322.200 238.800 327.000 ;
        RECT 241.200 322.200 242.000 327.000 ;
        RECT 246.400 326.800 250.600 327.600 ;
        RECT 252.400 327.400 253.200 333.000 ;
        RECT 256.600 333.800 257.400 334.400 ;
        RECT 260.200 333.800 261.000 334.400 ;
        RECT 263.400 333.800 264.200 334.400 ;
        RECT 256.600 333.000 259.200 333.800 ;
        RECT 260.200 333.000 262.600 333.800 ;
        RECT 263.400 333.000 266.000 333.800 ;
        RECT 256.600 331.600 257.400 333.000 ;
        RECT 260.200 331.600 261.000 333.000 ;
        RECT 263.400 331.600 264.200 333.000 ;
        RECT 266.800 331.600 267.600 334.400 ;
        RECT 251.200 326.800 253.200 327.400 ;
        RECT 255.600 330.800 257.400 331.600 ;
        RECT 258.800 330.800 261.000 331.600 ;
        RECT 262.000 330.800 264.200 331.600 ;
        RECT 265.200 330.800 267.600 331.600 ;
        RECT 274.800 333.800 275.600 339.800 ;
        RECT 281.200 336.600 282.000 339.800 ;
        RECT 282.800 337.000 283.600 339.800 ;
        RECT 284.400 337.000 285.200 339.800 ;
        RECT 286.000 337.000 286.800 339.800 ;
        RECT 289.200 337.000 290.000 339.800 ;
        RECT 292.400 337.000 293.200 339.800 ;
        RECT 294.000 337.000 294.800 339.800 ;
        RECT 295.600 337.000 296.400 339.800 ;
        RECT 297.200 337.000 298.000 339.800 ;
        RECT 279.400 335.800 282.000 336.600 ;
        RECT 298.800 336.600 299.600 339.800 ;
        RECT 285.400 335.800 290.000 336.400 ;
        RECT 279.400 335.200 280.200 335.800 ;
        RECT 277.200 334.400 280.200 335.200 ;
        RECT 274.800 333.000 283.600 333.800 ;
        RECT 285.400 333.400 286.200 335.800 ;
        RECT 289.200 335.600 290.000 335.800 ;
        RECT 290.800 335.600 292.400 336.400 ;
        RECT 295.400 335.600 296.400 336.400 ;
        RECT 298.800 335.800 301.200 336.600 ;
        RECT 287.600 333.600 288.400 335.200 ;
        RECT 289.200 334.800 290.000 335.000 ;
        RECT 289.200 334.200 293.600 334.800 ;
        RECT 292.800 334.000 293.600 334.200 ;
        RECT 242.800 322.200 243.600 325.000 ;
        RECT 244.400 322.200 245.200 325.000 ;
        RECT 247.600 322.200 248.400 326.800 ;
        RECT 251.200 326.200 251.800 326.800 ;
        RECT 250.800 325.600 251.800 326.200 ;
        RECT 250.800 322.200 251.600 325.600 ;
        RECT 255.600 322.200 256.400 330.800 ;
        RECT 258.800 322.200 259.600 330.800 ;
        RECT 262.000 322.200 262.800 330.800 ;
        RECT 265.200 322.200 266.000 330.800 ;
        RECT 274.800 327.400 275.600 333.000 ;
        RECT 284.200 332.600 286.200 333.400 ;
        RECT 290.000 332.600 293.200 333.400 ;
        RECT 295.600 332.800 296.400 335.600 ;
        RECT 300.400 335.200 301.200 335.800 ;
        RECT 300.400 334.600 302.200 335.200 ;
        RECT 301.400 333.400 302.200 334.600 ;
        RECT 305.200 334.600 306.000 339.800 ;
        RECT 306.800 336.000 307.600 339.800 ;
        RECT 306.800 335.200 307.800 336.000 ;
        RECT 305.200 334.000 306.400 334.600 ;
        RECT 301.400 332.600 305.200 333.400 ;
        RECT 276.200 332.000 277.000 332.200 ;
        RECT 281.200 332.000 282.000 332.400 ;
        RECT 298.800 332.000 299.600 332.600 ;
        RECT 305.800 332.000 306.400 334.000 ;
        RECT 276.200 331.400 299.600 332.000 ;
        RECT 305.600 331.400 306.400 332.000 ;
        RECT 305.600 329.600 306.200 331.400 ;
        RECT 307.000 330.800 307.800 335.200 ;
        RECT 284.400 329.400 285.200 329.600 ;
        RECT 279.800 329.000 285.200 329.400 ;
        RECT 279.000 328.800 285.200 329.000 ;
        RECT 286.200 329.000 294.800 329.600 ;
        RECT 276.400 328.000 278.000 328.800 ;
        RECT 279.000 328.200 280.400 328.800 ;
        RECT 286.200 328.200 286.800 329.000 ;
        RECT 294.000 328.800 294.800 329.000 ;
        RECT 297.200 329.000 306.200 329.600 ;
        RECT 297.200 328.800 298.000 329.000 ;
        RECT 277.400 327.600 278.000 328.000 ;
        RECT 281.000 327.600 286.800 328.200 ;
        RECT 287.400 327.600 290.000 328.400 ;
        RECT 274.800 326.800 276.800 327.400 ;
        RECT 277.400 326.800 281.600 327.600 ;
        RECT 276.200 326.200 276.800 326.800 ;
        RECT 276.200 325.600 277.200 326.200 ;
        RECT 276.400 322.200 277.200 325.600 ;
        RECT 279.600 322.200 280.400 326.800 ;
        RECT 282.800 322.200 283.600 325.000 ;
        RECT 284.400 322.200 285.200 325.000 ;
        RECT 286.000 322.200 286.800 327.000 ;
        RECT 289.200 322.200 290.000 327.000 ;
        RECT 292.400 322.200 293.200 328.400 ;
        RECT 300.400 327.600 303.000 328.400 ;
        RECT 295.600 326.800 299.800 327.600 ;
        RECT 294.000 322.200 294.800 325.000 ;
        RECT 295.600 322.200 296.400 325.000 ;
        RECT 297.200 322.200 298.000 325.000 ;
        RECT 300.400 322.200 301.200 327.600 ;
        RECT 305.600 327.400 306.200 329.000 ;
        RECT 303.600 326.800 306.200 327.400 ;
        RECT 306.800 330.000 307.800 330.800 ;
        RECT 310.000 333.800 310.800 339.800 ;
        RECT 316.400 336.600 317.200 339.800 ;
        RECT 318.000 337.000 318.800 339.800 ;
        RECT 319.600 337.000 320.400 339.800 ;
        RECT 321.200 337.000 322.000 339.800 ;
        RECT 324.400 337.000 325.200 339.800 ;
        RECT 327.600 337.000 328.400 339.800 ;
        RECT 329.200 337.000 330.000 339.800 ;
        RECT 330.800 337.000 331.600 339.800 ;
        RECT 332.400 337.000 333.200 339.800 ;
        RECT 314.600 335.800 317.200 336.600 ;
        RECT 334.000 336.600 334.800 339.800 ;
        RECT 320.600 335.800 325.200 336.400 ;
        RECT 314.600 335.200 315.400 335.800 ;
        RECT 312.400 334.400 315.400 335.200 ;
        RECT 310.000 333.000 318.800 333.800 ;
        RECT 320.600 333.400 321.400 335.800 ;
        RECT 324.400 335.600 325.200 335.800 ;
        RECT 326.000 335.600 327.600 336.400 ;
        RECT 330.600 335.600 331.600 336.400 ;
        RECT 334.000 335.800 336.400 336.600 ;
        RECT 322.800 333.600 323.600 335.200 ;
        RECT 324.400 334.800 325.200 335.000 ;
        RECT 324.400 334.200 328.800 334.800 ;
        RECT 328.000 334.000 328.800 334.200 ;
        RECT 303.600 322.200 304.400 326.800 ;
        RECT 306.800 322.200 307.600 330.000 ;
        RECT 310.000 327.400 310.800 333.000 ;
        RECT 319.400 332.600 321.400 333.400 ;
        RECT 325.200 332.600 328.400 333.400 ;
        RECT 330.800 332.800 331.600 335.600 ;
        RECT 335.600 335.200 336.400 335.800 ;
        RECT 335.600 334.600 337.400 335.200 ;
        RECT 336.600 333.400 337.400 334.600 ;
        RECT 340.400 334.600 341.200 339.800 ;
        RECT 342.000 336.000 342.800 339.800 ;
        RECT 342.000 335.200 343.000 336.000 ;
        RECT 340.400 334.000 341.600 334.600 ;
        RECT 336.600 332.600 340.400 333.400 ;
        RECT 311.600 332.200 312.400 332.400 ;
        RECT 311.400 332.000 312.400 332.200 ;
        RECT 314.800 332.000 315.600 332.400 ;
        RECT 316.400 332.000 317.200 332.400 ;
        RECT 334.000 332.000 334.800 332.600 ;
        RECT 341.000 332.000 341.600 334.000 ;
        RECT 311.400 331.400 334.800 332.000 ;
        RECT 340.800 331.400 341.600 332.000 ;
        RECT 340.800 329.600 341.400 331.400 ;
        RECT 342.200 330.800 343.000 335.200 ;
        RECT 343.600 334.300 344.400 334.400 ;
        RECT 345.200 334.300 346.000 335.200 ;
        RECT 343.600 333.700 346.000 334.300 ;
        RECT 343.600 333.600 344.400 333.700 ;
        RECT 345.200 333.600 346.000 333.700 ;
        RECT 319.600 329.400 320.400 329.600 ;
        RECT 315.000 329.000 320.400 329.400 ;
        RECT 314.200 328.800 320.400 329.000 ;
        RECT 321.400 329.000 330.000 329.600 ;
        RECT 311.600 328.000 313.200 328.800 ;
        RECT 314.200 328.200 315.600 328.800 ;
        RECT 321.400 328.200 322.000 329.000 ;
        RECT 329.200 328.800 330.000 329.000 ;
        RECT 332.400 329.000 341.400 329.600 ;
        RECT 332.400 328.800 333.200 329.000 ;
        RECT 312.600 327.600 313.200 328.000 ;
        RECT 316.200 327.600 322.000 328.200 ;
        RECT 322.600 327.600 325.200 328.400 ;
        RECT 310.000 326.800 312.000 327.400 ;
        RECT 312.600 326.800 316.800 327.600 ;
        RECT 311.400 326.200 312.000 326.800 ;
        RECT 311.400 325.600 312.400 326.200 ;
        RECT 311.600 322.200 312.400 325.600 ;
        RECT 314.800 322.200 315.600 326.800 ;
        RECT 318.000 322.200 318.800 325.000 ;
        RECT 319.600 322.200 320.400 325.000 ;
        RECT 321.200 322.200 322.000 327.000 ;
        RECT 324.400 322.200 325.200 327.000 ;
        RECT 327.600 322.200 328.400 328.400 ;
        RECT 335.600 327.600 338.200 328.400 ;
        RECT 330.800 326.800 335.000 327.600 ;
        RECT 329.200 322.200 330.000 325.000 ;
        RECT 330.800 322.200 331.600 325.000 ;
        RECT 332.400 322.200 333.200 325.000 ;
        RECT 335.600 322.200 336.400 327.600 ;
        RECT 340.800 327.400 341.400 329.000 ;
        RECT 338.800 326.800 341.400 327.400 ;
        RECT 342.000 330.000 343.000 330.800 ;
        RECT 342.000 328.300 342.800 330.000 ;
        RECT 343.600 328.300 344.400 328.400 ;
        RECT 342.000 327.700 344.400 328.300 ;
        RECT 338.800 322.200 339.600 326.800 ;
        RECT 342.000 322.200 342.800 327.700 ;
        RECT 343.600 327.600 344.400 327.700 ;
        RECT 346.800 322.200 347.600 339.800 ;
        RECT 351.000 338.400 351.800 339.800 ;
        RECT 351.000 337.600 352.400 338.400 ;
        RECT 351.000 336.400 351.800 337.600 ;
        RECT 350.000 335.800 351.800 336.400 ;
        RECT 348.400 333.600 349.200 335.200 ;
        RECT 350.000 322.200 350.800 335.800 ;
        RECT 356.400 335.600 357.200 339.800 ;
        RECT 357.800 336.400 358.600 337.200 ;
        RECT 358.000 336.300 358.800 336.400 ;
        RECT 359.600 336.300 360.400 339.800 ;
        RECT 358.000 335.700 360.400 336.300 ;
        RECT 361.200 336.000 362.000 339.800 ;
        RECT 364.400 336.000 365.200 339.800 ;
        RECT 361.200 335.800 365.200 336.000 ;
        RECT 366.000 335.800 366.800 339.800 ;
        RECT 367.600 336.000 368.400 339.800 ;
        RECT 370.800 336.000 371.600 339.800 ;
        RECT 367.600 335.800 371.600 336.000 ;
        RECT 358.000 335.600 358.800 335.700 ;
        RECT 354.800 332.800 355.600 334.400 ;
        RECT 353.200 332.200 354.000 332.400 ;
        RECT 356.400 332.200 357.000 335.600 ;
        RECT 359.800 334.400 360.400 335.700 ;
        RECT 361.400 335.400 365.000 335.800 ;
        RECT 363.600 334.400 364.400 334.800 ;
        RECT 366.200 334.400 366.800 335.800 ;
        RECT 367.800 335.400 371.400 335.800 ;
        RECT 370.000 334.400 370.800 334.800 ;
        RECT 359.600 333.600 362.200 334.400 ;
        RECT 363.600 333.800 365.200 334.400 ;
        RECT 364.400 333.600 365.200 333.800 ;
        RECT 366.000 333.600 368.600 334.400 ;
        RECT 370.000 334.300 371.600 334.400 ;
        RECT 372.400 334.300 373.200 339.800 ;
        RECT 374.000 335.600 374.800 337.200 ;
        RECT 376.200 336.400 377.000 339.800 ;
        RECT 383.000 338.400 383.800 339.800 ;
        RECT 382.000 337.600 383.800 338.400 ;
        RECT 383.000 336.400 383.800 337.600 ;
        RECT 376.200 335.800 378.000 336.400 ;
        RECT 370.000 333.800 373.200 334.300 ;
        RECT 370.800 333.700 373.200 333.800 ;
        RECT 370.800 333.600 371.600 333.700 ;
        RECT 358.000 332.200 358.800 332.400 ;
        RECT 353.200 331.600 354.800 332.200 ;
        RECT 356.400 331.600 358.800 332.200 ;
        RECT 354.000 331.200 354.800 331.600 ;
        RECT 351.600 328.800 352.400 330.400 ;
        RECT 358.000 330.200 358.600 331.600 ;
        RECT 359.600 330.200 360.400 330.400 ;
        RECT 361.600 330.200 362.200 333.600 ;
        RECT 362.800 331.600 363.600 333.200 ;
        RECT 366.000 330.200 366.800 330.400 ;
        RECT 368.000 330.200 368.600 333.600 ;
        RECT 369.200 332.300 370.000 333.200 ;
        RECT 370.800 332.300 371.600 332.400 ;
        RECT 369.200 331.700 371.600 332.300 ;
        RECT 369.200 331.600 370.000 331.700 ;
        RECT 370.800 331.600 371.600 331.700 ;
        RECT 353.200 329.600 357.200 330.200 ;
        RECT 353.200 322.200 354.000 329.600 ;
        RECT 356.400 322.200 357.200 329.600 ;
        RECT 358.000 322.200 358.800 330.200 ;
        RECT 359.600 329.600 361.000 330.200 ;
        RECT 361.600 329.600 362.600 330.200 ;
        RECT 366.000 329.600 367.400 330.200 ;
        RECT 368.000 329.600 369.000 330.200 ;
        RECT 360.400 328.400 361.000 329.600 ;
        RECT 360.400 327.600 361.200 328.400 ;
        RECT 361.800 322.200 362.600 329.600 ;
        RECT 366.800 328.400 367.400 329.600 ;
        RECT 366.800 327.600 367.600 328.400 ;
        RECT 368.200 324.400 369.000 329.600 ;
        RECT 368.200 323.600 370.000 324.400 ;
        RECT 368.200 322.200 369.000 323.600 ;
        RECT 372.400 322.200 373.200 333.700 ;
        RECT 374.000 334.300 374.800 334.400 ;
        RECT 377.200 334.300 378.000 335.800 ;
        RECT 382.000 335.800 383.800 336.400 ;
        RECT 374.000 333.700 378.000 334.300 ;
        RECT 374.000 333.600 374.800 333.700 ;
        RECT 375.600 328.800 376.400 330.400 ;
        RECT 377.200 322.200 378.000 333.700 ;
        RECT 378.800 334.300 379.600 335.200 ;
        RECT 380.400 334.300 381.200 335.200 ;
        RECT 378.800 333.700 381.200 334.300 ;
        RECT 378.800 333.600 379.600 333.700 ;
        RECT 380.400 333.600 381.200 333.700 ;
        RECT 382.000 334.300 382.800 335.800 ;
        RECT 385.200 334.300 386.000 335.200 ;
        RECT 382.000 333.700 386.000 334.300 ;
        RECT 382.000 322.200 382.800 333.700 ;
        RECT 385.200 333.600 386.000 333.700 ;
        RECT 383.600 328.800 384.400 330.400 ;
        RECT 386.800 322.200 387.600 339.800 ;
        RECT 388.400 335.800 389.200 339.800 ;
        RECT 390.000 336.000 390.800 339.800 ;
        RECT 393.200 336.000 394.000 339.800 ;
        RECT 395.400 338.400 396.200 339.800 ;
        RECT 394.800 337.600 396.200 338.400 ;
        RECT 390.000 335.800 394.000 336.000 ;
        RECT 395.400 336.400 396.200 337.600 ;
        RECT 400.200 336.400 401.000 339.800 ;
        RECT 395.400 335.800 397.200 336.400 ;
        RECT 400.200 335.800 402.000 336.400 ;
        RECT 404.400 335.800 405.200 339.800 ;
        RECT 406.000 336.000 406.800 339.800 ;
        RECT 409.200 336.000 410.000 339.800 ;
        RECT 406.000 335.800 410.000 336.000 ;
        RECT 412.400 337.600 413.200 339.800 ;
        RECT 388.600 334.400 389.200 335.800 ;
        RECT 390.200 335.400 393.800 335.800 ;
        RECT 392.400 334.400 393.200 334.800 ;
        RECT 388.400 333.600 391.000 334.400 ;
        RECT 392.400 333.800 394.000 334.400 ;
        RECT 393.200 333.600 394.000 333.800 ;
        RECT 388.400 330.200 389.200 330.400 ;
        RECT 390.400 330.200 391.000 333.600 ;
        RECT 391.600 331.600 392.400 333.200 ;
        RECT 388.400 329.600 389.800 330.200 ;
        RECT 390.400 329.600 391.400 330.200 ;
        RECT 389.200 328.400 389.800 329.600 ;
        RECT 389.200 327.600 390.000 328.400 ;
        RECT 390.600 322.200 391.400 329.600 ;
        RECT 394.800 328.800 395.600 330.400 ;
        RECT 396.400 322.200 397.200 335.800 ;
        RECT 398.000 333.600 398.800 335.200 ;
        RECT 398.000 330.300 398.800 330.400 ;
        RECT 399.600 330.300 400.400 330.400 ;
        RECT 398.000 329.700 400.400 330.300 ;
        RECT 398.000 329.600 398.800 329.700 ;
        RECT 399.600 328.800 400.400 329.700 ;
        RECT 401.200 330.300 402.000 335.800 ;
        RECT 402.800 333.600 403.600 335.200 ;
        RECT 404.600 334.400 405.200 335.800 ;
        RECT 406.200 335.400 409.800 335.800 ;
        RECT 408.400 334.400 409.200 334.800 ;
        RECT 412.400 334.400 413.000 337.600 ;
        RECT 414.000 336.300 414.800 337.200 ;
        RECT 415.600 336.300 416.400 339.800 ;
        RECT 428.400 338.400 429.200 339.800 ;
        RECT 428.400 337.600 429.400 338.400 ;
        RECT 431.600 337.800 432.400 339.800 ;
        RECT 431.600 337.600 432.800 337.800 ;
        RECT 414.000 335.700 416.400 336.300 ;
        RECT 414.000 335.600 414.800 335.700 ;
        RECT 404.400 333.600 407.000 334.400 ;
        RECT 408.400 333.800 410.000 334.400 ;
        RECT 409.200 333.600 410.000 333.800 ;
        RECT 412.400 333.600 413.200 334.400 ;
        RECT 404.400 330.300 405.200 330.400 ;
        RECT 401.200 330.200 405.200 330.300 ;
        RECT 406.400 330.200 407.000 333.600 ;
        RECT 407.600 331.600 408.400 333.200 ;
        RECT 409.300 332.300 409.900 333.600 ;
        RECT 410.800 332.300 411.600 332.400 ;
        RECT 409.300 331.700 411.600 332.300 ;
        RECT 410.800 330.800 411.600 331.700 ;
        RECT 412.400 330.200 413.000 333.600 ;
        RECT 414.000 332.300 414.800 332.400 ;
        RECT 415.600 332.300 416.400 335.700 ;
        RECT 417.200 336.300 418.000 337.200 ;
        RECT 428.800 337.000 432.800 337.600 ;
        RECT 418.800 336.300 419.600 336.400 ;
        RECT 423.600 336.300 424.400 336.400 ;
        RECT 426.800 336.300 428.600 336.400 ;
        RECT 417.200 335.700 428.600 336.300 ;
        RECT 417.200 335.600 418.000 335.700 ;
        RECT 418.800 335.600 419.600 335.700 ;
        RECT 423.600 335.600 424.400 335.700 ;
        RECT 426.800 335.600 428.600 335.700 ;
        RECT 417.200 334.300 418.000 334.400 ;
        RECT 428.400 334.300 430.000 334.400 ;
        RECT 417.200 333.700 430.000 334.300 ;
        RECT 417.200 333.600 418.000 333.700 ;
        RECT 428.400 333.600 430.000 333.700 ;
        RECT 414.000 331.700 416.400 332.300 ;
        RECT 414.000 331.600 414.800 331.700 ;
        RECT 401.200 329.700 405.800 330.200 ;
        RECT 401.200 322.200 402.000 329.700 ;
        RECT 404.400 329.600 405.800 329.700 ;
        RECT 406.400 329.600 407.400 330.200 ;
        RECT 405.200 328.400 405.800 329.600 ;
        RECT 405.200 327.600 406.000 328.400 ;
        RECT 406.600 326.400 407.400 329.600 ;
        RECT 411.400 329.400 413.200 330.200 ;
        RECT 406.600 325.600 408.400 326.400 ;
        RECT 406.600 322.200 407.400 325.600 ;
        RECT 411.400 322.200 412.200 329.400 ;
        RECT 415.600 322.200 416.400 331.700 ;
        RECT 430.000 331.600 431.600 332.400 ;
        RECT 432.200 330.400 432.800 337.000 ;
        RECT 441.600 334.200 442.400 339.800 ;
        RECT 444.400 335.800 445.200 339.800 ;
        RECT 446.000 336.000 446.800 339.800 ;
        RECT 449.200 336.000 450.000 339.800 ;
        RECT 446.000 335.800 450.000 336.000 ;
        RECT 444.600 334.400 445.200 335.800 ;
        RECT 446.200 335.400 449.800 335.800 ;
        RECT 448.400 334.400 449.200 334.800 ;
        RECT 441.600 333.800 443.400 334.200 ;
        RECT 441.800 333.600 443.400 333.800 ;
        RECT 444.400 333.600 447.000 334.400 ;
        RECT 448.400 333.800 450.000 334.400 ;
        RECT 449.200 333.600 450.000 333.800 ;
        RECT 439.600 331.600 441.200 332.400 ;
        RECT 432.200 329.800 435.600 330.400 ;
        RECT 434.800 329.600 435.600 329.800 ;
        RECT 438.000 329.600 438.800 331.200 ;
        RECT 442.800 330.400 443.400 333.600 ;
        RECT 446.400 332.400 447.000 333.600 ;
        RECT 446.000 331.600 447.000 332.400 ;
        RECT 447.600 331.600 448.400 333.200 ;
        RECT 442.800 329.600 443.600 330.400 ;
        RECT 444.400 330.200 445.200 330.400 ;
        RECT 446.400 330.200 447.000 331.600 ;
        RECT 444.400 329.600 445.800 330.200 ;
        RECT 446.400 329.600 447.400 330.200 ;
        RECT 425.400 328.800 429.000 329.400 ;
        RECT 425.400 328.200 426.000 328.800 ;
        RECT 425.200 322.200 426.000 328.200 ;
        RECT 428.400 328.200 429.000 328.800 ;
        RECT 430.200 329.000 433.800 329.200 ;
        RECT 434.800 329.000 435.400 329.600 ;
        RECT 430.200 328.600 434.000 329.000 ;
        RECT 430.200 328.200 430.800 328.600 ;
        RECT 428.400 322.800 429.200 328.200 ;
        RECT 430.000 323.400 430.800 328.200 ;
        RECT 431.600 322.800 432.400 328.000 ;
        RECT 433.200 323.000 434.000 328.600 ;
        RECT 434.800 323.400 435.600 329.000 ;
        RECT 428.400 322.200 432.400 322.800 ;
        RECT 433.400 322.800 434.000 323.000 ;
        RECT 436.400 323.000 437.200 329.000 ;
        RECT 441.200 327.600 442.000 329.200 ;
        RECT 442.800 327.000 443.400 329.600 ;
        RECT 445.200 328.400 445.800 329.600 ;
        RECT 445.200 327.600 446.000 328.400 ;
        RECT 439.800 326.400 443.400 327.000 ;
        RECT 439.800 326.200 440.400 326.400 ;
        RECT 436.400 322.800 437.000 323.000 ;
        RECT 433.400 322.200 437.000 322.800 ;
        RECT 439.600 322.200 440.400 326.200 ;
        RECT 442.800 326.200 443.400 326.400 ;
        RECT 442.800 322.200 443.600 326.200 ;
        RECT 446.600 322.200 447.400 329.600 ;
        RECT 450.800 322.200 451.600 339.800 ;
        RECT 455.600 337.800 456.400 339.800 ;
        RECT 452.400 333.600 453.200 335.200 ;
        RECT 455.600 334.400 456.200 337.800 ;
        RECT 457.200 335.600 458.000 337.200 ;
        RECT 455.600 333.600 456.400 334.400 ;
        RECT 458.800 333.800 459.600 339.800 ;
        RECT 465.200 336.600 466.000 339.800 ;
        RECT 466.800 337.000 467.600 339.800 ;
        RECT 468.400 337.000 469.200 339.800 ;
        RECT 470.000 337.000 470.800 339.800 ;
        RECT 473.200 337.000 474.000 339.800 ;
        RECT 476.400 337.000 477.200 339.800 ;
        RECT 478.000 337.000 478.800 339.800 ;
        RECT 479.600 337.000 480.400 339.800 ;
        RECT 481.200 337.000 482.000 339.800 ;
        RECT 463.400 335.800 466.000 336.600 ;
        RECT 482.800 336.600 483.600 339.800 ;
        RECT 469.400 335.800 474.000 336.400 ;
        RECT 463.400 335.200 464.200 335.800 ;
        RECT 461.200 334.400 464.200 335.200 ;
        RECT 452.500 332.400 453.100 333.600 ;
        RECT 455.600 332.400 456.200 333.600 ;
        RECT 458.800 333.000 467.600 333.800 ;
        RECT 469.400 333.400 470.200 335.800 ;
        RECT 473.200 335.600 474.000 335.800 ;
        RECT 474.800 335.600 476.400 336.400 ;
        RECT 479.400 335.600 480.400 336.400 ;
        RECT 482.800 335.800 485.200 336.600 ;
        RECT 471.600 333.600 472.400 335.200 ;
        RECT 473.200 334.800 474.000 335.000 ;
        RECT 473.200 334.200 477.600 334.800 ;
        RECT 476.800 334.000 477.600 334.200 ;
        RECT 452.400 332.300 453.200 332.400 ;
        RECT 454.000 332.300 454.800 332.400 ;
        RECT 452.400 331.700 454.800 332.300 ;
        RECT 452.400 331.600 453.200 331.700 ;
        RECT 454.000 330.800 454.800 331.700 ;
        RECT 455.600 331.600 456.400 332.400 ;
        RECT 455.600 330.200 456.200 331.600 ;
        RECT 454.600 329.400 456.400 330.200 ;
        RECT 454.600 322.200 455.400 329.400 ;
        RECT 458.800 327.400 459.600 333.000 ;
        RECT 468.200 332.600 470.200 333.400 ;
        RECT 474.000 332.600 477.200 333.400 ;
        RECT 479.600 332.800 480.400 335.600 ;
        RECT 484.400 335.200 485.200 335.800 ;
        RECT 484.400 334.600 486.200 335.200 ;
        RECT 485.400 333.400 486.200 334.600 ;
        RECT 489.200 334.600 490.000 339.800 ;
        RECT 490.800 336.000 491.600 339.800 ;
        RECT 494.600 336.400 495.400 339.800 ;
        RECT 490.800 335.200 491.800 336.000 ;
        RECT 494.600 335.800 496.400 336.400 ;
        RECT 498.800 335.800 499.600 339.800 ;
        RECT 500.400 336.000 501.200 339.800 ;
        RECT 503.600 336.000 504.400 339.800 ;
        RECT 500.400 335.800 504.400 336.000 ;
        RECT 489.200 334.000 490.400 334.600 ;
        RECT 485.400 332.600 489.200 333.400 ;
        RECT 460.200 332.000 461.000 332.200 ;
        RECT 463.600 332.000 464.400 332.400 ;
        RECT 465.200 332.000 466.000 332.400 ;
        RECT 482.800 332.000 483.600 332.600 ;
        RECT 489.800 332.000 490.400 334.000 ;
        RECT 460.200 331.400 483.600 332.000 ;
        RECT 489.600 331.400 490.400 332.000 ;
        RECT 489.600 329.600 490.200 331.400 ;
        RECT 491.000 330.800 491.800 335.200 ;
        RECT 468.400 329.400 469.200 329.600 ;
        RECT 463.800 329.000 469.200 329.400 ;
        RECT 463.000 328.800 469.200 329.000 ;
        RECT 470.200 329.000 478.800 329.600 ;
        RECT 460.400 328.000 462.000 328.800 ;
        RECT 463.000 328.200 464.400 328.800 ;
        RECT 470.200 328.200 470.800 329.000 ;
        RECT 478.000 328.800 478.800 329.000 ;
        RECT 481.200 329.000 490.200 329.600 ;
        RECT 481.200 328.800 482.000 329.000 ;
        RECT 461.400 327.600 462.000 328.000 ;
        RECT 465.000 327.600 470.800 328.200 ;
        RECT 471.400 327.600 474.000 328.400 ;
        RECT 458.800 326.800 460.800 327.400 ;
        RECT 461.400 326.800 465.600 327.600 ;
        RECT 460.200 326.200 460.800 326.800 ;
        RECT 460.200 325.600 461.200 326.200 ;
        RECT 460.400 322.200 461.200 325.600 ;
        RECT 463.600 322.200 464.400 326.800 ;
        RECT 466.800 322.200 467.600 325.000 ;
        RECT 468.400 322.200 469.200 325.000 ;
        RECT 470.000 322.200 470.800 327.000 ;
        RECT 473.200 322.200 474.000 327.000 ;
        RECT 476.400 322.200 477.200 328.400 ;
        RECT 484.400 327.600 487.000 328.400 ;
        RECT 479.600 326.800 483.800 327.600 ;
        RECT 478.000 322.200 478.800 325.000 ;
        RECT 479.600 322.200 480.400 325.000 ;
        RECT 481.200 322.200 482.000 325.000 ;
        RECT 484.400 322.200 485.200 327.600 ;
        RECT 489.600 327.400 490.200 329.000 ;
        RECT 487.600 326.800 490.200 327.400 ;
        RECT 490.800 330.000 491.800 330.800 ;
        RECT 495.600 332.300 496.400 335.800 ;
        RECT 497.200 334.300 498.000 335.200 ;
        RECT 499.000 334.400 499.600 335.800 ;
        RECT 500.600 335.400 504.200 335.800 ;
        RECT 502.800 334.400 503.600 334.800 ;
        RECT 498.800 334.300 501.400 334.400 ;
        RECT 497.200 333.700 501.400 334.300 ;
        RECT 502.800 333.800 504.400 334.400 ;
        RECT 497.200 333.600 498.000 333.700 ;
        RECT 498.800 333.600 501.400 333.700 ;
        RECT 503.600 333.600 504.400 333.800 ;
        RECT 497.200 332.300 498.000 332.400 ;
        RECT 495.600 331.700 498.000 332.300 ;
        RECT 487.600 322.200 488.400 326.800 ;
        RECT 490.800 322.200 491.600 330.000 ;
        RECT 494.000 328.800 494.800 330.400 ;
        RECT 495.600 322.200 496.400 331.700 ;
        RECT 497.200 331.600 498.000 331.700 ;
        RECT 497.200 330.300 498.000 330.400 ;
        RECT 498.800 330.300 499.600 330.400 ;
        RECT 497.200 330.200 499.600 330.300 ;
        RECT 500.800 330.200 501.400 333.600 ;
        RECT 502.000 331.600 502.800 333.200 ;
        RECT 497.200 329.700 500.200 330.200 ;
        RECT 497.200 329.600 498.000 329.700 ;
        RECT 498.800 329.600 500.200 329.700 ;
        RECT 500.800 329.600 501.800 330.200 ;
        RECT 499.600 328.400 500.200 329.600 ;
        RECT 499.600 327.600 500.400 328.400 ;
        RECT 501.000 322.200 501.800 329.600 ;
        RECT 505.200 322.200 506.000 339.800 ;
        RECT 506.800 335.600 507.600 337.200 ;
        RECT 508.400 336.000 509.200 339.800 ;
        RECT 511.600 336.000 512.400 339.800 ;
        RECT 508.400 335.800 512.400 336.000 ;
        RECT 513.200 335.800 514.000 339.800 ;
        RECT 514.800 336.000 515.600 339.800 ;
        RECT 518.000 336.000 518.800 339.800 ;
        RECT 514.800 335.800 518.800 336.000 ;
        RECT 519.600 336.300 520.400 339.800 ;
        RECT 522.800 337.600 523.600 339.800 ;
        RECT 521.200 336.300 522.000 336.400 ;
        RECT 508.600 335.400 512.200 335.800 ;
        RECT 509.200 334.400 510.000 334.800 ;
        RECT 513.200 334.400 513.800 335.800 ;
        RECT 515.000 335.400 518.600 335.800 ;
        RECT 519.600 335.700 522.000 336.300 ;
        RECT 515.600 334.400 516.400 334.800 ;
        RECT 519.600 334.400 520.200 335.700 ;
        RECT 521.200 335.600 522.000 335.700 ;
        RECT 522.800 334.400 523.400 337.600 ;
        RECT 524.400 336.300 525.200 337.200 ;
        RECT 526.000 336.300 526.800 337.200 ;
        RECT 524.400 335.700 526.800 336.300 ;
        RECT 524.400 335.600 525.200 335.700 ;
        RECT 526.000 335.600 526.800 335.700 ;
        RECT 508.400 333.800 510.000 334.400 ;
        RECT 508.400 333.600 509.200 333.800 ;
        RECT 511.400 333.600 514.000 334.400 ;
        RECT 514.800 333.800 516.400 334.400 ;
        RECT 514.800 333.600 515.600 333.800 ;
        RECT 517.800 333.600 520.400 334.400 ;
        RECT 522.800 333.600 523.600 334.400 ;
        RECT 527.600 334.300 528.400 339.800 ;
        RECT 529.200 336.000 530.000 339.800 ;
        RECT 532.400 336.000 533.200 339.800 ;
        RECT 529.200 335.800 533.200 336.000 ;
        RECT 534.000 335.800 534.800 339.800 ;
        RECT 535.600 336.000 536.400 339.800 ;
        RECT 538.800 336.000 539.600 339.800 ;
        RECT 535.600 335.800 539.600 336.000 ;
        RECT 540.400 335.800 541.200 339.800 ;
        RECT 529.400 335.400 533.000 335.800 ;
        RECT 530.000 334.400 530.800 334.800 ;
        RECT 534.000 334.400 534.600 335.800 ;
        RECT 535.800 335.400 539.400 335.800 ;
        RECT 536.400 334.400 537.200 334.800 ;
        RECT 540.400 334.400 541.000 335.800 ;
        RECT 529.200 334.300 530.800 334.400 ;
        RECT 527.600 333.800 530.800 334.300 ;
        RECT 527.600 333.700 530.000 333.800 ;
        RECT 510.000 331.600 510.800 333.200 ;
        RECT 511.400 332.300 512.000 333.600 ;
        RECT 514.800 332.300 515.600 332.400 ;
        RECT 511.400 331.700 515.600 332.300 ;
        RECT 511.400 330.200 512.000 331.700 ;
        RECT 514.800 331.600 515.600 331.700 ;
        RECT 516.400 331.600 517.200 333.200 ;
        RECT 517.800 332.400 518.400 333.600 ;
        RECT 517.800 331.600 518.800 332.400 ;
        RECT 513.200 330.200 514.000 330.400 ;
        RECT 517.800 330.200 518.400 331.600 ;
        RECT 521.200 330.800 522.000 332.400 ;
        RECT 519.600 330.200 520.400 330.400 ;
        RECT 522.800 330.200 523.400 333.600 ;
        RECT 511.000 329.600 512.000 330.200 ;
        RECT 512.600 329.600 514.000 330.200 ;
        RECT 517.400 329.600 518.400 330.200 ;
        RECT 519.000 329.600 520.400 330.200 ;
        RECT 511.000 322.200 511.800 329.600 ;
        RECT 512.600 328.400 513.200 329.600 ;
        RECT 512.400 327.600 513.200 328.400 ;
        RECT 517.400 322.200 518.200 329.600 ;
        RECT 519.000 328.400 519.600 329.600 ;
        RECT 518.800 327.600 519.600 328.400 ;
        RECT 521.800 329.400 523.600 330.200 ;
        RECT 521.800 322.200 522.600 329.400 ;
        RECT 527.600 322.200 528.400 333.700 ;
        RECT 529.200 333.600 530.000 333.700 ;
        RECT 532.200 333.600 534.800 334.400 ;
        RECT 535.600 333.800 537.200 334.400 ;
        RECT 535.600 333.600 536.400 333.800 ;
        RECT 538.600 333.600 541.200 334.400 ;
        RECT 530.800 331.600 531.600 333.200 ;
        RECT 532.200 330.200 532.800 333.600 ;
        RECT 537.200 331.600 538.000 333.200 ;
        RECT 538.600 330.400 539.200 333.600 ;
        RECT 534.000 330.200 534.800 330.400 ;
        RECT 531.800 329.600 532.800 330.200 ;
        RECT 533.400 329.600 534.800 330.200 ;
        RECT 537.200 329.600 539.200 330.400 ;
        RECT 540.400 330.300 541.200 330.400 ;
        RECT 542.000 330.300 542.800 339.800 ;
        RECT 543.600 335.600 544.400 337.200 ;
        RECT 548.400 335.200 549.200 339.800 ;
        RECT 547.000 334.600 549.200 335.200 ;
        RECT 547.000 331.600 547.600 334.600 ;
        RECT 548.400 331.600 549.200 333.200 ;
        RECT 546.400 330.800 547.600 331.600 ;
        RECT 540.400 330.200 542.800 330.300 ;
        RECT 539.800 329.700 542.800 330.200 ;
        RECT 539.800 329.600 541.200 329.700 ;
        RECT 531.800 322.200 532.600 329.600 ;
        RECT 533.400 328.400 534.000 329.600 ;
        RECT 533.200 327.600 534.000 328.400 ;
        RECT 538.200 322.200 539.000 329.600 ;
        RECT 539.800 328.400 540.400 329.600 ;
        RECT 539.600 327.600 541.200 328.400 ;
        RECT 542.000 322.200 542.800 329.700 ;
        RECT 547.000 330.200 547.600 330.800 ;
        RECT 547.000 329.600 549.200 330.200 ;
        RECT 548.400 322.200 549.200 329.600 ;
        RECT 1.800 312.600 2.600 319.800 ;
        RECT 7.600 315.800 8.400 319.800 ;
        RECT 7.800 315.600 8.400 315.800 ;
        RECT 10.800 315.800 11.600 319.800 ;
        RECT 10.800 315.600 11.400 315.800 ;
        RECT 7.800 315.000 11.400 315.600 ;
        RECT 9.200 312.800 10.000 314.400 ;
        RECT 1.800 311.800 3.600 312.600 ;
        RECT 10.800 312.400 11.400 315.000 ;
        RECT 1.200 309.600 2.000 311.200 ;
        RECT 2.800 308.400 3.400 311.800 ;
        RECT 6.000 310.800 6.800 312.400 ;
        RECT 10.800 311.600 11.600 312.400 ;
        RECT 7.600 309.600 9.200 310.400 ;
        RECT 10.800 308.400 11.400 311.600 ;
        RECT 2.800 307.600 3.600 308.400 ;
        RECT 9.800 308.200 11.400 308.400 ;
        RECT 9.600 307.800 11.400 308.200 ;
        RECT 1.200 306.300 2.000 306.400 ;
        RECT 2.800 306.300 3.400 307.600 ;
        RECT 1.200 305.700 3.500 306.300 ;
        RECT 1.200 305.600 2.000 305.700 ;
        RECT 2.800 304.200 3.400 305.700 ;
        RECT 4.400 304.800 5.200 306.400 ;
        RECT 9.600 304.400 10.400 307.800 ;
        RECT 2.800 302.200 3.600 304.200 ;
        RECT 9.600 303.600 11.600 304.400 ;
        RECT 9.600 302.200 10.400 303.600 ;
        RECT 12.400 302.200 13.200 319.800 ;
        RECT 15.600 315.800 16.400 319.800 ;
        RECT 15.800 315.600 16.400 315.800 ;
        RECT 18.800 315.800 19.600 319.800 ;
        RECT 18.800 315.600 19.400 315.800 ;
        RECT 15.800 315.000 19.400 315.600 ;
        RECT 15.800 312.400 16.400 315.000 ;
        RECT 17.200 312.800 18.000 314.400 ;
        RECT 15.600 311.600 16.400 312.400 ;
        RECT 15.800 308.400 16.400 311.600 ;
        RECT 20.400 312.300 21.200 312.400 ;
        RECT 22.000 312.300 22.800 312.400 ;
        RECT 20.400 311.700 22.800 312.300 ;
        RECT 20.400 310.800 21.200 311.700 ;
        RECT 22.000 311.600 22.800 311.700 ;
        RECT 18.000 309.600 19.600 310.400 ;
        RECT 15.800 308.200 17.400 308.400 ;
        RECT 15.800 307.800 17.600 308.200 ;
        RECT 14.000 304.800 14.800 306.400 ;
        RECT 16.800 304.300 17.600 307.800 ;
        RECT 22.000 306.800 22.800 308.400 ;
        RECT 23.600 306.200 24.400 319.800 ;
        RECT 29.000 318.400 29.800 319.800 ;
        RECT 29.000 317.600 30.800 318.400 ;
        RECT 27.600 313.600 28.400 314.400 ;
        RECT 25.200 311.600 26.000 313.200 ;
        RECT 27.600 312.400 28.200 313.600 ;
        RECT 29.000 312.400 29.800 317.600 ;
        RECT 35.800 312.600 36.600 319.800 ;
        RECT 40.600 314.400 41.400 319.800 ;
        RECT 45.400 318.400 47.400 319.800 ;
        RECT 44.400 317.600 47.400 318.400 ;
        RECT 40.600 313.600 42.000 314.400 ;
        RECT 40.600 312.600 41.400 313.600 ;
        RECT 26.800 311.800 28.200 312.400 ;
        RECT 28.800 311.800 29.800 312.400 ;
        RECT 34.800 311.800 36.600 312.600 ;
        RECT 39.600 311.800 41.400 312.600 ;
        RECT 45.400 311.800 47.400 317.600 ;
        RECT 26.800 311.600 27.600 311.800 ;
        RECT 28.800 308.400 29.400 311.800 ;
        RECT 30.000 308.800 30.800 310.400 ;
        RECT 35.000 308.400 35.600 311.800 ;
        RECT 36.400 309.600 37.200 311.200 ;
        RECT 39.800 308.400 40.400 311.800 ;
        RECT 41.200 309.600 42.000 311.200 ;
        RECT 44.400 308.800 45.200 310.400 ;
        RECT 46.000 308.400 46.600 311.800 ;
        RECT 47.600 308.800 48.400 310.400 ;
        RECT 26.800 307.600 29.400 308.400 ;
        RECT 31.600 308.200 32.400 308.400 ;
        RECT 30.800 307.600 32.400 308.200 ;
        RECT 34.800 307.600 35.600 308.400 ;
        RECT 39.600 307.600 40.400 308.400 ;
        RECT 42.800 308.200 43.600 308.400 ;
        RECT 46.000 308.200 46.800 308.400 ;
        RECT 42.800 307.600 44.400 308.200 ;
        RECT 46.000 307.600 48.400 308.200 ;
        RECT 49.200 307.600 50.000 309.200 ;
        RECT 27.000 306.200 27.600 307.600 ;
        RECT 30.800 307.200 31.600 307.600 ;
        RECT 28.600 306.200 32.200 306.600 ;
        RECT 35.000 306.400 35.600 307.600 ;
        RECT 23.600 305.600 25.400 306.200 ;
        RECT 18.800 304.300 19.600 304.400 ;
        RECT 16.800 303.700 19.600 304.300 ;
        RECT 16.800 302.200 17.600 303.700 ;
        RECT 18.800 303.600 19.600 303.700 ;
        RECT 24.600 302.200 25.400 305.600 ;
        RECT 26.800 302.200 27.600 306.200 ;
        RECT 28.400 306.000 32.400 306.200 ;
        RECT 28.400 302.200 29.200 306.000 ;
        RECT 31.600 302.200 32.400 306.000 ;
        RECT 33.200 304.800 34.000 306.400 ;
        RECT 34.800 305.600 35.600 306.400 ;
        RECT 35.000 304.200 35.600 305.600 ;
        RECT 38.000 304.800 38.800 306.400 ;
        RECT 39.800 304.200 40.400 307.600 ;
        RECT 43.600 307.200 44.400 307.600 ;
        RECT 43.000 306.200 46.600 306.600 ;
        RECT 47.800 306.200 48.400 307.600 ;
        RECT 50.800 306.800 51.600 308.400 ;
        RECT 52.400 306.200 53.200 319.800 ;
        RECT 57.200 315.800 58.000 319.800 ;
        RECT 57.400 315.600 58.000 315.800 ;
        RECT 60.400 315.800 61.200 319.800 ;
        RECT 60.400 315.600 61.000 315.800 ;
        RECT 57.400 315.000 61.000 315.600 ;
        RECT 58.800 314.300 59.600 314.400 ;
        RECT 54.000 313.700 59.600 314.300 ;
        RECT 54.000 311.600 54.800 313.700 ;
        RECT 58.800 312.800 59.600 313.700 ;
        RECT 60.400 312.400 61.000 315.000 ;
        RECT 55.600 310.800 56.400 312.400 ;
        RECT 60.400 311.600 61.200 312.400 ;
        RECT 57.200 309.600 58.800 310.400 ;
        RECT 60.400 308.400 61.000 311.600 ;
        RECT 59.400 308.200 61.000 308.400 ;
        RECT 59.200 307.800 61.000 308.200 ;
        RECT 34.800 302.200 35.600 304.200 ;
        RECT 39.600 302.200 40.400 304.200 ;
        RECT 42.800 306.000 46.800 306.200 ;
        RECT 42.800 302.200 43.600 306.000 ;
        RECT 46.000 302.800 46.800 306.000 ;
        RECT 47.600 303.400 48.400 306.200 ;
        RECT 49.200 302.800 50.000 306.200 ;
        RECT 52.400 305.600 54.200 306.200 ;
        RECT 46.000 302.200 50.000 302.800 ;
        RECT 53.400 302.200 54.200 305.600 ;
        RECT 57.200 304.300 58.000 304.400 ;
        RECT 59.200 304.300 60.000 307.800 ;
        RECT 62.000 306.800 62.800 308.400 ;
        RECT 63.600 306.200 64.400 319.800 ;
        RECT 69.400 318.400 71.400 319.800 ;
        RECT 68.400 317.600 71.400 318.400 ;
        RECT 65.200 311.600 66.000 313.200 ;
        RECT 69.400 311.800 71.400 317.600 ;
        RECT 66.800 310.300 67.600 310.400 ;
        RECT 68.400 310.300 69.200 310.400 ;
        RECT 66.800 309.700 69.200 310.300 ;
        RECT 66.800 309.600 67.600 309.700 ;
        RECT 68.400 308.800 69.200 309.700 ;
        RECT 70.000 308.400 70.600 311.800 ;
        RECT 71.600 308.800 72.400 310.400 ;
        RECT 66.800 308.200 67.600 308.400 ;
        RECT 70.000 308.200 70.800 308.400 ;
        RECT 66.800 307.600 68.400 308.200 ;
        RECT 70.000 307.600 72.400 308.200 ;
        RECT 73.200 307.600 74.000 309.200 ;
        RECT 67.600 307.200 68.400 307.600 ;
        RECT 67.000 306.200 70.600 306.600 ;
        RECT 71.800 306.200 72.400 307.600 ;
        RECT 63.600 305.600 65.400 306.200 ;
        RECT 57.200 303.700 60.000 304.300 ;
        RECT 57.200 303.600 58.000 303.700 ;
        RECT 59.200 302.200 60.000 303.700 ;
        RECT 64.600 302.200 65.400 305.600 ;
        RECT 66.800 306.000 70.800 306.200 ;
        RECT 66.800 302.200 67.600 306.000 ;
        RECT 70.000 302.800 70.800 306.000 ;
        RECT 71.600 303.400 72.400 306.200 ;
        RECT 73.200 302.800 74.000 306.200 ;
        RECT 74.800 304.800 75.600 306.400 ;
        RECT 70.000 302.200 74.000 302.800 ;
        RECT 76.400 302.200 77.200 319.800 ;
        RECT 79.600 311.200 80.400 319.800 ;
        RECT 82.800 311.200 83.600 319.800 ;
        RECT 86.000 311.200 86.800 319.800 ;
        RECT 89.200 311.200 90.000 319.800 ;
        RECT 95.000 312.400 95.800 319.800 ;
        RECT 96.400 313.600 97.200 314.400 ;
        RECT 96.600 312.400 97.200 313.600 ;
        RECT 94.000 311.600 96.000 312.400 ;
        RECT 96.600 311.800 98.000 312.400 ;
        RECT 97.200 311.600 98.000 311.800 ;
        RECT 98.800 311.600 99.600 313.200 ;
        RECT 79.600 310.400 81.400 311.200 ;
        RECT 82.800 310.400 85.000 311.200 ;
        RECT 86.000 310.400 88.200 311.200 ;
        RECT 89.200 310.400 91.600 311.200 ;
        RECT 80.600 309.000 81.400 310.400 ;
        RECT 84.200 309.000 85.000 310.400 ;
        RECT 87.400 309.000 88.200 310.400 ;
        RECT 80.600 308.200 83.200 309.000 ;
        RECT 84.200 308.200 86.600 309.000 ;
        RECT 87.400 308.200 90.000 309.000 ;
        RECT 80.600 307.600 81.400 308.200 ;
        RECT 84.200 307.600 85.000 308.200 ;
        RECT 87.400 307.600 88.200 308.200 ;
        RECT 90.800 307.600 91.600 310.400 ;
        RECT 92.400 310.300 93.200 310.400 ;
        RECT 94.000 310.300 94.800 310.400 ;
        RECT 92.400 309.700 94.800 310.300 ;
        RECT 92.400 309.600 93.200 309.700 ;
        RECT 94.000 308.800 94.800 309.700 ;
        RECT 95.400 308.400 96.000 311.600 ;
        RECT 97.300 310.300 97.900 311.600 ;
        RECT 100.400 310.300 101.200 319.800 ;
        RECT 97.300 309.700 101.200 310.300 ;
        RECT 92.400 308.200 93.200 308.400 ;
        RECT 92.400 307.600 94.000 308.200 ;
        RECT 95.400 307.600 98.000 308.400 ;
        RECT 79.600 306.800 81.400 307.600 ;
        RECT 82.800 306.800 85.000 307.600 ;
        RECT 86.000 306.800 88.200 307.600 ;
        RECT 89.200 306.800 91.600 307.600 ;
        RECT 93.200 307.200 94.000 307.600 ;
        RECT 79.600 302.200 80.400 306.800 ;
        RECT 82.800 302.200 83.600 306.800 ;
        RECT 86.000 302.200 86.800 306.800 ;
        RECT 89.200 302.200 90.000 306.800 ;
        RECT 92.600 306.200 96.200 306.600 ;
        RECT 97.200 306.200 97.800 307.600 ;
        RECT 100.400 306.200 101.200 309.700 ;
        RECT 102.000 306.800 102.800 308.400 ;
        RECT 103.600 306.800 104.400 308.400 ;
        RECT 92.400 306.000 96.400 306.200 ;
        RECT 92.400 302.200 93.200 306.000 ;
        RECT 95.600 302.200 96.400 306.000 ;
        RECT 97.200 302.200 98.000 306.200 ;
        RECT 99.400 305.600 101.200 306.200 ;
        RECT 99.400 302.200 100.200 305.600 ;
        RECT 105.200 302.200 106.000 319.800 ;
        RECT 108.400 304.800 109.200 306.400 ;
        RECT 110.000 302.200 110.800 319.800 ;
        RECT 113.200 310.300 114.000 319.800 ;
        RECT 117.400 312.600 118.200 319.800 ;
        RECT 121.200 315.800 122.000 319.800 ;
        RECT 116.400 311.800 118.200 312.600 ;
        RECT 114.800 310.300 115.600 310.400 ;
        RECT 113.200 309.700 115.600 310.300 ;
        RECT 111.600 304.800 112.400 306.400 ;
        RECT 113.200 306.300 114.000 309.700 ;
        RECT 114.800 309.600 115.600 309.700 ;
        RECT 116.600 308.400 117.200 311.800 ;
        RECT 121.400 311.600 122.000 315.800 ;
        RECT 124.400 311.800 125.200 319.800 ;
        RECT 132.400 315.800 133.200 319.800 ;
        RECT 132.600 315.600 133.200 315.800 ;
        RECT 135.600 315.800 136.400 319.800 ;
        RECT 141.400 318.400 142.200 319.800 ;
        RECT 140.400 317.600 142.200 318.400 ;
        RECT 135.600 315.600 136.200 315.800 ;
        RECT 132.600 315.000 136.200 315.600 ;
        RECT 132.600 312.400 133.200 315.000 ;
        RECT 134.000 312.800 134.800 314.400 ;
        RECT 141.400 312.400 142.200 317.600 ;
        RECT 142.800 313.600 143.600 314.400 ;
        RECT 143.000 312.400 143.600 313.600 ;
        RECT 118.000 310.300 118.800 311.200 ;
        RECT 121.400 311.000 123.800 311.600 ;
        RECT 118.000 309.700 120.400 310.300 ;
        RECT 118.000 309.600 118.800 309.700 ;
        RECT 116.400 307.600 117.200 308.400 ;
        RECT 119.600 307.600 120.400 309.700 ;
        RECT 121.200 309.600 122.000 310.400 ;
        RECT 121.400 308.800 122.000 309.600 ;
        RECT 121.400 308.200 122.400 308.800 ;
        RECT 121.600 308.000 122.400 308.200 ;
        RECT 123.200 307.600 123.800 311.000 ;
        RECT 124.600 310.400 125.200 311.800 ;
        RECT 132.400 311.600 133.200 312.400 ;
        RECT 124.400 309.600 125.200 310.400 ;
        RECT 114.800 306.300 115.600 306.400 ;
        RECT 116.600 306.300 117.200 307.600 ;
        RECT 123.200 307.400 124.000 307.600 ;
        RECT 121.000 307.000 124.000 307.400 ;
        RECT 119.800 306.800 124.000 307.000 ;
        RECT 119.800 306.400 121.600 306.800 ;
        RECT 118.000 306.300 118.800 306.400 ;
        RECT 113.200 305.700 115.600 306.300 ;
        RECT 116.500 305.700 118.800 306.300 ;
        RECT 119.800 306.200 120.400 306.400 ;
        RECT 124.600 306.200 125.200 309.600 ;
        RECT 132.600 308.400 133.200 311.600 ;
        RECT 134.800 309.600 136.400 310.400 ;
        RECT 137.200 310.300 138.000 312.400 ;
        RECT 141.400 311.800 142.400 312.400 ;
        RECT 143.000 311.800 144.400 312.400 ;
        RECT 137.200 309.700 139.500 310.300 ;
        RECT 138.900 308.400 139.500 309.700 ;
        RECT 140.400 308.800 141.200 310.400 ;
        RECT 141.800 308.400 142.400 311.800 ;
        RECT 143.600 311.600 144.400 311.800 ;
        RECT 146.800 311.200 147.600 319.800 ;
        RECT 150.000 311.200 150.800 319.800 ;
        RECT 153.200 311.200 154.000 319.800 ;
        RECT 156.400 311.200 157.200 319.800 ;
        RECT 159.600 312.400 160.400 319.800 ;
        RECT 162.800 312.400 163.600 319.800 ;
        RECT 159.600 311.800 163.600 312.400 ;
        RECT 164.400 311.800 165.200 319.800 ;
        RECT 166.800 313.600 167.600 314.400 ;
        RECT 166.800 312.400 167.400 313.600 ;
        RECT 168.200 312.400 169.000 319.800 ;
        RECT 173.200 313.600 174.000 314.400 ;
        RECT 173.200 312.400 173.800 313.600 ;
        RECT 174.600 312.400 175.400 319.800 ;
        RECT 166.000 311.800 167.400 312.400 ;
        RECT 168.000 311.800 169.000 312.400 ;
        RECT 172.400 311.800 173.800 312.400 ;
        RECT 174.400 311.800 175.400 312.400 ;
        RECT 146.800 310.400 148.600 311.200 ;
        RECT 150.000 310.400 152.200 311.200 ;
        RECT 153.200 310.400 155.400 311.200 ;
        RECT 156.400 310.400 158.800 311.200 ;
        RECT 160.400 310.400 161.200 310.800 ;
        RECT 164.400 310.400 165.000 311.800 ;
        RECT 166.000 311.600 166.800 311.800 ;
        RECT 168.000 310.400 168.600 311.800 ;
        RECT 172.400 311.600 173.200 311.800 ;
        RECT 147.800 309.000 148.600 310.400 ;
        RECT 151.400 309.000 152.200 310.400 ;
        RECT 154.600 309.000 155.400 310.400 ;
        RECT 132.600 308.200 134.200 308.400 ;
        RECT 138.800 308.200 139.600 308.400 ;
        RECT 132.600 307.800 134.400 308.200 ;
        RECT 113.200 302.200 114.000 305.700 ;
        RECT 114.800 304.800 115.600 305.700 ;
        RECT 116.600 304.200 117.200 305.700 ;
        RECT 118.000 305.600 118.800 305.700 ;
        RECT 116.400 302.200 117.200 304.200 ;
        RECT 119.600 302.200 120.400 306.200 ;
        RECT 123.800 305.200 125.200 306.200 ;
        RECT 123.800 304.300 124.600 305.200 ;
        RECT 126.000 304.300 126.800 304.400 ;
        RECT 123.800 303.700 126.800 304.300 ;
        RECT 123.800 302.200 124.600 303.700 ;
        RECT 126.000 303.600 126.800 303.700 ;
        RECT 133.600 304.300 134.400 307.800 ;
        RECT 138.800 307.600 140.400 308.200 ;
        RECT 141.800 307.600 144.400 308.400 ;
        RECT 147.800 308.200 150.400 309.000 ;
        RECT 151.400 308.200 153.800 309.000 ;
        RECT 154.600 308.200 157.200 309.000 ;
        RECT 147.800 307.600 148.600 308.200 ;
        RECT 151.400 307.600 152.200 308.200 ;
        RECT 154.600 307.600 155.400 308.200 ;
        RECT 158.000 307.600 158.800 310.400 ;
        RECT 159.600 309.800 161.200 310.400 ;
        RECT 162.800 309.800 165.200 310.400 ;
        RECT 159.600 309.600 160.400 309.800 ;
        RECT 161.200 307.600 162.000 309.200 ;
        RECT 139.600 307.200 140.400 307.600 ;
        RECT 139.000 306.200 142.600 306.600 ;
        RECT 143.600 306.200 144.200 307.600 ;
        RECT 146.800 306.800 148.600 307.600 ;
        RECT 150.000 306.800 152.200 307.600 ;
        RECT 153.200 306.800 155.400 307.600 ;
        RECT 156.400 306.800 158.800 307.600 ;
        RECT 138.800 306.000 142.800 306.200 ;
        RECT 135.600 304.300 136.400 304.400 ;
        RECT 133.600 303.700 136.400 304.300 ;
        RECT 133.600 302.200 134.400 303.700 ;
        RECT 135.600 303.600 136.400 303.700 ;
        RECT 138.800 302.200 139.600 306.000 ;
        RECT 142.000 302.200 142.800 306.000 ;
        RECT 143.600 302.200 144.400 306.200 ;
        RECT 146.800 302.200 147.600 306.800 ;
        RECT 150.000 302.200 150.800 306.800 ;
        RECT 153.200 302.200 154.000 306.800 ;
        RECT 156.400 302.200 157.200 306.800 ;
        RECT 162.800 306.200 163.400 309.800 ;
        RECT 164.400 309.600 165.200 309.800 ;
        RECT 167.600 309.600 168.600 310.400 ;
        RECT 168.000 308.400 168.600 309.600 ;
        RECT 169.200 308.800 170.000 310.400 ;
        RECT 170.800 310.300 171.600 310.400 ;
        RECT 174.400 310.300 175.000 311.800 ;
        RECT 170.800 309.700 175.000 310.300 ;
        RECT 170.800 309.600 171.600 309.700 ;
        RECT 174.400 308.400 175.000 309.700 ;
        RECT 175.600 308.800 176.400 310.400 ;
        RECT 166.000 307.600 168.600 308.400 ;
        RECT 170.800 308.200 171.600 308.400 ;
        RECT 170.000 307.600 171.600 308.200 ;
        RECT 172.400 307.600 175.000 308.400 ;
        RECT 177.200 308.300 178.000 308.400 ;
        RECT 180.400 308.300 181.200 319.800 ;
        RECT 182.000 308.300 182.800 308.400 ;
        RECT 177.200 308.200 182.800 308.300 ;
        RECT 176.400 307.700 182.800 308.200 ;
        RECT 176.400 307.600 178.000 307.700 ;
        RECT 162.800 302.200 163.600 306.200 ;
        RECT 164.400 305.600 165.200 306.400 ;
        RECT 166.200 306.200 166.800 307.600 ;
        RECT 170.000 307.200 170.800 307.600 ;
        RECT 167.800 306.200 171.400 306.600 ;
        RECT 172.600 306.200 173.200 307.600 ;
        RECT 176.400 307.200 177.200 307.600 ;
        RECT 174.200 306.200 177.800 306.600 ;
        RECT 164.200 304.800 165.000 305.600 ;
        RECT 166.000 302.200 166.800 306.200 ;
        RECT 167.600 306.000 171.600 306.200 ;
        RECT 167.600 302.200 168.400 306.000 ;
        RECT 170.800 302.200 171.600 306.000 ;
        RECT 172.400 302.200 173.200 306.200 ;
        RECT 174.000 306.000 178.000 306.200 ;
        RECT 174.000 302.200 174.800 306.000 ;
        RECT 177.200 302.200 178.000 306.000 ;
        RECT 178.800 304.800 179.600 306.400 ;
        RECT 180.400 302.200 181.200 307.700 ;
        RECT 182.000 306.800 182.800 307.700 ;
        RECT 183.600 306.200 184.400 319.800 ;
        RECT 185.200 311.600 186.000 313.200 ;
        RECT 189.400 312.600 190.200 319.800 ;
        RECT 193.800 318.400 194.600 319.800 ;
        RECT 193.800 317.600 195.600 318.400 ;
        RECT 188.400 311.800 190.200 312.600 ;
        RECT 192.400 313.600 193.200 314.400 ;
        RECT 192.400 312.400 193.000 313.600 ;
        RECT 193.800 312.400 194.600 317.600 ;
        RECT 191.600 311.800 193.000 312.400 ;
        RECT 193.600 311.800 194.600 312.400 ;
        RECT 185.300 310.300 185.900 311.600 ;
        RECT 188.600 310.300 189.200 311.800 ;
        RECT 191.600 311.600 192.400 311.800 ;
        RECT 185.300 309.700 189.200 310.300 ;
        RECT 188.600 308.400 189.200 309.700 ;
        RECT 190.000 309.600 190.800 311.200 ;
        RECT 193.600 308.400 194.200 311.800 ;
        RECT 194.800 308.800 195.600 310.400 ;
        RECT 188.400 307.600 189.200 308.400 ;
        RECT 191.600 307.600 194.200 308.400 ;
        RECT 196.400 308.300 197.200 308.400 ;
        RECT 198.000 308.300 198.800 319.800 ;
        RECT 196.400 308.200 198.800 308.300 ;
        RECT 195.600 307.700 198.800 308.200 ;
        RECT 195.600 307.600 197.200 307.700 ;
        RECT 183.600 305.600 185.400 306.200 ;
        RECT 184.600 304.400 185.400 305.600 ;
        RECT 186.800 304.800 187.600 306.400 ;
        RECT 183.600 303.600 185.400 304.400 ;
        RECT 188.600 304.200 189.200 307.600 ;
        RECT 191.800 306.200 192.400 307.600 ;
        RECT 195.600 307.200 196.400 307.600 ;
        RECT 193.400 306.200 197.000 306.600 ;
        RECT 184.600 302.200 185.400 303.600 ;
        RECT 188.400 302.200 189.200 304.200 ;
        RECT 191.600 302.200 192.400 306.200 ;
        RECT 193.200 306.000 197.200 306.200 ;
        RECT 193.200 302.200 194.000 306.000 ;
        RECT 196.400 302.200 197.200 306.000 ;
        RECT 198.000 302.200 198.800 307.700 ;
        RECT 199.600 308.300 200.400 308.400 ;
        RECT 201.200 308.300 202.000 308.400 ;
        RECT 199.600 307.700 202.000 308.300 ;
        RECT 199.600 307.600 200.400 307.700 ;
        RECT 201.200 306.800 202.000 307.700 ;
        RECT 199.600 304.800 200.400 306.400 ;
        RECT 202.800 306.200 203.600 319.800 ;
        RECT 206.800 313.600 207.600 314.400 ;
        RECT 204.400 311.600 205.200 313.200 ;
        RECT 206.800 312.400 207.400 313.600 ;
        RECT 208.200 312.400 209.000 319.800 ;
        RECT 206.000 311.800 207.400 312.400 ;
        RECT 208.000 311.800 209.000 312.400 ;
        RECT 215.000 312.400 215.800 319.800 ;
        RECT 216.400 313.600 217.200 314.400 ;
        RECT 216.600 312.400 217.200 313.600 ;
        RECT 215.000 311.800 216.000 312.400 ;
        RECT 216.600 311.800 218.000 312.400 ;
        RECT 206.000 311.600 206.800 311.800 ;
        RECT 204.500 310.300 205.100 311.600 ;
        RECT 208.000 310.300 208.600 311.800 ;
        RECT 204.500 309.700 208.600 310.300 ;
        RECT 208.000 308.400 208.600 309.700 ;
        RECT 209.200 308.800 210.000 310.400 ;
        RECT 214.000 308.800 214.800 310.400 ;
        RECT 215.400 308.400 216.000 311.800 ;
        RECT 217.200 311.600 218.000 311.800 ;
        RECT 218.800 311.600 219.600 313.200 ;
        RECT 206.000 307.600 208.600 308.400 ;
        RECT 210.800 308.200 211.600 308.400 ;
        RECT 210.000 307.600 211.600 308.200 ;
        RECT 212.400 308.200 213.200 308.400 ;
        RECT 212.400 307.600 214.000 308.200 ;
        RECT 215.400 307.600 218.000 308.400 ;
        RECT 206.200 306.200 206.800 307.600 ;
        RECT 210.000 307.200 210.800 307.600 ;
        RECT 213.200 307.200 214.000 307.600 ;
        RECT 207.800 306.200 211.400 306.600 ;
        RECT 212.600 306.200 216.200 306.600 ;
        RECT 217.200 306.200 217.800 307.600 ;
        RECT 220.400 306.200 221.200 319.800 ;
        RECT 222.000 312.300 222.800 312.400 ;
        RECT 223.600 312.300 224.400 313.200 ;
        RECT 222.000 311.700 224.400 312.300 ;
        RECT 222.000 311.600 222.800 311.700 ;
        RECT 223.600 311.600 224.400 311.700 ;
        RECT 222.000 308.300 222.800 308.400 ;
        RECT 225.200 308.300 226.000 319.800 ;
        RECT 228.400 311.600 229.200 313.200 ;
        RECT 222.000 307.700 226.000 308.300 ;
        RECT 222.000 306.800 222.800 307.700 ;
        RECT 225.200 306.200 226.000 307.700 ;
        RECT 226.800 306.800 227.600 308.400 ;
        RECT 230.000 306.200 230.800 319.800 ;
        RECT 234.000 313.600 234.800 314.400 ;
        RECT 234.000 312.400 234.600 313.600 ;
        RECT 235.400 312.400 236.200 319.800 ;
        RECT 233.200 311.800 234.600 312.400 ;
        RECT 235.200 311.800 236.200 312.400 ;
        RECT 233.200 311.600 234.000 311.800 ;
        RECT 235.200 308.400 235.800 311.800 ;
        RECT 236.400 308.800 237.200 310.400 ;
        RECT 231.600 308.300 232.400 308.400 ;
        RECT 233.200 308.300 235.800 308.400 ;
        RECT 231.600 307.700 235.800 308.300 ;
        RECT 238.000 308.300 238.800 308.400 ;
        RECT 241.200 308.300 242.000 319.800 ;
        RECT 245.400 318.400 246.200 319.800 ;
        RECT 244.400 317.600 246.200 318.400 ;
        RECT 245.400 312.400 246.200 317.600 ;
        RECT 246.800 313.600 247.600 314.400 ;
        RECT 247.000 312.400 247.600 313.600 ;
        RECT 245.400 311.800 246.400 312.400 ;
        RECT 247.000 311.800 248.400 312.400 ;
        RECT 250.800 312.000 251.600 319.800 ;
        RECT 254.000 315.200 254.800 319.800 ;
        RECT 244.400 308.800 245.200 310.400 ;
        RECT 245.800 308.400 246.400 311.800 ;
        RECT 247.600 311.600 248.400 311.800 ;
        RECT 250.600 311.200 251.600 312.000 ;
        RECT 252.200 314.600 254.800 315.200 ;
        RECT 252.200 313.000 252.800 314.600 ;
        RECT 257.200 314.400 258.000 319.800 ;
        RECT 260.400 317.000 261.200 319.800 ;
        RECT 262.000 317.000 262.800 319.800 ;
        RECT 263.600 317.000 264.400 319.800 ;
        RECT 258.600 314.400 262.800 315.200 ;
        RECT 255.400 313.600 258.000 314.400 ;
        RECT 265.200 313.600 266.000 319.800 ;
        RECT 268.400 315.000 269.200 319.800 ;
        RECT 271.600 315.000 272.400 319.800 ;
        RECT 273.200 317.000 274.000 319.800 ;
        RECT 274.800 317.000 275.600 319.800 ;
        RECT 278.000 315.200 278.800 319.800 ;
        RECT 281.200 316.400 282.000 319.800 ;
        RECT 281.200 315.800 282.200 316.400 ;
        RECT 281.600 315.200 282.200 315.800 ;
        RECT 276.800 314.400 281.000 315.200 ;
        RECT 281.600 314.600 283.600 315.200 ;
        RECT 268.400 313.600 271.000 314.400 ;
        RECT 271.600 313.800 277.400 314.400 ;
        RECT 280.400 314.000 281.000 314.400 ;
        RECT 260.400 313.000 261.200 313.200 ;
        RECT 252.200 312.400 261.200 313.000 ;
        RECT 263.600 313.000 264.400 313.200 ;
        RECT 271.600 313.000 272.200 313.800 ;
        RECT 278.000 313.200 279.400 313.800 ;
        RECT 280.400 313.200 282.000 314.000 ;
        RECT 263.600 312.400 272.200 313.000 ;
        RECT 273.200 313.000 279.400 313.200 ;
        RECT 273.200 312.600 278.600 313.000 ;
        RECT 273.200 312.400 274.000 312.600 ;
        RECT 242.800 308.300 243.600 308.400 ;
        RECT 238.000 308.200 240.300 308.300 ;
        RECT 231.600 306.800 232.400 307.700 ;
        RECT 233.200 307.600 235.800 307.700 ;
        RECT 237.200 307.700 240.300 308.200 ;
        RECT 237.200 307.600 238.800 307.700 ;
        RECT 233.400 306.200 234.000 307.600 ;
        RECT 237.200 307.200 238.000 307.600 ;
        RECT 235.000 306.200 238.600 306.600 ;
        RECT 239.700 306.400 240.300 307.700 ;
        RECT 241.200 308.200 243.600 308.300 ;
        RECT 241.200 307.700 244.400 308.200 ;
        RECT 202.800 305.600 204.600 306.200 ;
        RECT 203.800 304.400 204.600 305.600 ;
        RECT 202.800 303.600 204.600 304.400 ;
        RECT 203.800 302.200 204.600 303.600 ;
        RECT 206.000 302.200 206.800 306.200 ;
        RECT 207.600 306.000 211.600 306.200 ;
        RECT 207.600 302.200 208.400 306.000 ;
        RECT 210.800 302.200 211.600 306.000 ;
        RECT 212.400 306.000 216.400 306.200 ;
        RECT 212.400 302.200 213.200 306.000 ;
        RECT 215.600 302.200 216.400 306.000 ;
        RECT 217.200 302.200 218.000 306.200 ;
        RECT 219.400 305.600 221.200 306.200 ;
        RECT 224.200 305.600 226.000 306.200 ;
        RECT 229.000 305.600 230.800 306.200 ;
        RECT 219.400 304.400 220.200 305.600 ;
        RECT 218.800 303.600 220.200 304.400 ;
        RECT 219.400 302.200 220.200 303.600 ;
        RECT 224.200 302.200 225.000 305.600 ;
        RECT 229.000 304.400 229.800 305.600 ;
        RECT 228.400 303.600 229.800 304.400 ;
        RECT 229.000 302.200 229.800 303.600 ;
        RECT 233.200 302.200 234.000 306.200 ;
        RECT 234.800 306.000 238.800 306.200 ;
        RECT 234.800 302.200 235.600 306.000 ;
        RECT 238.000 302.200 238.800 306.000 ;
        RECT 239.600 304.800 240.400 306.400 ;
        RECT 241.200 302.200 242.000 307.700 ;
        RECT 242.800 307.600 244.400 307.700 ;
        RECT 245.800 307.600 248.400 308.400 ;
        RECT 243.600 307.200 244.400 307.600 ;
        RECT 243.000 306.200 246.600 306.600 ;
        RECT 247.600 306.200 248.200 307.600 ;
        RECT 250.600 306.800 251.400 311.200 ;
        RECT 252.200 310.600 252.800 312.400 ;
        RECT 252.000 310.000 252.800 310.600 ;
        RECT 258.800 310.000 282.200 310.600 ;
        RECT 252.000 308.000 252.600 310.000 ;
        RECT 258.800 309.400 259.600 310.000 ;
        RECT 270.000 309.600 270.800 310.000 ;
        RECT 276.400 309.600 277.200 310.000 ;
        RECT 281.200 309.800 282.200 310.000 ;
        RECT 281.200 309.600 282.000 309.800 ;
        RECT 253.200 308.600 257.000 309.400 ;
        RECT 252.000 307.400 253.200 308.000 ;
        RECT 242.800 306.000 246.800 306.200 ;
        RECT 242.800 302.200 243.600 306.000 ;
        RECT 246.000 302.200 246.800 306.000 ;
        RECT 247.600 302.200 248.400 306.200 ;
        RECT 250.600 306.000 251.600 306.800 ;
        RECT 250.800 302.200 251.600 306.000 ;
        RECT 252.400 302.200 253.200 307.400 ;
        RECT 256.200 307.400 257.000 308.600 ;
        RECT 256.200 306.800 258.000 307.400 ;
        RECT 257.200 306.200 258.000 306.800 ;
        RECT 262.000 306.400 262.800 309.200 ;
        RECT 265.200 308.600 268.400 309.400 ;
        RECT 272.200 308.600 274.200 309.400 ;
        RECT 282.800 309.000 283.600 314.600 ;
        RECT 292.400 312.000 293.200 319.800 ;
        RECT 295.600 315.200 296.400 319.800 ;
        RECT 264.800 307.800 265.600 308.000 ;
        RECT 264.800 307.200 269.200 307.800 ;
        RECT 268.400 307.000 269.200 307.200 ;
        RECT 270.000 306.800 270.800 308.400 ;
        RECT 257.200 305.400 259.600 306.200 ;
        RECT 262.000 305.600 263.000 306.400 ;
        RECT 266.000 305.600 267.600 306.400 ;
        RECT 268.400 306.200 269.200 306.400 ;
        RECT 272.200 306.200 273.000 308.600 ;
        RECT 274.800 308.200 283.600 309.000 ;
        RECT 278.200 306.800 281.200 307.600 ;
        RECT 278.200 306.200 279.000 306.800 ;
        RECT 268.400 305.600 273.000 306.200 ;
        RECT 258.800 302.200 259.600 305.400 ;
        RECT 276.400 305.400 279.000 306.200 ;
        RECT 260.400 302.200 261.200 305.000 ;
        RECT 262.000 302.200 262.800 305.000 ;
        RECT 263.600 302.200 264.400 305.000 ;
        RECT 265.200 302.200 266.000 305.000 ;
        RECT 268.400 302.200 269.200 305.000 ;
        RECT 271.600 302.200 272.400 305.000 ;
        RECT 273.200 302.200 274.000 305.000 ;
        RECT 274.800 302.200 275.600 305.000 ;
        RECT 276.400 302.200 277.200 305.400 ;
        RECT 282.800 302.200 283.600 308.200 ;
        RECT 292.200 311.200 293.200 312.000 ;
        RECT 293.800 314.600 296.400 315.200 ;
        RECT 293.800 313.000 294.400 314.600 ;
        RECT 298.800 314.400 299.600 319.800 ;
        RECT 302.000 317.000 302.800 319.800 ;
        RECT 303.600 317.000 304.400 319.800 ;
        RECT 305.200 317.000 306.000 319.800 ;
        RECT 300.200 314.400 304.400 315.200 ;
        RECT 297.000 313.600 299.600 314.400 ;
        RECT 306.800 313.600 307.600 319.800 ;
        RECT 310.000 315.000 310.800 319.800 ;
        RECT 313.200 315.000 314.000 319.800 ;
        RECT 314.800 317.000 315.600 319.800 ;
        RECT 316.400 317.000 317.200 319.800 ;
        RECT 319.600 315.200 320.400 319.800 ;
        RECT 322.800 316.400 323.600 319.800 ;
        RECT 322.800 315.800 323.800 316.400 ;
        RECT 323.200 315.200 323.800 315.800 ;
        RECT 318.400 314.400 322.600 315.200 ;
        RECT 323.200 314.600 325.200 315.200 ;
        RECT 310.000 313.600 312.600 314.400 ;
        RECT 313.200 313.800 319.000 314.400 ;
        RECT 322.000 314.000 322.600 314.400 ;
        RECT 302.000 313.000 302.800 313.200 ;
        RECT 293.800 312.400 302.800 313.000 ;
        RECT 305.200 313.000 306.000 313.200 ;
        RECT 313.200 313.000 313.800 313.800 ;
        RECT 319.600 313.200 321.000 313.800 ;
        RECT 322.000 313.200 323.600 314.000 ;
        RECT 305.200 312.400 313.800 313.000 ;
        RECT 314.800 313.000 321.000 313.200 ;
        RECT 314.800 312.600 320.200 313.000 ;
        RECT 314.800 312.400 315.600 312.600 ;
        RECT 292.200 306.800 293.000 311.200 ;
        RECT 293.800 310.600 294.400 312.400 ;
        RECT 317.800 311.800 318.800 312.000 ;
        RECT 321.200 311.800 322.000 312.400 ;
        RECT 295.000 311.200 322.000 311.800 ;
        RECT 295.000 311.000 295.800 311.200 ;
        RECT 293.600 310.000 294.400 310.600 ;
        RECT 293.600 308.000 294.200 310.000 ;
        RECT 294.800 308.600 298.600 309.400 ;
        RECT 293.600 307.400 294.800 308.000 ;
        RECT 292.200 306.000 293.200 306.800 ;
        RECT 292.400 302.200 293.200 306.000 ;
        RECT 294.000 302.200 294.800 307.400 ;
        RECT 297.800 307.400 298.600 308.600 ;
        RECT 297.800 306.800 299.600 307.400 ;
        RECT 298.800 306.200 299.600 306.800 ;
        RECT 303.600 306.400 304.400 309.200 ;
        RECT 306.800 308.600 310.000 309.400 ;
        RECT 313.800 308.600 315.800 309.400 ;
        RECT 324.400 309.000 325.200 314.600 ;
        RECT 326.000 312.400 326.800 319.800 ;
        RECT 329.200 312.400 330.000 319.800 ;
        RECT 326.000 311.800 330.000 312.400 ;
        RECT 330.800 311.800 331.600 319.800 ;
        RECT 334.600 314.400 335.400 319.800 ;
        RECT 332.400 313.600 334.000 314.400 ;
        RECT 334.600 313.600 336.400 314.400 ;
        RECT 333.200 312.400 333.800 313.600 ;
        RECT 334.600 312.400 335.400 313.600 ;
        RECT 332.400 311.800 333.800 312.400 ;
        RECT 334.400 311.800 335.400 312.400 ;
        RECT 326.800 310.400 327.600 310.800 ;
        RECT 330.800 310.400 331.400 311.800 ;
        RECT 332.400 311.600 333.200 311.800 ;
        RECT 326.000 309.800 327.600 310.400 ;
        RECT 329.200 309.800 331.600 310.400 ;
        RECT 326.000 309.600 326.800 309.800 ;
        RECT 306.400 307.800 307.200 308.000 ;
        RECT 306.400 307.200 310.800 307.800 ;
        RECT 310.000 307.000 310.800 307.200 ;
        RECT 311.600 306.800 312.400 308.400 ;
        RECT 298.800 305.400 301.200 306.200 ;
        RECT 303.600 305.600 304.600 306.400 ;
        RECT 307.600 305.600 309.200 306.400 ;
        RECT 310.000 306.200 310.800 306.400 ;
        RECT 313.800 306.200 314.600 308.600 ;
        RECT 316.400 308.200 325.200 309.000 ;
        RECT 319.800 306.800 322.800 307.600 ;
        RECT 319.800 306.200 320.600 306.800 ;
        RECT 310.000 305.600 314.600 306.200 ;
        RECT 300.400 302.200 301.200 305.400 ;
        RECT 318.000 305.400 320.600 306.200 ;
        RECT 302.000 302.200 302.800 305.000 ;
        RECT 303.600 302.200 304.400 305.000 ;
        RECT 305.200 302.200 306.000 305.000 ;
        RECT 306.800 302.200 307.600 305.000 ;
        RECT 310.000 302.200 310.800 305.000 ;
        RECT 313.200 302.200 314.000 305.000 ;
        RECT 314.800 302.200 315.600 305.000 ;
        RECT 316.400 302.200 317.200 305.000 ;
        RECT 318.000 302.200 318.800 305.400 ;
        RECT 324.400 302.200 325.200 308.200 ;
        RECT 327.600 307.600 328.400 309.200 ;
        RECT 329.200 306.200 329.800 309.800 ;
        RECT 330.800 309.600 331.600 309.800 ;
        RECT 334.400 308.400 335.000 311.800 ;
        RECT 335.600 308.800 336.400 310.400 ;
        RECT 332.400 307.600 335.000 308.400 ;
        RECT 337.200 308.200 338.000 308.400 ;
        RECT 336.400 307.600 338.000 308.200 ;
        RECT 338.800 308.300 339.600 319.800 ;
        RECT 345.200 312.400 346.000 319.800 ;
        RECT 349.400 312.400 350.200 319.800 ;
        RECT 350.800 313.600 351.600 314.400 ;
        RECT 351.000 312.400 351.600 313.600 ;
        RECT 343.800 311.800 346.000 312.400 ;
        RECT 343.800 311.200 344.400 311.800 ;
        RECT 348.400 311.600 350.400 312.400 ;
        RECT 351.000 311.800 352.400 312.400 ;
        RECT 351.600 311.600 352.400 311.800 ;
        RECT 353.200 311.600 354.000 313.200 ;
        RECT 343.200 310.400 344.400 311.200 ;
        RECT 340.400 308.300 341.200 308.400 ;
        RECT 338.800 307.700 341.200 308.300 ;
        RECT 329.200 302.200 330.000 306.200 ;
        RECT 330.800 305.600 331.600 306.400 ;
        RECT 332.600 306.200 333.200 307.600 ;
        RECT 336.400 307.200 337.200 307.600 ;
        RECT 334.200 306.200 337.800 306.600 ;
        RECT 330.600 304.800 331.400 305.600 ;
        RECT 332.400 302.200 333.200 306.200 ;
        RECT 334.000 306.000 338.000 306.200 ;
        RECT 334.000 302.200 334.800 306.000 ;
        RECT 337.200 302.200 338.000 306.000 ;
        RECT 338.800 302.200 339.600 307.700 ;
        RECT 340.400 307.600 341.200 307.700 ;
        RECT 343.800 307.400 344.400 310.400 ;
        RECT 345.200 308.800 346.000 310.400 ;
        RECT 348.400 308.800 349.200 310.400 ;
        RECT 349.800 308.400 350.400 311.600 ;
        RECT 351.700 310.300 352.300 311.600 ;
        RECT 354.800 310.300 355.600 319.800 ;
        RECT 359.600 315.800 360.400 319.800 ;
        RECT 359.800 315.600 360.400 315.800 ;
        RECT 362.800 315.800 363.600 319.800 ;
        RECT 362.800 315.600 363.400 315.800 ;
        RECT 359.800 315.000 363.400 315.600 ;
        RECT 361.200 312.800 362.000 314.400 ;
        RECT 362.800 312.400 363.400 315.000 ;
        RECT 358.000 310.800 358.800 312.400 ;
        RECT 362.800 311.600 363.600 312.400 ;
        RECT 351.700 309.700 355.600 310.300 ;
        RECT 346.800 308.200 347.600 308.400 ;
        RECT 346.800 307.600 348.400 308.200 ;
        RECT 349.800 307.600 352.400 308.400 ;
        RECT 343.800 306.800 346.000 307.400 ;
        RECT 347.600 307.200 348.400 307.600 ;
        RECT 340.400 304.800 341.200 306.400 ;
        RECT 345.200 302.200 346.000 306.800 ;
        RECT 347.000 306.200 350.600 306.600 ;
        RECT 351.600 306.200 352.200 307.600 ;
        RECT 354.800 306.200 355.600 309.700 ;
        RECT 359.600 309.600 361.200 310.400 ;
        RECT 362.800 308.400 363.400 311.600 ;
        RECT 356.400 306.800 357.200 308.400 ;
        RECT 361.800 308.200 363.400 308.400 ;
        RECT 361.600 307.800 363.400 308.200 ;
        RECT 366.000 310.300 366.800 319.800 ;
        RECT 367.600 319.200 371.600 319.800 ;
        RECT 367.600 311.800 368.400 319.200 ;
        RECT 369.200 311.800 370.000 318.600 ;
        RECT 370.800 312.400 371.600 319.200 ;
        RECT 374.000 312.400 374.800 319.800 ;
        RECT 370.800 311.800 374.800 312.400 ;
        RECT 369.400 311.200 370.000 311.800 ;
        RECT 375.600 311.600 376.400 313.200 ;
        RECT 367.600 310.300 368.400 311.200 ;
        RECT 369.400 310.600 371.400 311.200 ;
        RECT 366.000 309.700 368.400 310.300 ;
        RECT 346.800 306.000 350.800 306.200 ;
        RECT 346.800 302.200 347.600 306.000 ;
        RECT 350.000 302.200 350.800 306.000 ;
        RECT 351.600 302.200 352.400 306.200 ;
        RECT 353.800 305.600 355.600 306.200 ;
        RECT 353.800 302.200 354.600 305.600 ;
        RECT 361.600 302.200 362.400 307.800 ;
        RECT 364.400 304.800 365.200 306.400 ;
        RECT 366.000 302.200 366.800 309.700 ;
        RECT 367.600 309.600 368.400 309.700 ;
        RECT 370.800 310.400 371.400 310.600 ;
        RECT 373.200 310.400 374.000 310.800 ;
        RECT 370.800 309.600 371.600 310.400 ;
        RECT 373.200 310.300 374.800 310.400 ;
        RECT 375.600 310.300 376.400 310.400 ;
        RECT 373.200 309.800 376.400 310.300 ;
        RECT 374.000 309.700 376.400 309.800 ;
        RECT 374.000 309.600 374.800 309.700 ;
        RECT 375.600 309.600 376.400 309.700 ;
        RECT 369.400 308.800 370.200 309.600 ;
        RECT 369.400 308.400 370.000 308.800 ;
        RECT 369.200 307.600 370.000 308.400 ;
        RECT 370.800 306.200 371.400 309.600 ;
        RECT 372.400 307.600 373.200 309.200 ;
        RECT 377.200 306.400 378.000 319.800 ;
        RECT 380.400 312.400 381.200 319.800 ;
        RECT 383.600 319.200 387.600 319.800 ;
        RECT 383.600 312.400 384.400 319.200 ;
        RECT 380.400 311.800 384.400 312.400 ;
        RECT 385.200 311.800 386.000 318.600 ;
        RECT 386.800 311.800 387.600 319.200 ;
        RECT 388.400 312.300 389.200 319.800 ;
        RECT 392.400 313.600 393.200 314.400 ;
        RECT 392.400 312.400 393.000 313.600 ;
        RECT 393.800 312.400 394.600 319.800 ;
        RECT 399.600 315.800 400.400 319.800 ;
        RECT 399.800 315.600 400.400 315.800 ;
        RECT 402.800 315.800 403.600 319.800 ;
        RECT 404.400 315.800 405.200 319.800 ;
        RECT 402.800 315.600 403.400 315.800 ;
        RECT 399.800 315.000 403.400 315.600 ;
        RECT 401.200 312.800 402.000 314.400 ;
        RECT 402.800 312.400 403.400 315.000 ;
        RECT 404.600 315.600 405.200 315.800 ;
        RECT 407.600 315.800 408.400 319.800 ;
        RECT 407.600 315.600 408.200 315.800 ;
        RECT 404.600 315.000 408.200 315.600 ;
        RECT 404.600 312.400 405.200 315.000 ;
        RECT 406.000 312.800 406.800 314.400 ;
        RECT 407.600 314.300 408.400 314.400 ;
        RECT 410.800 314.300 411.600 319.800 ;
        RECT 407.600 313.700 411.600 314.300 ;
        RECT 407.600 313.600 408.400 313.700 ;
        RECT 391.600 312.300 393.000 312.400 ;
        RECT 388.400 311.800 393.000 312.300 ;
        RECT 393.600 311.800 394.600 312.400 ;
        RECT 385.200 311.200 385.800 311.800 ;
        RECT 388.400 311.700 392.400 311.800 ;
        RECT 381.200 310.400 382.000 310.800 ;
        RECT 383.800 310.600 385.800 311.200 ;
        RECT 383.800 310.400 384.400 310.600 ;
        RECT 378.800 310.300 379.600 310.400 ;
        RECT 380.400 310.300 382.000 310.400 ;
        RECT 378.800 309.800 382.000 310.300 ;
        RECT 378.800 309.700 381.200 309.800 ;
        RECT 378.800 309.600 379.600 309.700 ;
        RECT 380.400 309.600 381.200 309.700 ;
        RECT 383.600 309.600 384.400 310.400 ;
        RECT 386.800 309.600 387.600 311.200 ;
        RECT 378.800 306.800 379.600 308.400 ;
        RECT 382.000 307.600 382.800 309.200 ;
        RECT 370.200 302.200 371.800 306.200 ;
        RECT 375.600 305.600 378.000 306.400 ;
        RECT 383.800 306.200 384.400 309.600 ;
        RECT 385.000 308.800 385.800 309.600 ;
        RECT 385.200 308.400 385.800 308.800 ;
        RECT 385.200 307.600 386.000 308.400 ;
        RECT 376.200 302.200 377.000 305.600 ;
        RECT 383.400 302.200 385.000 306.200 ;
        RECT 388.400 302.200 389.200 311.700 ;
        RECT 391.600 311.600 392.400 311.700 ;
        RECT 393.600 308.400 394.200 311.800 ;
        RECT 398.000 310.800 398.800 312.400 ;
        RECT 402.800 311.600 403.600 312.400 ;
        RECT 404.400 311.600 405.200 312.400 ;
        RECT 394.800 308.800 395.600 310.400 ;
        RECT 399.600 309.600 401.200 310.400 ;
        RECT 402.800 308.400 403.400 311.600 ;
        RECT 390.000 308.300 390.800 308.400 ;
        RECT 391.600 308.300 394.200 308.400 ;
        RECT 390.000 307.700 394.200 308.300 ;
        RECT 396.400 308.200 397.200 308.400 ;
        RECT 401.800 308.200 403.400 308.400 ;
        RECT 390.000 307.600 390.800 307.700 ;
        RECT 391.600 307.600 394.200 307.700 ;
        RECT 395.600 307.600 397.200 308.200 ;
        RECT 401.600 307.800 403.400 308.200 ;
        RECT 404.600 308.400 405.200 311.600 ;
        RECT 409.200 310.800 410.000 312.400 ;
        RECT 406.800 309.600 408.400 310.400 ;
        RECT 404.600 308.200 406.200 308.400 ;
        RECT 404.600 307.800 406.400 308.200 ;
        RECT 390.000 304.800 390.800 306.400 ;
        RECT 391.800 306.200 392.400 307.600 ;
        RECT 395.600 307.200 396.400 307.600 ;
        RECT 393.400 306.200 397.000 306.600 ;
        RECT 391.600 302.200 392.400 306.200 ;
        RECT 393.200 306.000 397.200 306.200 ;
        RECT 393.200 302.200 394.000 306.000 ;
        RECT 396.400 302.200 397.200 306.000 ;
        RECT 401.600 302.200 402.400 307.800 ;
        RECT 405.600 302.200 406.400 307.800 ;
        RECT 410.800 302.200 411.600 313.700 ;
        RECT 414.600 312.600 415.400 319.800 ;
        RECT 425.200 313.800 426.000 319.800 ;
        RECT 425.400 313.200 426.000 313.800 ;
        RECT 428.400 319.200 432.400 319.800 ;
        RECT 428.400 313.800 429.200 319.200 ;
        RECT 430.000 313.800 430.800 318.600 ;
        RECT 431.600 314.000 432.400 319.200 ;
        RECT 433.400 319.200 437.000 319.800 ;
        RECT 433.400 319.000 434.000 319.200 ;
        RECT 428.400 313.200 429.000 313.800 ;
        RECT 425.400 312.600 429.000 313.200 ;
        RECT 430.200 313.400 430.800 313.800 ;
        RECT 433.200 313.400 434.000 319.000 ;
        RECT 436.400 319.000 437.000 319.200 ;
        RECT 430.200 313.000 434.000 313.400 ;
        RECT 434.800 313.000 435.600 318.600 ;
        RECT 436.400 313.000 437.200 319.000 ;
        RECT 430.200 312.800 433.800 313.000 ;
        RECT 414.600 311.800 416.400 312.600 ;
        RECT 434.800 312.400 435.400 313.000 ;
        RECT 434.800 312.200 435.600 312.400 ;
        RECT 414.000 309.600 414.800 311.200 ;
        RECT 415.600 308.400 416.200 311.800 ;
        RECT 432.200 311.600 435.600 312.200 ;
        RECT 436.400 312.300 437.200 312.400 ;
        RECT 438.000 312.300 438.800 319.800 ;
        RECT 442.800 316.400 443.600 319.800 ;
        RECT 442.600 315.800 443.600 316.400 ;
        RECT 442.600 315.200 443.200 315.800 ;
        RECT 446.000 315.200 446.800 319.800 ;
        RECT 449.200 317.000 450.000 319.800 ;
        RECT 450.800 317.000 451.600 319.800 ;
        RECT 436.400 311.700 438.800 312.300 ;
        RECT 436.400 311.600 437.200 311.700 ;
        RECT 432.200 310.400 432.800 311.600 ;
        RECT 430.000 309.600 431.600 310.400 ;
        RECT 432.200 309.600 434.000 310.400 ;
        RECT 412.400 308.300 413.200 308.400 ;
        RECT 415.600 308.300 416.400 308.400 ;
        RECT 428.400 308.300 430.000 308.400 ;
        RECT 412.400 307.700 416.400 308.300 ;
        RECT 412.400 307.600 413.200 307.700 ;
        RECT 415.600 307.600 416.400 307.700 ;
        RECT 417.300 307.700 430.000 308.300 ;
        RECT 412.400 306.300 413.200 306.400 ;
        RECT 414.000 306.300 414.800 306.400 ;
        RECT 412.400 305.700 414.800 306.300 ;
        RECT 412.400 304.800 413.200 305.700 ;
        RECT 414.000 305.600 414.800 305.700 ;
        RECT 415.600 304.200 416.200 307.600 ;
        RECT 417.300 306.400 417.900 307.700 ;
        RECT 428.400 307.600 430.000 307.700 ;
        RECT 417.200 304.800 418.000 306.400 ;
        RECT 418.800 306.300 419.600 306.400 ;
        RECT 426.800 306.300 429.200 306.400 ;
        RECT 418.800 305.700 429.200 306.300 ;
        RECT 418.800 305.600 419.600 305.700 ;
        RECT 426.800 305.600 429.200 305.700 ;
        RECT 432.200 305.000 432.800 309.600 ;
        RECT 428.800 304.400 432.800 305.000 ;
        RECT 428.800 304.200 429.400 304.400 ;
        RECT 415.600 302.200 416.400 304.200 ;
        RECT 428.400 303.600 429.400 304.200 ;
        RECT 431.600 304.200 432.800 304.400 ;
        RECT 428.400 302.200 429.200 303.600 ;
        RECT 431.600 302.200 432.400 304.200 ;
        RECT 438.000 302.200 438.800 311.700 ;
        RECT 441.200 314.600 443.200 315.200 ;
        RECT 441.200 309.000 442.000 314.600 ;
        RECT 443.800 314.400 448.000 315.200 ;
        RECT 452.400 315.000 453.200 319.800 ;
        RECT 455.600 315.000 456.400 319.800 ;
        RECT 443.800 314.000 444.400 314.400 ;
        RECT 442.800 313.200 444.400 314.000 ;
        RECT 447.400 313.800 453.200 314.400 ;
        RECT 445.400 313.200 446.800 313.800 ;
        RECT 445.400 313.000 451.600 313.200 ;
        RECT 446.200 312.600 451.600 313.000 ;
        RECT 450.800 312.400 451.600 312.600 ;
        RECT 452.600 313.000 453.200 313.800 ;
        RECT 453.800 313.600 456.400 314.400 ;
        RECT 458.800 313.600 459.600 319.800 ;
        RECT 460.400 317.000 461.200 319.800 ;
        RECT 462.000 317.000 462.800 319.800 ;
        RECT 463.600 317.000 464.400 319.800 ;
        RECT 462.000 314.400 466.200 315.200 ;
        RECT 466.800 314.400 467.600 319.800 ;
        RECT 470.000 315.200 470.800 319.800 ;
        RECT 470.000 314.600 472.600 315.200 ;
        RECT 466.800 313.600 469.400 314.400 ;
        RECT 460.400 313.000 461.200 313.200 ;
        RECT 452.600 312.400 461.200 313.000 ;
        RECT 463.600 313.000 464.400 313.200 ;
        RECT 472.000 313.000 472.600 314.600 ;
        RECT 463.600 312.400 472.600 313.000 ;
        RECT 472.000 310.600 472.600 312.400 ;
        RECT 473.200 312.000 474.000 319.800 ;
        RECT 473.200 311.200 474.200 312.000 ;
        RECT 442.600 310.000 466.000 310.600 ;
        RECT 472.000 310.000 472.800 310.600 ;
        RECT 442.600 309.800 443.400 310.000 ;
        RECT 444.400 309.600 445.200 310.000 ;
        RECT 447.600 309.600 448.400 310.000 ;
        RECT 465.200 309.400 466.000 310.000 ;
        RECT 441.200 308.200 450.000 309.000 ;
        RECT 450.600 308.600 452.600 309.400 ;
        RECT 456.400 308.600 459.600 309.400 ;
        RECT 439.600 304.800 440.400 306.400 ;
        RECT 441.200 302.200 442.000 308.200 ;
        RECT 443.600 306.800 446.600 307.600 ;
        RECT 445.800 306.200 446.600 306.800 ;
        RECT 451.800 306.200 452.600 308.600 ;
        RECT 454.000 306.800 454.800 308.400 ;
        RECT 459.200 307.800 460.000 308.000 ;
        RECT 455.600 307.200 460.000 307.800 ;
        RECT 455.600 307.000 456.400 307.200 ;
        RECT 462.000 306.400 462.800 309.200 ;
        RECT 467.800 308.600 471.600 309.400 ;
        RECT 467.800 307.400 468.600 308.600 ;
        RECT 472.200 308.000 472.800 310.000 ;
        RECT 455.600 306.200 456.400 306.400 ;
        RECT 445.800 305.400 448.400 306.200 ;
        RECT 451.800 305.600 456.400 306.200 ;
        RECT 457.200 305.600 458.800 306.400 ;
        RECT 461.800 305.600 462.800 306.400 ;
        RECT 466.800 306.800 468.600 307.400 ;
        RECT 471.600 307.400 472.800 308.000 ;
        RECT 466.800 306.200 467.600 306.800 ;
        RECT 447.600 302.200 448.400 305.400 ;
        RECT 465.200 305.400 467.600 306.200 ;
        RECT 449.200 302.200 450.000 305.000 ;
        RECT 450.800 302.200 451.600 305.000 ;
        RECT 452.400 302.200 453.200 305.000 ;
        RECT 455.600 302.200 456.400 305.000 ;
        RECT 458.800 302.200 459.600 305.000 ;
        RECT 460.400 302.200 461.200 305.000 ;
        RECT 462.000 302.200 462.800 305.000 ;
        RECT 463.600 302.200 464.400 305.000 ;
        RECT 465.200 302.200 466.000 305.400 ;
        RECT 471.600 302.200 472.400 307.400 ;
        RECT 473.400 306.800 474.200 311.200 ;
        RECT 473.200 306.300 474.200 306.800 ;
        RECT 476.400 306.300 477.200 306.400 ;
        RECT 473.200 305.700 477.200 306.300 ;
        RECT 473.200 302.200 474.000 305.700 ;
        RECT 476.400 304.800 477.200 305.700 ;
        RECT 478.000 302.200 478.800 319.800 ;
        RECT 481.200 311.200 482.000 319.800 ;
        RECT 484.400 311.200 485.200 319.800 ;
        RECT 487.600 311.200 488.400 319.800 ;
        RECT 490.800 311.200 491.600 319.800 ;
        RECT 479.600 310.400 482.000 311.200 ;
        RECT 483.000 310.400 485.200 311.200 ;
        RECT 486.200 310.400 488.400 311.200 ;
        RECT 489.800 310.400 491.600 311.200 ;
        RECT 479.600 307.600 480.400 310.400 ;
        RECT 483.000 309.000 483.800 310.400 ;
        RECT 486.200 309.000 487.000 310.400 ;
        RECT 489.800 309.000 490.600 310.400 ;
        RECT 481.200 308.200 483.800 309.000 ;
        RECT 484.600 308.200 487.000 309.000 ;
        RECT 488.000 308.200 490.600 309.000 ;
        RECT 483.000 307.600 483.800 308.200 ;
        RECT 486.200 307.600 487.000 308.200 ;
        RECT 489.800 307.600 490.600 308.200 ;
        RECT 479.600 306.800 482.000 307.600 ;
        RECT 483.000 306.800 485.200 307.600 ;
        RECT 486.200 306.800 488.400 307.600 ;
        RECT 489.800 306.800 491.600 307.600 ;
        RECT 481.200 302.200 482.000 306.800 ;
        RECT 484.400 302.200 485.200 306.800 ;
        RECT 487.600 302.200 488.400 306.800 ;
        RECT 490.800 302.200 491.600 306.800 ;
        RECT 494.000 304.800 494.800 306.400 ;
        RECT 495.600 302.200 496.400 319.800 ;
        RECT 497.400 319.200 501.000 319.800 ;
        RECT 497.400 319.000 498.000 319.200 ;
        RECT 497.200 313.000 498.000 319.000 ;
        RECT 500.400 319.000 501.000 319.200 ;
        RECT 502.000 319.200 506.000 319.800 ;
        RECT 498.800 313.000 499.600 318.600 ;
        RECT 500.400 313.400 501.200 319.000 ;
        RECT 502.000 314.000 502.800 319.200 ;
        RECT 503.600 313.800 504.400 318.600 ;
        RECT 505.200 313.800 506.000 319.200 ;
        RECT 503.600 313.400 504.200 313.800 ;
        RECT 500.400 313.000 504.200 313.400 ;
        RECT 499.000 312.400 499.600 313.000 ;
        RECT 500.600 312.800 504.200 313.000 ;
        RECT 505.400 313.200 506.000 313.800 ;
        RECT 508.400 313.800 509.200 319.800 ;
        RECT 508.400 313.200 509.000 313.800 ;
        RECT 505.400 312.600 509.000 313.200 ;
        RECT 498.800 312.200 499.600 312.400 ;
        RECT 512.600 312.400 513.400 319.800 ;
        RECT 514.000 313.600 514.800 314.400 ;
        RECT 514.200 312.400 514.800 313.600 ;
        RECT 498.800 311.600 502.200 312.200 ;
        RECT 512.600 311.800 513.600 312.400 ;
        RECT 514.200 311.800 515.600 312.400 ;
        RECT 501.600 305.000 502.200 311.600 ;
        RECT 502.800 309.600 504.400 310.400 ;
        RECT 510.000 309.600 510.800 310.400 ;
        RECT 510.100 308.400 510.700 309.600 ;
        RECT 511.600 308.800 512.400 310.400 ;
        RECT 513.000 308.400 513.600 311.800 ;
        RECT 514.800 311.600 515.600 311.800 ;
        RECT 518.000 310.300 518.800 319.800 ;
        RECT 519.600 312.400 520.400 319.800 ;
        RECT 522.800 312.400 523.600 319.800 ;
        RECT 519.600 311.800 523.600 312.400 ;
        RECT 524.400 311.800 525.200 319.800 ;
        RECT 520.400 310.400 521.200 310.800 ;
        RECT 524.400 310.400 525.000 311.800 ;
        RECT 519.600 310.300 521.200 310.400 ;
        RECT 518.000 309.800 521.200 310.300 ;
        RECT 522.800 309.800 525.200 310.400 ;
        RECT 518.000 309.700 520.400 309.800 ;
        RECT 504.400 308.300 506.000 308.400 ;
        RECT 508.400 308.300 509.200 308.400 ;
        RECT 504.400 307.700 509.200 308.300 ;
        RECT 504.400 307.600 506.000 307.700 ;
        RECT 508.400 307.600 509.200 307.700 ;
        RECT 510.000 308.200 510.800 308.400 ;
        RECT 510.000 307.600 511.600 308.200 ;
        RECT 513.000 307.600 515.600 308.400 ;
        RECT 510.800 307.200 511.600 307.600 ;
        RECT 505.800 305.600 507.600 306.400 ;
        RECT 510.200 306.200 513.800 306.600 ;
        RECT 514.800 306.200 515.400 307.600 ;
        RECT 510.000 306.000 514.000 306.200 ;
        RECT 501.600 304.400 505.600 305.000 ;
        RECT 501.600 304.200 502.800 304.400 ;
        RECT 502.000 302.200 502.800 304.200 ;
        RECT 505.000 304.200 505.600 304.400 ;
        RECT 505.000 303.600 506.000 304.200 ;
        RECT 505.200 302.200 506.000 303.600 ;
        RECT 510.000 302.200 510.800 306.000 ;
        RECT 513.200 302.200 514.000 306.000 ;
        RECT 514.800 302.200 515.600 306.200 ;
        RECT 516.400 304.800 517.200 306.400 ;
        RECT 518.000 302.200 518.800 309.700 ;
        RECT 519.600 309.600 520.400 309.700 ;
        RECT 521.200 307.600 522.000 309.200 ;
        RECT 522.800 306.200 523.400 309.800 ;
        RECT 524.400 309.600 525.200 309.800 ;
        RECT 527.600 308.300 528.400 319.800 ;
        RECT 531.800 312.400 532.600 319.800 ;
        RECT 533.200 313.600 534.000 314.400 ;
        RECT 533.400 312.400 534.000 313.600 ;
        RECT 538.200 312.400 539.000 319.800 ;
        RECT 539.600 313.600 540.400 314.400 ;
        RECT 539.800 312.400 540.400 313.600 ;
        RECT 531.800 311.800 532.800 312.400 ;
        RECT 533.400 311.800 534.800 312.400 ;
        RECT 530.800 308.800 531.600 310.400 ;
        RECT 532.200 308.400 532.800 311.800 ;
        RECT 534.000 311.600 534.800 311.800 ;
        RECT 537.200 311.600 539.200 312.400 ;
        RECT 539.800 311.800 541.200 312.400 ;
        RECT 540.400 311.600 541.200 311.800 ;
        RECT 537.200 308.800 538.000 310.400 ;
        RECT 538.600 308.400 539.200 311.600 ;
        RECT 529.200 308.300 530.000 308.400 ;
        RECT 527.600 308.200 530.000 308.300 ;
        RECT 527.600 307.700 530.800 308.200 ;
        RECT 522.800 302.200 523.600 306.200 ;
        RECT 524.400 305.600 525.200 306.400 ;
        RECT 524.200 304.800 525.000 305.600 ;
        RECT 526.000 304.800 526.800 306.400 ;
        RECT 527.600 302.200 528.400 307.700 ;
        RECT 529.200 307.600 530.800 307.700 ;
        RECT 532.200 307.600 534.800 308.400 ;
        RECT 535.600 308.200 536.400 308.400 ;
        RECT 535.600 307.600 537.200 308.200 ;
        RECT 538.600 307.600 541.200 308.400 ;
        RECT 530.000 307.200 530.800 307.600 ;
        RECT 529.400 306.200 533.000 306.600 ;
        RECT 534.000 306.200 534.600 307.600 ;
        RECT 536.400 307.200 537.200 307.600 ;
        RECT 535.800 306.200 539.400 306.600 ;
        RECT 540.400 306.200 541.000 307.600 ;
        RECT 543.600 306.200 544.400 319.800 ;
        RECT 529.200 306.000 533.200 306.200 ;
        RECT 529.200 302.200 530.000 306.000 ;
        RECT 532.400 302.200 533.200 306.000 ;
        RECT 534.000 302.200 534.800 306.200 ;
        RECT 535.600 306.000 539.600 306.200 ;
        RECT 535.600 302.200 536.400 306.000 ;
        RECT 538.800 302.200 539.600 306.000 ;
        RECT 540.400 302.200 541.200 306.200 ;
        RECT 542.600 305.600 544.400 306.200 ;
        RECT 542.600 304.400 543.400 305.600 ;
        RECT 542.600 303.600 544.400 304.400 ;
        RECT 542.600 302.200 543.400 303.600 ;
        RECT 2.400 294.200 3.200 299.800 ;
        RECT 1.400 293.800 3.200 294.200 ;
        RECT 1.400 293.600 3.000 293.800 ;
        RECT 1.400 290.400 2.000 293.600 ;
        RECT 3.600 291.600 5.200 292.400 ;
        RECT 1.200 289.600 2.000 290.400 ;
        RECT 6.000 289.600 6.800 291.200 ;
        RECT 1.400 287.000 2.000 289.600 ;
        RECT 2.800 288.300 3.600 289.200 ;
        RECT 7.600 288.300 8.400 299.800 ;
        RECT 12.400 297.800 13.200 299.800 ;
        RECT 9.200 296.300 10.000 297.200 ;
        RECT 10.800 296.300 11.600 297.200 ;
        RECT 12.600 296.400 13.200 297.800 ;
        RECT 9.200 295.700 11.600 296.300 ;
        RECT 9.200 295.600 10.000 295.700 ;
        RECT 10.800 295.600 11.600 295.700 ;
        RECT 12.400 295.600 13.200 296.400 ;
        RECT 14.000 296.300 14.800 296.400 ;
        RECT 15.600 296.300 16.400 297.200 ;
        RECT 14.000 295.700 16.400 296.300 ;
        RECT 14.000 295.600 14.800 295.700 ;
        RECT 15.600 295.600 16.400 295.700 ;
        RECT 12.600 294.400 13.200 295.600 ;
        RECT 12.400 293.600 13.200 294.400 ;
        RECT 12.600 290.200 13.200 293.600 ;
        RECT 14.000 290.800 14.800 292.400 ;
        RECT 12.400 289.400 14.200 290.200 ;
        RECT 2.800 287.700 8.400 288.300 ;
        RECT 2.800 287.600 3.600 287.700 ;
        RECT 1.400 286.400 5.000 287.000 ;
        RECT 1.400 286.200 2.000 286.400 ;
        RECT 1.200 282.200 2.000 286.200 ;
        RECT 4.400 286.200 5.000 286.400 ;
        RECT 4.400 282.200 5.200 286.200 ;
        RECT 7.600 282.200 8.400 287.700 ;
        RECT 13.400 282.200 14.200 289.400 ;
        RECT 17.200 288.300 18.000 299.800 ;
        RECT 18.800 295.600 19.600 297.200 ;
        RECT 18.800 288.300 19.600 288.400 ;
        RECT 17.200 287.700 19.600 288.300 ;
        RECT 17.200 282.200 18.000 287.700 ;
        RECT 18.800 287.600 19.600 287.700 ;
        RECT 20.400 282.200 21.200 299.800 ;
        RECT 25.600 294.200 26.400 299.800 ;
        RECT 29.000 298.400 29.800 299.800 ;
        RECT 28.400 297.600 29.800 298.400 ;
        RECT 34.800 297.800 35.600 299.800 ;
        RECT 29.000 296.400 29.800 297.600 ;
        RECT 29.000 295.800 30.800 296.400 ;
        RECT 25.600 293.800 27.400 294.200 ;
        RECT 25.800 293.600 27.400 293.800 ;
        RECT 23.600 291.600 25.200 292.400 ;
        RECT 22.000 289.600 22.800 291.200 ;
        RECT 26.800 290.400 27.400 293.600 ;
        RECT 26.800 289.600 27.600 290.400 ;
        RECT 25.200 287.600 26.000 289.200 ;
        RECT 26.800 287.000 27.400 289.600 ;
        RECT 28.400 288.800 29.200 290.400 ;
        RECT 23.800 286.400 27.400 287.000 ;
        RECT 23.800 286.200 24.400 286.400 ;
        RECT 23.600 282.200 24.400 286.200 ;
        RECT 26.800 286.200 27.400 286.400 ;
        RECT 26.800 282.200 27.600 286.200 ;
        RECT 30.000 282.200 30.800 295.800 ;
        RECT 33.200 295.600 34.000 297.200 ;
        RECT 31.600 294.300 32.400 295.200 ;
        RECT 35.000 294.400 35.600 297.800 ;
        RECT 39.600 296.000 40.400 299.800 ;
        RECT 33.200 294.300 34.000 294.400 ;
        RECT 31.600 293.700 34.000 294.300 ;
        RECT 31.600 293.600 32.400 293.700 ;
        RECT 33.200 293.600 34.000 293.700 ;
        RECT 34.800 293.600 35.600 294.400 ;
        RECT 35.000 290.200 35.600 293.600 ;
        RECT 39.400 295.200 40.400 296.000 ;
        RECT 36.400 290.800 37.200 292.400 ;
        RECT 39.400 290.800 40.200 295.200 ;
        RECT 41.200 294.600 42.000 299.800 ;
        RECT 47.600 296.600 48.400 299.800 ;
        RECT 49.200 297.000 50.000 299.800 ;
        RECT 50.800 297.000 51.600 299.800 ;
        RECT 52.400 297.000 53.200 299.800 ;
        RECT 54.000 297.000 54.800 299.800 ;
        RECT 57.200 297.000 58.000 299.800 ;
        RECT 60.400 297.000 61.200 299.800 ;
        RECT 62.000 297.000 62.800 299.800 ;
        RECT 63.600 297.000 64.400 299.800 ;
        RECT 46.000 295.800 48.400 296.600 ;
        RECT 65.200 296.600 66.000 299.800 ;
        RECT 46.000 295.200 46.800 295.800 ;
        RECT 40.800 294.000 42.000 294.600 ;
        RECT 45.000 294.600 46.800 295.200 ;
        RECT 50.800 295.600 51.800 296.400 ;
        RECT 54.800 295.600 56.400 296.400 ;
        RECT 57.200 295.800 61.800 296.400 ;
        RECT 65.200 295.800 67.800 296.600 ;
        RECT 57.200 295.600 58.000 295.800 ;
        RECT 40.800 292.000 41.400 294.000 ;
        RECT 45.000 293.400 45.800 294.600 ;
        RECT 42.000 292.600 45.800 293.400 ;
        RECT 50.800 292.800 51.600 295.600 ;
        RECT 57.200 294.800 58.000 295.000 ;
        RECT 53.600 294.200 58.000 294.800 ;
        RECT 53.600 294.000 54.400 294.200 ;
        RECT 58.800 293.600 59.600 295.200 ;
        RECT 61.000 293.400 61.800 295.800 ;
        RECT 67.000 295.200 67.800 295.800 ;
        RECT 67.000 294.400 70.000 295.200 ;
        RECT 71.600 293.800 72.400 299.800 ;
        RECT 74.800 296.000 75.600 299.800 ;
        RECT 54.000 292.600 57.200 293.400 ;
        RECT 61.000 292.600 63.000 293.400 ;
        RECT 63.600 293.000 72.400 293.800 ;
        RECT 47.600 292.000 48.400 292.600 ;
        RECT 65.200 292.000 66.000 292.400 ;
        RECT 68.400 292.000 69.200 292.400 ;
        RECT 70.200 292.000 71.000 292.200 ;
        RECT 40.800 291.400 41.600 292.000 ;
        RECT 47.600 291.400 71.000 292.000 ;
        RECT 34.800 289.400 36.600 290.200 ;
        RECT 39.400 290.000 40.400 290.800 ;
        RECT 35.800 284.400 36.600 289.400 ;
        RECT 35.800 283.600 37.200 284.400 ;
        RECT 35.800 282.200 36.600 283.600 ;
        RECT 39.600 282.200 40.400 290.000 ;
        RECT 41.000 289.600 41.600 291.400 ;
        RECT 41.000 289.000 50.000 289.600 ;
        RECT 41.000 287.400 41.600 289.000 ;
        RECT 49.200 288.800 50.000 289.000 ;
        RECT 52.400 289.000 61.000 289.600 ;
        RECT 52.400 288.800 53.200 289.000 ;
        RECT 44.200 287.600 46.800 288.400 ;
        RECT 41.000 286.800 43.600 287.400 ;
        RECT 42.800 282.200 43.600 286.800 ;
        RECT 46.000 282.200 46.800 287.600 ;
        RECT 47.400 286.800 51.600 287.600 ;
        RECT 49.200 282.200 50.000 285.000 ;
        RECT 50.800 282.200 51.600 285.000 ;
        RECT 52.400 282.200 53.200 285.000 ;
        RECT 54.000 282.200 54.800 288.400 ;
        RECT 57.200 287.600 59.800 288.400 ;
        RECT 60.400 288.200 61.000 289.000 ;
        RECT 62.000 289.400 62.800 289.600 ;
        RECT 62.000 289.000 67.400 289.400 ;
        RECT 62.000 288.800 68.200 289.000 ;
        RECT 66.800 288.200 68.200 288.800 ;
        RECT 60.400 287.600 66.200 288.200 ;
        RECT 69.200 288.000 70.800 288.800 ;
        RECT 69.200 287.600 69.800 288.000 ;
        RECT 57.200 282.200 58.000 287.000 ;
        RECT 60.400 282.200 61.200 287.000 ;
        RECT 65.600 286.800 69.800 287.600 ;
        RECT 71.600 287.400 72.400 293.000 ;
        RECT 74.600 295.200 75.600 296.000 ;
        RECT 74.600 290.800 75.400 295.200 ;
        RECT 76.400 294.600 77.200 299.800 ;
        RECT 82.800 296.600 83.600 299.800 ;
        RECT 84.400 297.000 85.200 299.800 ;
        RECT 86.000 297.000 86.800 299.800 ;
        RECT 87.600 297.000 88.400 299.800 ;
        RECT 89.200 297.000 90.000 299.800 ;
        RECT 92.400 297.000 93.200 299.800 ;
        RECT 95.600 297.000 96.400 299.800 ;
        RECT 97.200 297.000 98.000 299.800 ;
        RECT 98.800 297.000 99.600 299.800 ;
        RECT 81.200 295.800 83.600 296.600 ;
        RECT 100.400 296.600 101.200 299.800 ;
        RECT 81.200 295.200 82.000 295.800 ;
        RECT 76.000 294.000 77.200 294.600 ;
        RECT 80.200 294.600 82.000 295.200 ;
        RECT 86.000 295.600 87.000 296.400 ;
        RECT 90.000 295.600 91.600 296.400 ;
        RECT 92.400 295.800 97.000 296.400 ;
        RECT 100.400 295.800 103.000 296.600 ;
        RECT 92.400 295.600 93.200 295.800 ;
        RECT 76.000 292.000 76.600 294.000 ;
        RECT 80.200 293.400 81.000 294.600 ;
        RECT 77.200 292.600 81.000 293.400 ;
        RECT 86.000 292.800 86.800 295.600 ;
        RECT 92.400 294.800 93.200 295.000 ;
        RECT 88.800 294.200 93.200 294.800 ;
        RECT 88.800 294.000 89.600 294.200 ;
        RECT 94.000 293.600 94.800 295.200 ;
        RECT 96.200 293.400 97.000 295.800 ;
        RECT 102.200 295.200 103.000 295.800 ;
        RECT 102.200 294.400 105.200 295.200 ;
        RECT 106.800 293.800 107.600 299.800 ;
        RECT 109.000 296.400 109.800 299.800 ;
        RECT 108.400 295.600 110.800 296.400 ;
        RECT 113.200 295.800 114.000 299.800 ;
        RECT 114.800 296.000 115.600 299.800 ;
        RECT 118.000 296.000 118.800 299.800 ;
        RECT 121.200 297.800 122.000 299.800 ;
        RECT 114.800 295.800 118.800 296.000 ;
        RECT 89.200 292.600 92.400 293.400 ;
        RECT 96.200 292.600 98.200 293.400 ;
        RECT 98.800 293.000 107.600 293.800 ;
        RECT 82.800 292.000 83.600 292.600 ;
        RECT 100.400 292.000 101.200 292.400 ;
        RECT 103.600 292.000 104.400 292.400 ;
        RECT 105.400 292.000 106.200 292.200 ;
        RECT 76.000 291.400 76.800 292.000 ;
        RECT 82.800 291.400 106.200 292.000 ;
        RECT 74.600 290.000 75.600 290.800 ;
        RECT 70.400 286.800 72.400 287.400 ;
        RECT 62.000 282.200 62.800 285.000 ;
        RECT 63.600 282.200 64.400 285.000 ;
        RECT 66.800 282.200 67.600 286.800 ;
        RECT 70.400 286.200 71.000 286.800 ;
        RECT 70.000 285.600 71.000 286.200 ;
        RECT 70.000 282.200 70.800 285.600 ;
        RECT 74.800 282.200 75.600 290.000 ;
        RECT 76.200 289.600 76.800 291.400 ;
        RECT 76.200 289.000 85.200 289.600 ;
        RECT 76.200 287.400 76.800 289.000 ;
        RECT 84.400 288.800 85.200 289.000 ;
        RECT 87.600 289.000 96.200 289.600 ;
        RECT 87.600 288.800 88.400 289.000 ;
        RECT 79.400 287.600 82.000 288.400 ;
        RECT 76.200 286.800 78.800 287.400 ;
        RECT 78.000 282.200 78.800 286.800 ;
        RECT 81.200 282.200 82.000 287.600 ;
        RECT 82.600 286.800 86.800 287.600 ;
        RECT 84.400 282.200 85.200 285.000 ;
        RECT 86.000 282.200 86.800 285.000 ;
        RECT 87.600 282.200 88.400 285.000 ;
        RECT 89.200 282.200 90.000 288.400 ;
        RECT 92.400 287.600 95.000 288.400 ;
        RECT 95.600 288.200 96.200 289.000 ;
        RECT 97.200 289.400 98.000 289.600 ;
        RECT 97.200 289.000 102.600 289.400 ;
        RECT 97.200 288.800 103.400 289.000 ;
        RECT 102.000 288.200 103.400 288.800 ;
        RECT 95.600 287.600 101.400 288.200 ;
        RECT 104.400 288.000 106.000 288.800 ;
        RECT 104.400 287.600 105.000 288.000 ;
        RECT 92.400 282.200 93.200 287.000 ;
        RECT 95.600 282.200 96.400 287.000 ;
        RECT 100.800 286.800 105.000 287.600 ;
        RECT 106.800 287.400 107.600 293.000 ;
        RECT 108.400 288.800 109.200 290.400 ;
        RECT 105.600 286.800 107.600 287.400 ;
        RECT 97.200 282.200 98.000 285.000 ;
        RECT 98.800 282.200 99.600 285.000 ;
        RECT 102.000 282.200 102.800 286.800 ;
        RECT 105.600 286.200 106.200 286.800 ;
        RECT 105.200 285.600 106.200 286.200 ;
        RECT 105.200 282.200 106.000 285.600 ;
        RECT 110.000 282.200 110.800 295.600 ;
        RECT 111.600 294.300 112.400 295.200 ;
        RECT 113.400 294.400 114.000 295.800 ;
        RECT 115.000 295.400 118.600 295.800 ;
        RECT 119.600 295.600 120.400 297.200 ;
        RECT 117.200 294.400 118.000 294.800 ;
        RECT 121.400 294.400 122.000 297.800 ;
        RECT 130.800 296.000 131.600 299.800 ;
        RECT 134.000 296.000 134.800 299.800 ;
        RECT 130.800 295.800 134.800 296.000 ;
        RECT 135.600 295.800 136.400 299.800 ;
        RECT 131.000 295.400 134.600 295.800 ;
        RECT 131.600 294.400 132.400 294.800 ;
        RECT 135.600 294.400 136.200 295.800 ;
        RECT 137.200 295.600 138.000 297.200 ;
        RECT 113.200 294.300 115.800 294.400 ;
        RECT 111.600 293.700 115.800 294.300 ;
        RECT 117.200 293.800 118.800 294.400 ;
        RECT 111.600 293.600 112.400 293.700 ;
        RECT 113.200 293.600 115.800 293.700 ;
        RECT 118.000 293.600 118.800 293.800 ;
        RECT 121.200 293.600 122.000 294.400 ;
        RECT 129.200 294.300 130.000 294.400 ;
        RECT 130.800 294.300 132.400 294.400 ;
        RECT 129.200 293.800 132.400 294.300 ;
        RECT 129.200 293.700 131.600 293.800 ;
        RECT 129.200 293.600 130.000 293.700 ;
        RECT 130.800 293.600 131.600 293.700 ;
        RECT 133.800 293.600 136.400 294.400 ;
        RECT 138.800 294.300 139.600 299.800 ;
        RECT 140.400 296.000 141.200 299.800 ;
        RECT 143.600 296.000 144.400 299.800 ;
        RECT 140.400 295.800 144.400 296.000 ;
        RECT 145.200 295.800 146.000 299.800 ;
        RECT 140.600 295.400 144.200 295.800 ;
        RECT 141.200 294.400 142.000 294.800 ;
        RECT 145.200 294.400 145.800 295.800 ;
        RECT 140.400 294.300 142.000 294.400 ;
        RECT 138.800 293.800 142.000 294.300 ;
        RECT 138.800 293.700 141.200 293.800 ;
        RECT 113.200 290.200 114.000 290.400 ;
        RECT 115.200 290.200 115.800 293.600 ;
        RECT 116.400 291.600 117.200 293.200 ;
        RECT 121.400 290.200 122.000 293.600 ;
        RECT 122.800 290.800 123.600 292.400 ;
        RECT 126.000 292.300 126.800 292.400 ;
        RECT 132.400 292.300 133.200 293.200 ;
        RECT 126.000 291.700 133.200 292.300 ;
        RECT 126.000 291.600 126.800 291.700 ;
        RECT 132.400 291.600 133.200 291.700 ;
        RECT 133.800 292.300 134.400 293.600 ;
        RECT 137.200 292.300 138.000 292.400 ;
        RECT 133.800 291.700 138.000 292.300 ;
        RECT 133.800 290.200 134.400 291.700 ;
        RECT 137.200 291.600 138.000 291.700 ;
        RECT 135.600 290.200 136.400 290.400 ;
        RECT 113.200 289.600 114.600 290.200 ;
        RECT 115.200 289.600 116.200 290.200 ;
        RECT 114.000 288.400 114.600 289.600 ;
        RECT 114.000 287.600 114.800 288.400 ;
        RECT 115.400 282.200 116.200 289.600 ;
        RECT 121.200 289.400 123.000 290.200 ;
        RECT 122.200 288.300 123.000 289.400 ;
        RECT 133.400 289.600 134.400 290.200 ;
        RECT 135.000 289.600 136.400 290.200 ;
        RECT 129.200 288.300 130.000 288.400 ;
        RECT 122.200 287.700 130.000 288.300 ;
        RECT 122.200 282.200 123.000 287.700 ;
        RECT 129.200 287.600 130.000 287.700 ;
        RECT 133.400 282.200 134.200 289.600 ;
        RECT 135.000 288.400 135.600 289.600 ;
        RECT 134.800 287.600 135.600 288.400 ;
        RECT 138.800 282.200 139.600 293.700 ;
        RECT 140.400 293.600 141.200 293.700 ;
        RECT 143.400 293.600 146.000 294.400 ;
        RECT 148.000 294.200 148.800 299.800 ;
        RECT 147.000 293.800 148.800 294.200 ;
        RECT 154.800 297.800 155.600 299.800 ;
        RECT 154.800 294.400 155.400 297.800 ;
        RECT 156.400 295.600 157.200 297.200 ;
        RECT 158.000 296.000 158.800 299.800 ;
        RECT 161.200 296.000 162.000 299.800 ;
        RECT 158.000 295.800 162.000 296.000 ;
        RECT 162.800 295.800 163.600 299.800 ;
        RECT 167.000 298.400 167.800 299.800 ;
        RECT 166.000 297.600 167.800 298.400 ;
        RECT 170.800 297.800 171.600 299.800 ;
        RECT 167.000 296.400 167.800 297.600 ;
        RECT 166.000 295.800 167.800 296.400 ;
        RECT 158.200 295.400 161.800 295.800 ;
        RECT 158.800 294.400 159.600 294.800 ;
        RECT 162.800 294.400 163.400 295.800 ;
        RECT 147.000 293.600 148.600 293.800 ;
        RECT 154.800 293.600 155.600 294.400 ;
        RECT 158.000 293.800 159.600 294.400 ;
        RECT 158.000 293.600 158.800 293.800 ;
        RECT 161.000 293.600 163.600 294.400 ;
        RECT 164.400 293.600 165.200 295.200 ;
        RECT 142.000 291.600 142.800 293.200 ;
        RECT 143.400 290.200 144.000 293.600 ;
        RECT 147.000 290.400 147.600 293.600 ;
        RECT 154.800 292.400 155.400 293.600 ;
        RECT 149.200 291.600 150.800 292.400 ;
        RECT 145.200 290.200 146.000 290.400 ;
        RECT 143.000 289.600 144.000 290.200 ;
        RECT 144.600 289.600 146.000 290.200 ;
        RECT 146.800 289.600 147.600 290.400 ;
        RECT 151.600 289.600 152.400 291.200 ;
        RECT 153.200 290.800 154.000 292.400 ;
        RECT 154.800 291.600 155.600 292.400 ;
        RECT 159.600 291.600 160.400 293.200 ;
        RECT 154.800 290.200 155.400 291.600 ;
        RECT 161.000 290.200 161.600 293.600 ;
        RECT 162.800 290.200 163.600 290.400 ;
        RECT 143.000 282.200 143.800 289.600 ;
        RECT 144.600 288.400 145.200 289.600 ;
        RECT 144.400 287.600 145.200 288.400 ;
        RECT 147.000 287.000 147.600 289.600 ;
        RECT 153.800 289.400 155.600 290.200 ;
        RECT 160.600 289.600 161.600 290.200 ;
        RECT 162.200 289.600 163.600 290.200 ;
        RECT 148.400 287.600 149.200 289.200 ;
        RECT 147.000 286.400 150.600 287.000 ;
        RECT 147.000 286.200 147.600 286.400 ;
        RECT 146.800 282.200 147.600 286.200 ;
        RECT 150.000 286.200 150.600 286.400 ;
        RECT 150.000 282.200 150.800 286.200 ;
        RECT 153.800 282.200 154.600 289.400 ;
        RECT 160.600 282.200 161.400 289.600 ;
        RECT 162.200 288.400 162.800 289.600 ;
        RECT 162.000 287.600 162.800 288.400 ;
        RECT 166.000 282.200 166.800 295.800 ;
        RECT 169.200 295.600 170.000 297.200 ;
        RECT 171.000 294.400 171.600 297.800 ;
        RECT 177.000 295.800 178.600 299.800 ;
        RECT 182.600 296.400 183.400 299.800 ;
        RECT 182.600 295.800 184.400 296.400 ;
        RECT 186.800 295.800 187.600 299.800 ;
        RECT 188.400 296.000 189.200 299.800 ;
        RECT 191.600 296.000 192.400 299.800 ;
        RECT 188.400 295.800 192.400 296.000 ;
        RECT 193.200 295.800 194.000 299.800 ;
        RECT 196.400 297.800 197.200 299.800 ;
        RECT 202.200 298.400 203.800 299.800 ;
        RECT 170.800 293.600 171.600 294.400 ;
        RECT 167.600 292.300 168.400 292.400 ;
        RECT 171.000 292.300 171.600 293.600 ;
        RECT 175.600 292.800 176.400 294.400 ;
        RECT 177.400 292.400 178.000 295.800 ;
        RECT 178.800 294.300 179.600 294.400 ;
        RECT 180.400 294.300 181.200 294.400 ;
        RECT 178.800 293.700 181.200 294.300 ;
        RECT 178.800 293.600 179.600 293.700 ;
        RECT 180.400 293.600 181.200 293.700 ;
        RECT 178.800 293.200 179.400 293.600 ;
        RECT 178.600 292.400 179.400 293.200 ;
        RECT 167.600 291.700 171.600 292.300 ;
        RECT 167.600 291.600 168.400 291.700 ;
        RECT 167.600 288.800 168.400 290.400 ;
        RECT 171.000 290.200 171.600 291.700 ;
        RECT 172.400 290.800 173.200 292.400 ;
        RECT 174.000 292.200 174.800 292.400 ;
        RECT 174.000 291.600 175.600 292.200 ;
        RECT 177.200 291.600 178.000 292.400 ;
        RECT 174.800 291.200 175.600 291.600 ;
        RECT 177.400 291.400 178.000 291.600 ;
        RECT 180.400 292.300 181.200 292.400 ;
        RECT 183.600 292.300 184.400 295.800 ;
        RECT 185.200 294.300 186.000 295.200 ;
        RECT 187.000 294.400 187.600 295.800 ;
        RECT 188.600 295.400 192.200 295.800 ;
        RECT 190.800 294.400 191.600 294.800 ;
        RECT 186.800 294.300 189.400 294.400 ;
        RECT 185.200 293.700 189.400 294.300 ;
        RECT 190.800 293.800 192.400 294.400 ;
        RECT 185.200 293.600 186.000 293.700 ;
        RECT 186.800 293.600 189.400 293.700 ;
        RECT 191.600 293.600 192.400 293.800 ;
        RECT 180.400 291.700 184.400 292.300 ;
        RECT 177.400 290.800 179.400 291.400 ;
        RECT 180.400 290.800 181.200 291.700 ;
        RECT 178.800 290.200 179.400 290.800 ;
        RECT 170.800 289.400 172.600 290.200 ;
        RECT 171.800 282.200 172.600 289.400 ;
        RECT 174.000 289.600 178.000 290.200 ;
        RECT 174.000 282.200 174.800 289.600 ;
        RECT 177.200 282.800 178.000 289.600 ;
        RECT 178.800 283.400 179.600 290.200 ;
        RECT 180.400 282.800 181.200 290.200 ;
        RECT 182.000 288.800 182.800 290.400 ;
        RECT 177.200 282.200 181.200 282.800 ;
        RECT 183.600 282.200 184.400 291.700 ;
        RECT 185.200 290.300 186.000 290.400 ;
        RECT 186.800 290.300 187.600 290.400 ;
        RECT 185.200 290.200 187.600 290.300 ;
        RECT 188.800 290.200 189.400 293.600 ;
        RECT 190.000 291.600 190.800 293.200 ;
        RECT 193.200 292.400 193.800 295.800 ;
        RECT 196.400 295.600 197.000 297.800 ;
        RECT 201.200 297.600 203.800 298.400 ;
        RECT 198.000 295.600 198.800 297.200 ;
        RECT 202.200 295.800 203.800 297.600 ;
        RECT 207.600 295.800 208.400 299.800 ;
        RECT 210.800 297.800 211.600 299.800 ;
        RECT 194.600 295.000 197.000 295.600 ;
        RECT 193.200 291.600 194.000 292.400 ;
        RECT 194.600 292.000 195.200 295.000 ;
        RECT 196.200 293.600 197.200 294.400 ;
        RECT 201.200 293.600 202.000 294.400 ;
        RECT 196.000 292.800 196.800 293.600 ;
        RECT 201.400 293.200 202.000 293.600 ;
        RECT 201.400 292.400 202.200 293.200 ;
        RECT 202.800 292.400 203.400 295.800 ;
        RECT 204.400 292.800 205.200 294.400 ;
        RECT 207.600 292.400 208.200 295.800 ;
        RECT 210.800 295.600 211.400 297.800 ;
        RECT 212.400 295.600 213.200 297.200 ;
        RECT 214.600 296.400 215.400 299.800 ;
        RECT 221.400 298.400 223.000 299.800 ;
        RECT 220.400 297.600 223.000 298.400 ;
        RECT 214.600 295.800 216.400 296.400 ;
        RECT 221.400 295.800 223.000 297.600 ;
        RECT 229.400 295.800 231.000 299.800 ;
        RECT 237.400 295.800 239.000 299.800 ;
        RECT 242.800 295.800 243.600 299.800 ;
        RECT 247.000 296.800 247.800 299.800 ;
        RECT 247.000 295.800 248.400 296.800 ;
        RECT 209.000 295.000 211.400 295.600 ;
        RECT 193.200 290.200 193.800 291.600 ;
        RECT 194.600 291.400 195.400 292.000 ;
        RECT 194.600 291.200 198.800 291.400 ;
        RECT 194.800 290.800 198.800 291.200 ;
        RECT 199.600 290.800 200.400 292.400 ;
        RECT 202.800 291.600 203.600 292.400 ;
        RECT 206.000 292.200 206.800 292.400 ;
        RECT 205.200 291.600 206.800 292.200 ;
        RECT 207.600 291.600 208.400 292.400 ;
        RECT 209.000 292.000 209.600 295.000 ;
        RECT 210.600 294.300 211.600 294.400 ;
        RECT 214.000 294.300 214.800 294.400 ;
        RECT 210.600 293.700 214.800 294.300 ;
        RECT 210.600 293.600 211.600 293.700 ;
        RECT 214.000 293.600 214.800 293.700 ;
        RECT 210.400 292.800 211.200 293.600 ;
        RECT 215.600 292.300 216.400 295.800 ;
        RECT 217.200 293.600 218.000 295.200 ;
        RECT 220.400 293.600 221.200 294.400 ;
        RECT 220.600 293.200 221.200 293.600 ;
        RECT 220.600 292.400 221.400 293.200 ;
        RECT 222.000 292.400 222.600 295.800 ;
        RECT 223.600 292.800 224.400 294.400 ;
        RECT 228.400 293.600 229.200 294.400 ;
        RECT 228.600 293.200 229.200 293.600 ;
        RECT 228.600 292.400 229.400 293.200 ;
        RECT 230.000 292.400 230.600 295.800 ;
        RECT 231.600 292.800 232.400 294.400 ;
        RECT 236.400 293.600 237.200 294.400 ;
        RECT 236.600 293.200 237.200 293.600 ;
        RECT 236.600 292.400 237.400 293.200 ;
        RECT 238.000 292.400 238.600 295.800 ;
        RECT 243.000 295.600 243.600 295.800 ;
        RECT 243.000 295.200 244.800 295.600 ;
        RECT 243.000 295.000 247.200 295.200 ;
        RECT 244.200 294.600 247.200 295.000 ;
        RECT 246.400 294.400 247.200 294.600 ;
        RECT 239.600 292.800 240.400 294.400 ;
        RECT 242.800 292.800 243.600 294.400 ;
        RECT 244.800 293.800 245.600 294.000 ;
        RECT 244.600 293.200 245.600 293.800 ;
        RECT 244.600 292.400 245.200 293.200 ;
        RECT 218.800 292.300 219.600 292.400 ;
        RECT 202.800 291.400 203.400 291.600 ;
        RECT 201.400 290.800 203.400 291.400 ;
        RECT 205.200 291.200 206.000 291.600 ;
        RECT 185.200 289.700 188.200 290.200 ;
        RECT 185.200 289.600 186.000 289.700 ;
        RECT 186.800 289.600 188.200 289.700 ;
        RECT 188.800 289.600 189.800 290.200 ;
        RECT 193.200 289.600 194.600 290.200 ;
        RECT 187.600 288.400 188.200 289.600 ;
        RECT 187.600 287.600 188.400 288.400 ;
        RECT 189.000 282.200 189.800 289.600 ;
        RECT 193.800 284.400 194.600 289.600 ;
        RECT 193.200 283.600 194.600 284.400 ;
        RECT 193.800 282.200 194.600 283.600 ;
        RECT 198.000 282.200 198.800 290.800 ;
        RECT 201.400 290.200 202.000 290.800 ;
        RECT 207.600 290.400 208.200 291.600 ;
        RECT 209.000 291.400 209.800 292.000 ;
        RECT 215.600 291.700 219.600 292.300 ;
        RECT 209.000 291.200 213.200 291.400 ;
        RECT 209.200 290.800 213.200 291.200 ;
        RECT 207.600 290.200 208.400 290.400 ;
        RECT 199.600 282.800 200.400 290.200 ;
        RECT 201.200 283.400 202.000 290.200 ;
        RECT 202.800 289.600 206.800 290.200 ;
        RECT 207.600 289.600 209.000 290.200 ;
        RECT 202.800 282.800 203.600 289.600 ;
        RECT 199.600 282.200 203.600 282.800 ;
        RECT 206.000 282.200 206.800 289.600 ;
        RECT 208.200 282.200 209.000 289.600 ;
        RECT 212.400 282.200 213.200 290.800 ;
        RECT 214.000 288.800 214.800 290.400 ;
        RECT 215.600 282.200 216.400 291.700 ;
        RECT 218.800 290.800 219.600 291.700 ;
        RECT 222.000 291.600 222.800 292.400 ;
        RECT 225.200 292.200 226.000 292.400 ;
        RECT 224.400 291.600 226.000 292.200 ;
        RECT 222.000 291.400 222.600 291.600 ;
        RECT 220.600 290.800 222.600 291.400 ;
        RECT 224.400 291.200 225.200 291.600 ;
        RECT 226.800 290.800 227.600 292.400 ;
        RECT 230.000 291.600 230.800 292.400 ;
        RECT 233.200 292.200 234.000 292.400 ;
        RECT 232.400 291.600 234.000 292.200 ;
        RECT 230.000 291.400 230.600 291.600 ;
        RECT 228.600 290.800 230.600 291.400 ;
        RECT 232.400 291.200 233.200 291.600 ;
        RECT 234.800 290.800 235.600 292.400 ;
        RECT 238.000 291.600 238.800 292.400 ;
        RECT 241.200 292.200 242.000 292.400 ;
        RECT 240.400 291.600 242.000 292.200 ;
        RECT 244.400 291.600 245.200 292.400 ;
        RECT 238.000 291.400 238.600 291.600 ;
        RECT 236.600 290.800 238.600 291.400 ;
        RECT 240.400 291.200 241.200 291.600 ;
        RECT 246.400 291.000 247.000 294.400 ;
        RECT 247.800 292.400 248.400 295.800 ;
        RECT 249.200 295.600 250.000 297.200 ;
        RECT 247.600 292.300 248.400 292.400 ;
        RECT 249.200 292.300 250.000 292.400 ;
        RECT 247.600 291.700 250.000 292.300 ;
        RECT 247.600 291.600 248.400 291.700 ;
        RECT 249.200 291.600 250.000 291.700 ;
        RECT 250.800 292.300 251.600 299.800 ;
        RECT 255.600 295.800 256.400 299.800 ;
        RECT 257.000 296.400 257.800 297.200 ;
        RECT 254.000 292.800 254.800 294.400 ;
        RECT 252.400 292.300 253.200 292.400 ;
        RECT 250.800 292.200 253.200 292.300 ;
        RECT 255.600 292.200 256.200 295.800 ;
        RECT 257.200 295.600 258.000 296.400 ;
        RECT 258.800 295.600 259.600 297.200 ;
        RECT 260.400 294.300 261.200 299.800 ;
        RECT 262.000 296.000 262.800 299.800 ;
        RECT 265.200 296.000 266.000 299.800 ;
        RECT 262.000 295.800 266.000 296.000 ;
        RECT 266.800 298.300 267.600 299.800 ;
        RECT 270.000 298.300 270.800 298.400 ;
        RECT 266.800 297.700 270.800 298.300 ;
        RECT 266.800 295.800 267.600 297.700 ;
        RECT 270.000 297.600 270.800 297.700 ;
        RECT 276.400 296.000 277.200 299.800 ;
        RECT 262.200 295.400 265.800 295.800 ;
        RECT 262.800 294.400 263.600 294.800 ;
        RECT 266.800 294.400 267.400 295.800 ;
        RECT 276.200 295.200 277.200 296.000 ;
        RECT 262.000 294.300 263.600 294.400 ;
        RECT 260.400 293.800 263.600 294.300 ;
        RECT 260.400 293.700 262.800 293.800 ;
        RECT 257.200 292.200 258.000 292.400 ;
        RECT 250.800 291.700 254.000 292.200 ;
        RECT 220.600 290.200 221.200 290.800 ;
        RECT 228.600 290.200 229.200 290.800 ;
        RECT 236.600 290.200 237.200 290.800 ;
        RECT 244.600 290.400 247.000 291.000 ;
        RECT 218.800 282.800 219.600 290.200 ;
        RECT 220.400 283.400 221.200 290.200 ;
        RECT 222.000 289.600 226.000 290.200 ;
        RECT 222.000 282.800 222.800 289.600 ;
        RECT 218.800 282.200 222.800 282.800 ;
        RECT 225.200 282.200 226.000 289.600 ;
        RECT 226.800 282.800 227.600 290.200 ;
        RECT 228.400 283.400 229.200 290.200 ;
        RECT 230.000 289.600 234.000 290.200 ;
        RECT 230.000 282.800 230.800 289.600 ;
        RECT 226.800 282.200 230.800 282.800 ;
        RECT 233.200 282.200 234.000 289.600 ;
        RECT 234.800 282.800 235.600 290.200 ;
        RECT 236.400 283.400 237.200 290.200 ;
        RECT 238.000 289.600 242.000 290.200 ;
        RECT 238.000 282.800 238.800 289.600 ;
        RECT 234.800 282.200 238.800 282.800 ;
        RECT 241.200 282.200 242.000 289.600 ;
        RECT 244.600 286.200 245.200 290.400 ;
        RECT 247.800 290.200 248.400 291.600 ;
        RECT 244.400 282.200 245.200 286.200 ;
        RECT 247.600 282.200 248.400 290.200 ;
        RECT 250.800 282.200 251.600 291.700 ;
        RECT 252.400 291.600 254.000 291.700 ;
        RECT 255.600 291.600 258.000 292.200 ;
        RECT 253.200 291.200 254.000 291.600 ;
        RECT 257.200 290.200 257.800 291.600 ;
        RECT 252.400 289.600 256.400 290.200 ;
        RECT 252.400 282.200 253.200 289.600 ;
        RECT 255.600 282.200 256.400 289.600 ;
        RECT 257.200 282.200 258.000 290.200 ;
        RECT 260.400 282.200 261.200 293.700 ;
        RECT 262.000 293.600 262.800 293.700 ;
        RECT 265.000 293.600 267.600 294.400 ;
        RECT 263.600 291.600 264.400 293.200 ;
        RECT 265.000 290.200 265.600 293.600 ;
        RECT 276.200 290.800 277.000 295.200 ;
        RECT 278.000 294.600 278.800 299.800 ;
        RECT 284.400 296.600 285.200 299.800 ;
        RECT 286.000 297.000 286.800 299.800 ;
        RECT 287.600 297.000 288.400 299.800 ;
        RECT 289.200 297.000 290.000 299.800 ;
        RECT 290.800 297.000 291.600 299.800 ;
        RECT 294.000 297.000 294.800 299.800 ;
        RECT 297.200 297.000 298.000 299.800 ;
        RECT 298.800 297.000 299.600 299.800 ;
        RECT 300.400 297.000 301.200 299.800 ;
        RECT 282.800 295.800 285.200 296.600 ;
        RECT 302.000 296.600 302.800 299.800 ;
        RECT 282.800 295.200 283.600 295.800 ;
        RECT 277.600 294.000 278.800 294.600 ;
        RECT 281.800 294.600 283.600 295.200 ;
        RECT 287.600 295.600 288.600 296.400 ;
        RECT 291.600 295.600 293.200 296.400 ;
        RECT 294.000 295.800 298.600 296.400 ;
        RECT 302.000 295.800 304.600 296.600 ;
        RECT 294.000 295.600 294.800 295.800 ;
        RECT 277.600 292.000 278.200 294.000 ;
        RECT 281.800 293.400 282.600 294.600 ;
        RECT 278.800 292.600 282.600 293.400 ;
        RECT 287.600 292.800 288.400 295.600 ;
        RECT 294.000 294.800 294.800 295.000 ;
        RECT 290.400 294.200 294.800 294.800 ;
        RECT 290.400 294.000 291.200 294.200 ;
        RECT 295.600 293.600 296.400 295.200 ;
        RECT 297.800 293.400 298.600 295.800 ;
        RECT 303.800 295.200 304.600 295.800 ;
        RECT 303.800 294.400 306.800 295.200 ;
        RECT 308.400 293.800 309.200 299.800 ;
        RECT 311.600 295.200 312.400 299.800 ;
        RECT 314.800 295.200 315.600 299.800 ;
        RECT 318.000 295.200 318.800 299.800 ;
        RECT 321.200 295.200 322.000 299.800 ;
        RECT 290.800 292.600 294.000 293.400 ;
        RECT 297.800 292.600 299.800 293.400 ;
        RECT 300.400 293.000 309.200 293.800 ;
        RECT 284.400 292.000 285.200 292.600 ;
        RECT 302.000 292.000 302.800 292.400 ;
        RECT 305.200 292.000 306.000 292.400 ;
        RECT 307.000 292.000 307.800 292.200 ;
        RECT 277.600 291.400 278.400 292.000 ;
        RECT 284.400 291.400 307.800 292.000 ;
        RECT 266.800 290.200 267.600 290.400 ;
        RECT 264.600 289.600 265.600 290.200 ;
        RECT 266.200 289.600 267.600 290.200 ;
        RECT 276.200 290.000 277.200 290.800 ;
        RECT 264.600 282.200 265.400 289.600 ;
        RECT 266.200 288.400 266.800 289.600 ;
        RECT 266.000 287.600 266.800 288.400 ;
        RECT 276.400 282.200 277.200 290.000 ;
        RECT 277.800 289.600 278.400 291.400 ;
        RECT 277.800 289.000 286.800 289.600 ;
        RECT 277.800 287.400 278.400 289.000 ;
        RECT 286.000 288.800 286.800 289.000 ;
        RECT 289.200 289.000 297.800 289.600 ;
        RECT 289.200 288.800 290.000 289.000 ;
        RECT 281.000 287.600 283.600 288.400 ;
        RECT 277.800 286.800 280.400 287.400 ;
        RECT 279.600 282.200 280.400 286.800 ;
        RECT 282.800 282.200 283.600 287.600 ;
        RECT 284.200 286.800 288.400 287.600 ;
        RECT 286.000 282.200 286.800 285.000 ;
        RECT 287.600 282.200 288.400 285.000 ;
        RECT 289.200 282.200 290.000 285.000 ;
        RECT 290.800 282.200 291.600 288.400 ;
        RECT 294.000 287.600 296.600 288.400 ;
        RECT 297.200 288.200 297.800 289.000 ;
        RECT 298.800 289.400 299.600 289.600 ;
        RECT 298.800 289.000 304.200 289.400 ;
        RECT 298.800 288.800 305.000 289.000 ;
        RECT 303.600 288.200 305.000 288.800 ;
        RECT 297.200 287.600 303.000 288.200 ;
        RECT 306.000 288.000 307.600 288.800 ;
        RECT 306.000 287.600 306.600 288.000 ;
        RECT 294.000 282.200 294.800 287.000 ;
        RECT 297.200 282.200 298.000 287.000 ;
        RECT 302.400 286.800 306.600 287.600 ;
        RECT 308.400 287.400 309.200 293.000 ;
        RECT 310.000 294.400 312.400 295.200 ;
        RECT 313.400 294.400 315.600 295.200 ;
        RECT 316.600 294.400 318.800 295.200 ;
        RECT 320.200 294.400 322.000 295.200 ;
        RECT 325.600 298.300 326.400 299.800 ;
        RECT 327.600 298.300 328.400 298.400 ;
        RECT 325.600 297.700 328.400 298.300 ;
        RECT 310.000 291.600 310.800 294.400 ;
        RECT 313.400 293.800 314.200 294.400 ;
        RECT 316.600 293.800 317.400 294.400 ;
        RECT 320.200 293.800 321.000 294.400 ;
        RECT 325.600 294.200 326.400 297.700 ;
        RECT 327.600 297.600 328.400 297.700 ;
        RECT 330.800 295.600 331.600 297.200 ;
        RECT 311.600 293.000 314.200 293.800 ;
        RECT 315.000 293.000 317.400 293.800 ;
        RECT 318.400 293.000 321.000 293.800 ;
        RECT 313.400 291.600 314.200 293.000 ;
        RECT 316.600 291.600 317.400 293.000 ;
        RECT 320.200 291.600 321.000 293.000 ;
        RECT 324.600 293.800 326.400 294.200 ;
        RECT 332.400 294.300 333.200 299.800 ;
        RECT 334.000 296.000 334.800 299.800 ;
        RECT 337.200 296.000 338.000 299.800 ;
        RECT 334.000 295.800 338.000 296.000 ;
        RECT 338.800 295.800 339.600 299.800 ;
        RECT 340.400 295.800 341.200 299.800 ;
        RECT 342.000 296.000 342.800 299.800 ;
        RECT 345.200 296.000 346.000 299.800 ;
        RECT 342.000 295.800 346.000 296.000 ;
        RECT 348.400 297.800 349.200 299.800 ;
        RECT 354.800 298.400 355.600 299.800 ;
        RECT 354.800 297.800 355.800 298.400 ;
        RECT 334.200 295.400 337.800 295.800 ;
        RECT 334.800 294.400 335.600 294.800 ;
        RECT 338.800 294.400 339.400 295.800 ;
        RECT 340.600 294.400 341.200 295.800 ;
        RECT 342.200 295.400 345.800 295.800 ;
        RECT 344.400 294.400 345.200 294.800 ;
        RECT 348.400 294.400 349.000 297.800 ;
        RECT 355.200 297.600 355.800 297.800 ;
        RECT 358.000 298.300 358.800 299.800 ;
        RECT 362.800 298.300 363.600 298.400 ;
        RECT 358.000 297.700 363.600 298.300 ;
        RECT 358.000 297.600 359.200 297.700 ;
        RECT 362.800 297.600 363.600 297.700 ;
        RECT 350.000 296.300 350.800 297.200 ;
        RECT 355.200 297.000 359.200 297.600 ;
        RECT 353.200 296.300 355.600 296.400 ;
        RECT 350.000 295.700 355.600 296.300 ;
        RECT 350.000 295.600 350.800 295.700 ;
        RECT 353.200 295.600 355.600 295.700 ;
        RECT 334.000 294.300 335.600 294.400 ;
        RECT 332.400 293.800 335.600 294.300 ;
        RECT 324.600 293.600 326.200 293.800 ;
        RECT 332.400 293.700 334.800 293.800 ;
        RECT 310.000 290.800 312.400 291.600 ;
        RECT 313.400 290.800 315.600 291.600 ;
        RECT 316.600 290.800 318.800 291.600 ;
        RECT 320.200 290.800 322.000 291.600 ;
        RECT 307.200 286.800 309.200 287.400 ;
        RECT 298.800 282.200 299.600 285.000 ;
        RECT 300.400 282.200 301.200 285.000 ;
        RECT 303.600 282.200 304.400 286.800 ;
        RECT 307.200 286.200 307.800 286.800 ;
        RECT 306.800 285.600 307.800 286.200 ;
        RECT 306.800 282.200 307.600 285.600 ;
        RECT 311.600 282.200 312.400 290.800 ;
        RECT 314.800 282.200 315.600 290.800 ;
        RECT 318.000 282.200 318.800 290.800 ;
        RECT 321.200 282.200 322.000 290.800 ;
        RECT 324.600 290.400 325.200 293.600 ;
        RECT 326.800 291.600 328.400 292.400 ;
        RECT 324.400 289.600 325.200 290.400 ;
        RECT 329.200 289.600 330.000 291.200 ;
        RECT 324.600 287.000 325.200 289.600 ;
        RECT 326.000 288.300 326.800 289.200 ;
        RECT 330.800 288.300 331.600 288.400 ;
        RECT 326.000 287.700 331.600 288.300 ;
        RECT 326.000 287.600 326.800 287.700 ;
        RECT 330.800 287.600 331.600 287.700 ;
        RECT 324.600 286.400 328.200 287.000 ;
        RECT 324.600 286.200 325.200 286.400 ;
        RECT 324.400 282.200 325.200 286.200 ;
        RECT 327.600 286.200 328.200 286.400 ;
        RECT 327.600 282.200 328.400 286.200 ;
        RECT 332.400 282.200 333.200 293.700 ;
        RECT 334.000 293.600 334.800 293.700 ;
        RECT 337.000 293.600 339.600 294.400 ;
        RECT 340.400 293.600 343.000 294.400 ;
        RECT 344.400 294.300 346.000 294.400 ;
        RECT 348.400 294.300 349.200 294.400 ;
        RECT 351.600 294.300 352.400 294.400 ;
        RECT 344.400 293.800 347.500 294.300 ;
        RECT 345.200 293.700 347.500 293.800 ;
        RECT 345.200 293.600 346.000 293.700 ;
        RECT 335.600 291.600 336.400 293.200 ;
        RECT 337.000 290.200 337.600 293.600 ;
        RECT 342.400 292.300 343.000 293.600 ;
        RECT 346.900 292.400 347.500 293.700 ;
        RECT 348.400 293.700 352.400 294.300 ;
        RECT 348.400 293.600 349.200 293.700 ;
        RECT 351.600 293.600 352.400 293.700 ;
        RECT 353.200 294.300 354.000 294.400 ;
        RECT 354.800 294.300 356.400 294.400 ;
        RECT 353.200 293.700 356.400 294.300 ;
        RECT 353.200 293.600 354.000 293.700 ;
        RECT 354.800 293.600 356.400 293.700 ;
        RECT 338.900 291.700 343.000 292.300 ;
        RECT 338.900 290.400 339.500 291.700 ;
        RECT 338.800 290.200 339.600 290.400 ;
        RECT 336.600 289.600 337.600 290.200 ;
        RECT 338.200 289.600 339.600 290.200 ;
        RECT 340.400 290.200 341.200 290.400 ;
        RECT 342.400 290.200 343.000 291.700 ;
        RECT 346.800 290.800 347.600 292.400 ;
        RECT 348.400 290.200 349.000 293.600 ;
        RECT 356.400 291.600 358.000 292.400 ;
        RECT 358.600 290.400 359.200 297.000 ;
        RECT 364.600 296.400 365.400 297.200 ;
        RECT 361.200 296.300 362.000 296.400 ;
        RECT 364.400 296.300 365.200 296.400 ;
        RECT 361.200 295.700 365.200 296.300 ;
        RECT 361.200 295.600 362.000 295.700 ;
        RECT 364.400 295.600 365.200 295.700 ;
        RECT 366.000 295.600 366.800 299.800 ;
        RECT 364.400 292.200 365.200 292.400 ;
        RECT 366.200 292.200 366.800 295.600 ;
        RECT 367.600 292.800 368.400 294.400 ;
        RECT 369.200 292.200 370.000 292.400 ;
        RECT 364.400 291.600 366.800 292.200 ;
        RECT 368.400 291.600 370.000 292.200 ;
        RECT 340.400 289.600 341.800 290.200 ;
        RECT 342.400 289.600 343.400 290.200 ;
        RECT 336.600 282.200 337.400 289.600 ;
        RECT 338.200 288.400 338.800 289.600 ;
        RECT 338.000 287.600 338.800 288.400 ;
        RECT 341.200 288.400 341.800 289.600 ;
        RECT 341.200 287.600 342.000 288.400 ;
        RECT 342.600 282.200 343.400 289.600 ;
        RECT 347.400 289.400 349.200 290.200 ;
        RECT 358.600 289.800 362.000 290.400 ;
        RECT 364.600 290.200 365.200 291.600 ;
        RECT 368.400 291.200 369.200 291.600 ;
        RECT 361.200 289.600 362.000 289.800 ;
        RECT 347.400 282.200 348.200 289.400 ;
        RECT 351.800 288.800 355.400 289.400 ;
        RECT 351.800 288.200 352.400 288.800 ;
        RECT 351.600 282.200 352.400 288.200 ;
        RECT 354.800 288.200 355.400 288.800 ;
        RECT 356.600 289.000 360.200 289.200 ;
        RECT 361.200 289.000 361.800 289.600 ;
        RECT 356.600 288.600 360.400 289.000 ;
        RECT 356.600 288.200 357.200 288.600 ;
        RECT 354.800 282.800 355.600 288.200 ;
        RECT 356.400 283.400 357.200 288.200 ;
        RECT 358.000 282.800 358.800 288.000 ;
        RECT 359.600 283.000 360.400 288.600 ;
        RECT 361.200 283.400 362.000 289.000 ;
        RECT 354.800 282.200 358.800 282.800 ;
        RECT 359.800 282.800 360.400 283.000 ;
        RECT 362.800 283.000 363.600 289.000 ;
        RECT 362.800 282.800 363.400 283.000 ;
        RECT 359.800 282.200 363.400 282.800 ;
        RECT 364.400 282.200 365.200 290.200 ;
        RECT 366.000 289.600 370.000 290.200 ;
        RECT 366.000 282.200 366.800 289.600 ;
        RECT 369.200 282.200 370.000 289.600 ;
        RECT 370.800 282.200 371.600 299.800 ;
        RECT 372.400 293.600 373.200 295.200 ;
        RECT 374.000 282.200 374.800 299.800 ;
        RECT 375.600 295.600 376.400 297.200 ;
        RECT 377.200 295.800 378.000 299.800 ;
        RECT 378.800 296.000 379.600 299.800 ;
        RECT 382.000 296.000 382.800 299.800 ;
        RECT 385.200 297.800 386.000 299.800 ;
        RECT 378.800 295.800 382.800 296.000 ;
        RECT 377.400 294.400 378.000 295.800 ;
        RECT 379.000 295.400 382.600 295.800 ;
        RECT 383.600 295.600 384.400 297.200 ;
        RECT 381.200 294.400 382.000 294.800 ;
        RECT 385.400 294.400 386.000 297.800 ;
        RECT 389.000 296.400 389.800 299.800 ;
        RECT 389.000 295.800 390.800 296.400 ;
        RECT 393.200 296.000 394.000 299.800 ;
        RECT 396.400 296.000 397.200 299.800 ;
        RECT 393.200 295.800 397.200 296.000 ;
        RECT 398.000 295.800 398.800 299.800 ;
        RECT 400.200 296.400 401.000 299.800 ;
        RECT 407.000 298.400 407.800 299.800 ;
        RECT 406.000 297.600 407.800 298.400 ;
        RECT 407.000 296.400 407.800 297.600 ;
        RECT 409.400 296.400 410.200 297.200 ;
        RECT 400.200 295.800 402.000 296.400 ;
        RECT 377.200 293.600 379.800 294.400 ;
        RECT 381.200 293.800 382.800 294.400 ;
        RECT 382.000 293.600 382.800 293.800 ;
        RECT 385.200 293.600 386.000 294.400 ;
        RECT 377.200 290.200 378.000 290.400 ;
        RECT 379.200 290.200 379.800 293.600 ;
        RECT 380.400 291.600 381.200 293.200 ;
        RECT 383.600 292.300 384.400 292.400 ;
        RECT 385.400 292.300 386.000 293.600 ;
        RECT 383.600 291.700 386.000 292.300 ;
        RECT 383.600 291.600 384.400 291.700 ;
        RECT 385.400 290.200 386.000 291.700 ;
        RECT 386.800 292.300 387.600 292.400 ;
        RECT 390.000 292.300 390.800 295.800 ;
        RECT 393.400 295.400 397.000 295.800 ;
        RECT 391.600 293.600 392.400 295.200 ;
        RECT 394.000 294.400 394.800 294.800 ;
        RECT 398.000 294.400 398.600 295.800 ;
        RECT 393.200 293.800 394.800 294.400 ;
        RECT 393.200 293.600 394.000 293.800 ;
        RECT 396.200 293.600 398.800 294.400 ;
        RECT 399.600 294.300 400.400 294.400 ;
        RECT 401.200 294.300 402.000 295.800 ;
        RECT 406.000 295.800 407.800 296.400 ;
        RECT 399.600 293.700 402.000 294.300 ;
        RECT 399.600 293.600 400.400 293.700 ;
        RECT 386.800 291.700 390.800 292.300 ;
        RECT 386.800 290.800 387.600 291.700 ;
        RECT 377.200 289.600 378.600 290.200 ;
        RECT 379.200 289.600 380.200 290.200 ;
        RECT 378.000 288.400 378.600 289.600 ;
        RECT 378.000 287.600 378.800 288.400 ;
        RECT 379.400 282.200 380.200 289.600 ;
        RECT 385.200 289.400 387.000 290.200 ;
        RECT 386.200 282.200 387.000 289.400 ;
        RECT 388.400 288.800 389.200 290.400 ;
        RECT 390.000 282.200 390.800 291.700 ;
        RECT 394.800 291.600 395.600 293.200 ;
        RECT 396.200 292.400 396.800 293.600 ;
        RECT 396.200 291.600 397.200 292.400 ;
        RECT 396.200 290.200 396.800 291.600 ;
        RECT 398.000 290.200 398.800 290.400 ;
        RECT 395.800 289.600 396.800 290.200 ;
        RECT 397.400 289.600 398.800 290.200 ;
        RECT 395.800 282.200 396.600 289.600 ;
        RECT 397.400 288.400 398.000 289.600 ;
        RECT 399.600 288.800 400.400 290.400 ;
        RECT 397.200 287.600 398.000 288.400 ;
        RECT 401.200 282.200 402.000 293.700 ;
        RECT 402.800 294.300 403.600 295.200 ;
        RECT 404.400 294.300 405.200 295.200 ;
        RECT 402.800 293.700 405.200 294.300 ;
        RECT 402.800 293.600 403.600 293.700 ;
        RECT 404.400 293.600 405.200 293.700 ;
        RECT 406.000 282.200 406.800 295.800 ;
        RECT 409.200 295.600 410.000 296.400 ;
        RECT 410.800 295.800 411.600 299.800 ;
        RECT 409.200 292.200 410.000 292.400 ;
        RECT 411.000 292.200 411.600 295.800 ;
        RECT 415.600 295.600 416.400 297.200 ;
        RECT 412.400 294.300 413.200 294.400 ;
        RECT 417.200 294.300 418.000 299.800 ;
        RECT 420.400 297.800 421.200 299.800 ;
        RECT 418.800 295.600 419.600 297.200 ;
        RECT 420.600 294.400 421.200 297.800 ;
        RECT 412.400 293.700 418.000 294.300 ;
        RECT 412.400 292.800 413.200 293.700 ;
        RECT 414.000 292.200 414.800 292.400 ;
        RECT 409.200 291.600 411.600 292.200 ;
        RECT 413.200 291.600 414.800 292.200 ;
        RECT 407.600 288.800 408.400 290.400 ;
        RECT 409.400 290.200 410.000 291.600 ;
        RECT 413.200 291.200 414.000 291.600 ;
        RECT 409.200 282.200 410.000 290.200 ;
        RECT 410.800 289.600 414.800 290.200 ;
        RECT 410.800 282.200 411.600 289.600 ;
        RECT 414.000 282.200 414.800 289.600 ;
        RECT 417.200 282.200 418.000 293.700 ;
        RECT 420.400 293.600 421.200 294.400 ;
        RECT 418.800 292.300 419.600 292.400 ;
        RECT 420.600 292.300 421.200 293.600 ;
        RECT 430.000 292.400 430.800 299.800 ;
        RECT 433.200 295.200 434.000 299.800 ;
        RECT 437.800 295.800 439.400 299.800 ;
        RECT 443.400 296.400 444.200 299.800 ;
        RECT 443.400 295.800 445.200 296.400 ;
        RECT 431.800 294.600 434.000 295.200 ;
        RECT 418.800 291.700 421.200 292.300 ;
        RECT 418.800 291.600 419.600 291.700 ;
        RECT 420.600 290.200 421.200 291.700 ;
        RECT 422.000 290.800 422.800 292.400 ;
        RECT 430.000 290.200 430.600 292.400 ;
        RECT 431.800 291.600 432.400 294.600 ;
        RECT 436.400 292.800 437.200 294.400 ;
        RECT 438.200 292.400 438.800 295.800 ;
        RECT 439.600 294.300 440.400 294.400 ;
        RECT 444.400 294.300 445.200 295.800 ;
        RECT 447.600 295.600 448.400 297.200 ;
        RECT 439.600 293.700 445.200 294.300 ;
        RECT 439.600 293.600 440.400 293.700 ;
        RECT 439.600 293.200 440.200 293.600 ;
        RECT 439.400 292.400 440.200 293.200 ;
        RECT 434.800 292.200 435.600 292.400 ;
        RECT 434.800 291.600 436.400 292.200 ;
        RECT 438.000 291.600 438.800 292.400 ;
        RECT 431.200 290.800 432.400 291.600 ;
        RECT 435.600 291.200 436.400 291.600 ;
        RECT 438.200 291.400 438.800 291.600 ;
        RECT 438.200 290.800 440.200 291.400 ;
        RECT 441.200 290.800 442.000 292.400 ;
        RECT 431.800 290.200 432.400 290.800 ;
        RECT 439.600 290.200 440.200 290.800 ;
        RECT 420.400 289.400 422.200 290.200 ;
        RECT 421.400 282.200 422.200 289.400 ;
        RECT 430.000 282.200 430.800 290.200 ;
        RECT 431.800 289.600 434.000 290.200 ;
        RECT 433.200 282.200 434.000 289.600 ;
        RECT 434.800 289.600 438.800 290.200 ;
        RECT 434.800 282.200 435.600 289.600 ;
        RECT 438.000 282.800 438.800 289.600 ;
        RECT 439.600 283.400 440.400 290.200 ;
        RECT 441.200 282.800 442.000 290.200 ;
        RECT 442.800 288.800 443.600 290.400 ;
        RECT 438.000 282.200 442.000 282.800 ;
        RECT 444.400 282.200 445.200 293.700 ;
        RECT 446.000 294.300 446.800 295.200 ;
        RECT 447.700 294.300 448.300 295.600 ;
        RECT 446.000 293.700 448.300 294.300 ;
        RECT 446.000 293.600 446.800 293.700 ;
        RECT 449.200 282.200 450.000 299.800 ;
        RECT 452.400 296.000 453.200 299.800 ;
        RECT 452.200 295.200 453.200 296.000 ;
        RECT 452.200 290.800 453.000 295.200 ;
        RECT 454.000 294.600 454.800 299.800 ;
        RECT 460.400 296.600 461.200 299.800 ;
        RECT 462.000 297.000 462.800 299.800 ;
        RECT 463.600 297.000 464.400 299.800 ;
        RECT 465.200 297.000 466.000 299.800 ;
        RECT 466.800 297.000 467.600 299.800 ;
        RECT 470.000 297.000 470.800 299.800 ;
        RECT 473.200 297.000 474.000 299.800 ;
        RECT 474.800 297.000 475.600 299.800 ;
        RECT 476.400 297.000 477.200 299.800 ;
        RECT 458.800 295.800 461.200 296.600 ;
        RECT 478.000 296.600 478.800 299.800 ;
        RECT 458.800 295.200 459.600 295.800 ;
        RECT 453.600 294.000 454.800 294.600 ;
        RECT 457.800 294.600 459.600 295.200 ;
        RECT 463.600 295.600 464.600 296.400 ;
        RECT 467.600 295.600 469.200 296.400 ;
        RECT 470.000 295.800 474.600 296.400 ;
        RECT 478.000 295.800 480.600 296.600 ;
        RECT 470.000 295.600 470.800 295.800 ;
        RECT 453.600 292.000 454.200 294.000 ;
        RECT 457.800 293.400 458.600 294.600 ;
        RECT 454.800 292.600 458.600 293.400 ;
        RECT 463.600 292.800 464.400 295.600 ;
        RECT 470.000 294.800 470.800 295.000 ;
        RECT 466.400 294.200 470.800 294.800 ;
        RECT 466.400 294.000 467.200 294.200 ;
        RECT 471.600 293.600 472.400 295.200 ;
        RECT 473.800 293.400 474.600 295.800 ;
        RECT 479.800 295.200 480.600 295.800 ;
        RECT 479.800 294.400 482.800 295.200 ;
        RECT 484.400 293.800 485.200 299.800 ;
        RECT 486.200 296.400 487.000 297.200 ;
        RECT 486.000 295.600 486.800 296.400 ;
        RECT 487.600 295.800 488.400 299.800 ;
        RECT 492.400 299.200 496.400 299.800 ;
        RECT 492.400 295.800 493.200 299.200 ;
        RECT 494.000 295.800 494.800 298.600 ;
        RECT 495.600 296.000 496.400 299.200 ;
        RECT 498.800 296.000 499.600 299.800 ;
        RECT 495.600 295.800 499.600 296.000 ;
        RECT 466.800 292.600 470.000 293.400 ;
        RECT 473.800 292.600 475.800 293.400 ;
        RECT 476.400 293.000 485.200 293.800 ;
        RECT 460.400 292.000 461.200 292.600 ;
        RECT 478.000 292.000 478.800 292.400 ;
        RECT 479.600 292.000 480.400 292.400 ;
        RECT 483.000 292.000 483.800 292.200 ;
        RECT 453.600 291.400 454.400 292.000 ;
        RECT 460.400 291.400 483.800 292.000 ;
        RECT 452.200 290.000 453.200 290.800 ;
        RECT 452.400 282.200 453.200 290.000 ;
        RECT 453.800 289.600 454.400 291.400 ;
        RECT 453.800 289.000 462.800 289.600 ;
        RECT 453.800 287.400 454.400 289.000 ;
        RECT 462.000 288.800 462.800 289.000 ;
        RECT 465.200 289.000 473.800 289.600 ;
        RECT 465.200 288.800 466.000 289.000 ;
        RECT 457.000 287.600 459.600 288.400 ;
        RECT 453.800 286.800 456.400 287.400 ;
        RECT 455.600 282.200 456.400 286.800 ;
        RECT 458.800 282.200 459.600 287.600 ;
        RECT 460.200 286.800 464.400 287.600 ;
        RECT 462.000 282.200 462.800 285.000 ;
        RECT 463.600 282.200 464.400 285.000 ;
        RECT 465.200 282.200 466.000 285.000 ;
        RECT 466.800 282.200 467.600 288.400 ;
        RECT 470.000 287.600 472.600 288.400 ;
        RECT 473.200 288.200 473.800 289.000 ;
        RECT 474.800 289.400 475.600 289.600 ;
        RECT 474.800 289.000 480.200 289.400 ;
        RECT 474.800 288.800 481.000 289.000 ;
        RECT 479.600 288.200 481.000 288.800 ;
        RECT 473.200 287.600 479.000 288.200 ;
        RECT 482.000 288.000 483.600 288.800 ;
        RECT 482.000 287.600 482.600 288.000 ;
        RECT 470.000 282.200 470.800 287.000 ;
        RECT 473.200 282.200 474.000 287.000 ;
        RECT 478.400 286.800 482.600 287.600 ;
        RECT 484.400 287.400 485.200 293.000 ;
        RECT 486.000 292.200 486.800 292.400 ;
        RECT 487.800 292.200 488.400 295.800 ;
        RECT 494.000 294.400 494.600 295.800 ;
        RECT 495.800 295.400 499.400 295.800 ;
        RECT 498.000 294.400 498.800 294.800 ;
        RECT 489.200 292.800 490.000 294.400 ;
        RECT 492.400 292.800 493.200 294.400 ;
        RECT 494.000 293.800 496.400 294.400 ;
        RECT 498.000 293.800 499.600 294.400 ;
        RECT 495.600 293.600 496.400 293.800 ;
        RECT 498.800 293.600 499.600 293.800 ;
        RECT 490.800 292.200 491.600 292.400 ;
        RECT 486.000 291.600 488.400 292.200 ;
        RECT 490.000 291.600 491.600 292.200 ;
        RECT 494.000 291.600 494.800 293.200 ;
        RECT 495.800 292.400 496.400 293.600 ;
        RECT 495.600 291.600 496.400 292.400 ;
        RECT 497.200 292.300 498.000 293.200 ;
        RECT 498.800 292.300 499.600 292.400 ;
        RECT 497.200 291.700 499.600 292.300 ;
        RECT 497.200 291.600 498.000 291.700 ;
        RECT 498.800 291.600 499.600 291.700 ;
        RECT 486.200 290.200 486.800 291.600 ;
        RECT 490.000 291.200 490.800 291.600 ;
        RECT 495.800 290.200 496.400 291.600 ;
        RECT 483.200 286.800 485.200 287.400 ;
        RECT 474.800 282.200 475.600 285.000 ;
        RECT 476.400 282.200 477.200 285.000 ;
        RECT 479.600 282.200 480.400 286.800 ;
        RECT 483.200 286.200 483.800 286.800 ;
        RECT 482.800 285.600 483.800 286.200 ;
        RECT 482.800 282.200 483.600 285.600 ;
        RECT 486.000 282.200 486.800 290.200 ;
        RECT 487.600 289.600 491.600 290.200 ;
        RECT 487.600 282.200 488.400 289.600 ;
        RECT 490.800 282.200 491.600 289.600 ;
        RECT 495.000 282.200 497.000 290.200 ;
        RECT 500.400 282.200 501.200 299.800 ;
        RECT 505.200 297.800 506.000 299.800 ;
        RECT 503.600 295.600 504.400 297.200 ;
        RECT 502.000 293.600 502.800 295.200 ;
        RECT 505.400 294.400 506.000 297.800 ;
        RECT 509.000 298.400 509.800 299.800 ;
        RECT 509.000 297.600 510.800 298.400 ;
        RECT 509.000 296.400 509.800 297.600 ;
        RECT 509.000 295.800 510.800 296.400 ;
        RECT 505.200 293.600 506.000 294.400 ;
        RECT 505.400 290.200 506.000 293.600 ;
        RECT 506.800 290.800 507.600 292.400 ;
        RECT 505.200 289.400 507.000 290.200 ;
        RECT 506.200 288.400 507.000 289.400 ;
        RECT 508.400 288.800 509.200 290.400 ;
        RECT 506.200 287.600 507.600 288.400 ;
        RECT 506.200 282.200 507.000 287.600 ;
        RECT 510.000 282.200 510.800 295.800 ;
        RECT 513.200 296.300 514.000 296.400 ;
        RECT 514.800 296.300 515.600 299.800 ;
        RECT 513.200 295.700 515.600 296.300 ;
        RECT 513.200 295.600 514.000 295.700 ;
        RECT 514.600 295.200 515.600 295.700 ;
        RECT 511.600 293.600 512.400 295.200 ;
        RECT 514.600 290.800 515.400 295.200 ;
        RECT 516.400 294.600 517.200 299.800 ;
        RECT 522.800 296.600 523.600 299.800 ;
        RECT 524.400 297.000 525.200 299.800 ;
        RECT 526.000 297.000 526.800 299.800 ;
        RECT 527.600 297.000 528.400 299.800 ;
        RECT 529.200 297.000 530.000 299.800 ;
        RECT 532.400 297.000 533.200 299.800 ;
        RECT 535.600 297.000 536.400 299.800 ;
        RECT 537.200 297.000 538.000 299.800 ;
        RECT 538.800 297.000 539.600 299.800 ;
        RECT 521.200 295.800 523.600 296.600 ;
        RECT 540.400 296.600 541.200 299.800 ;
        RECT 521.200 295.200 522.000 295.800 ;
        RECT 516.000 294.000 517.200 294.600 ;
        RECT 520.200 294.600 522.000 295.200 ;
        RECT 526.000 295.600 527.000 296.400 ;
        RECT 530.000 295.600 531.600 296.400 ;
        RECT 532.400 295.800 537.000 296.400 ;
        RECT 540.400 295.800 543.000 296.600 ;
        RECT 532.400 295.600 533.200 295.800 ;
        RECT 516.000 292.000 516.600 294.000 ;
        RECT 520.200 293.400 521.000 294.600 ;
        RECT 517.200 292.600 521.000 293.400 ;
        RECT 526.000 292.800 526.800 295.600 ;
        RECT 532.400 294.800 533.200 295.000 ;
        RECT 528.800 294.200 533.200 294.800 ;
        RECT 528.800 294.000 529.600 294.200 ;
        RECT 534.000 293.600 534.800 295.200 ;
        RECT 536.200 293.400 537.000 295.800 ;
        RECT 542.200 295.200 543.000 295.800 ;
        RECT 542.200 294.400 545.200 295.200 ;
        RECT 546.800 293.800 547.600 299.800 ;
        RECT 529.200 292.600 532.400 293.400 ;
        RECT 536.200 292.600 538.200 293.400 ;
        RECT 538.800 293.000 547.600 293.800 ;
        RECT 522.800 292.000 523.600 292.600 ;
        RECT 540.400 292.000 541.200 292.400 ;
        RECT 545.400 292.000 546.200 292.200 ;
        RECT 516.000 291.400 516.800 292.000 ;
        RECT 522.800 291.400 546.200 292.000 ;
        RECT 514.600 290.000 515.600 290.800 ;
        RECT 514.800 282.200 515.600 290.000 ;
        RECT 516.200 289.600 516.800 291.400 ;
        RECT 516.200 289.000 525.200 289.600 ;
        RECT 516.200 287.400 516.800 289.000 ;
        RECT 524.400 288.800 525.200 289.000 ;
        RECT 527.600 289.000 536.200 289.600 ;
        RECT 527.600 288.800 528.400 289.000 ;
        RECT 519.400 287.600 522.000 288.400 ;
        RECT 516.200 286.800 518.800 287.400 ;
        RECT 518.000 282.200 518.800 286.800 ;
        RECT 521.200 282.200 522.000 287.600 ;
        RECT 522.600 286.800 526.800 287.600 ;
        RECT 524.400 282.200 525.200 285.000 ;
        RECT 526.000 282.200 526.800 285.000 ;
        RECT 527.600 282.200 528.400 285.000 ;
        RECT 529.200 282.200 530.000 288.400 ;
        RECT 532.400 287.600 535.000 288.400 ;
        RECT 535.600 288.200 536.200 289.000 ;
        RECT 537.200 289.400 538.000 289.600 ;
        RECT 537.200 289.000 542.600 289.400 ;
        RECT 537.200 288.800 543.400 289.000 ;
        RECT 542.000 288.200 543.400 288.800 ;
        RECT 535.600 287.600 541.400 288.200 ;
        RECT 544.400 288.000 546.000 288.800 ;
        RECT 544.400 287.600 545.000 288.000 ;
        RECT 532.400 282.200 533.200 287.000 ;
        RECT 535.600 282.200 536.400 287.000 ;
        RECT 540.800 286.800 545.000 287.600 ;
        RECT 546.800 287.400 547.600 293.000 ;
        RECT 545.600 286.800 547.600 287.400 ;
        RECT 537.200 282.200 538.000 285.000 ;
        RECT 538.800 282.200 539.600 285.000 ;
        RECT 542.000 282.200 542.800 286.800 ;
        RECT 545.600 286.200 546.200 286.800 ;
        RECT 545.200 285.600 546.200 286.200 ;
        RECT 545.200 282.200 546.000 285.600 ;
        RECT 2.800 272.000 3.600 279.800 ;
        RECT 6.000 275.200 6.800 279.800 ;
        RECT 2.600 271.200 3.600 272.000 ;
        RECT 4.200 274.600 6.800 275.200 ;
        RECT 4.200 273.000 4.800 274.600 ;
        RECT 9.200 274.400 10.000 279.800 ;
        RECT 12.400 277.000 13.200 279.800 ;
        RECT 14.000 277.000 14.800 279.800 ;
        RECT 15.600 277.000 16.400 279.800 ;
        RECT 10.600 274.400 14.800 275.200 ;
        RECT 7.400 273.600 10.000 274.400 ;
        RECT 17.200 273.600 18.000 279.800 ;
        RECT 20.400 275.000 21.200 279.800 ;
        RECT 23.600 275.000 24.400 279.800 ;
        RECT 25.200 277.000 26.000 279.800 ;
        RECT 26.800 277.000 27.600 279.800 ;
        RECT 30.000 275.200 30.800 279.800 ;
        RECT 33.200 276.400 34.000 279.800 ;
        RECT 33.200 275.800 34.200 276.400 ;
        RECT 33.600 275.200 34.200 275.800 ;
        RECT 28.800 274.400 33.000 275.200 ;
        RECT 33.600 274.600 35.600 275.200 ;
        RECT 20.400 273.600 23.000 274.400 ;
        RECT 23.600 273.800 29.400 274.400 ;
        RECT 32.400 274.000 33.000 274.400 ;
        RECT 12.400 273.000 13.200 273.200 ;
        RECT 4.200 272.400 13.200 273.000 ;
        RECT 15.600 273.000 16.400 273.200 ;
        RECT 23.600 273.000 24.200 273.800 ;
        RECT 30.000 273.200 31.400 273.800 ;
        RECT 32.400 273.200 34.000 274.000 ;
        RECT 15.600 272.400 24.200 273.000 ;
        RECT 25.200 273.000 31.400 273.200 ;
        RECT 25.200 272.600 30.600 273.000 ;
        RECT 25.200 272.400 26.000 272.600 ;
        RECT 2.600 266.800 3.400 271.200 ;
        RECT 4.200 270.600 4.800 272.400 ;
        RECT 4.000 270.000 4.800 270.600 ;
        RECT 10.800 270.000 34.200 270.600 ;
        RECT 4.000 268.000 4.600 270.000 ;
        RECT 10.800 269.400 11.600 270.000 ;
        RECT 28.400 269.600 29.200 270.000 ;
        RECT 30.000 269.600 30.800 270.000 ;
        RECT 33.400 269.800 34.200 270.000 ;
        RECT 5.200 268.600 9.000 269.400 ;
        RECT 4.000 267.400 5.200 268.000 ;
        RECT 2.600 266.000 3.600 266.800 ;
        RECT 2.800 262.200 3.600 266.000 ;
        RECT 4.400 262.200 5.200 267.400 ;
        RECT 8.200 267.400 9.000 268.600 ;
        RECT 8.200 266.800 10.000 267.400 ;
        RECT 9.200 266.200 10.000 266.800 ;
        RECT 14.000 266.400 14.800 269.200 ;
        RECT 17.200 268.600 20.400 269.400 ;
        RECT 24.200 268.600 26.200 269.400 ;
        RECT 34.800 269.000 35.600 274.600 ;
        RECT 39.000 274.400 41.000 279.800 ;
        RECT 38.000 273.600 41.000 274.400 ;
        RECT 39.000 271.800 41.000 273.600 ;
        RECT 16.800 267.800 17.600 268.000 ;
        RECT 16.800 267.200 21.200 267.800 ;
        RECT 20.400 267.000 21.200 267.200 ;
        RECT 22.000 266.800 22.800 268.400 ;
        RECT 9.200 265.400 11.600 266.200 ;
        RECT 14.000 265.600 15.000 266.400 ;
        RECT 18.000 265.600 19.600 266.400 ;
        RECT 20.400 266.200 21.200 266.400 ;
        RECT 24.200 266.200 25.000 268.600 ;
        RECT 26.800 268.200 35.600 269.000 ;
        RECT 38.000 268.800 38.800 270.400 ;
        RECT 39.600 268.400 40.200 271.800 ;
        RECT 44.400 271.600 45.200 273.200 ;
        RECT 41.200 268.800 42.000 270.400 ;
        RECT 30.200 266.800 33.200 267.600 ;
        RECT 30.200 266.200 31.000 266.800 ;
        RECT 20.400 265.600 25.000 266.200 ;
        RECT 10.800 262.200 11.600 265.400 ;
        RECT 28.400 265.400 31.000 266.200 ;
        RECT 12.400 262.200 13.200 265.000 ;
        RECT 14.000 262.200 14.800 265.000 ;
        RECT 15.600 262.200 16.400 265.000 ;
        RECT 17.200 262.200 18.000 265.000 ;
        RECT 20.400 262.200 21.200 265.000 ;
        RECT 23.600 262.200 24.400 265.000 ;
        RECT 25.200 262.200 26.000 265.000 ;
        RECT 26.800 262.200 27.600 265.000 ;
        RECT 28.400 262.200 29.200 265.400 ;
        RECT 34.800 262.200 35.600 268.200 ;
        RECT 36.400 268.200 37.200 268.400 ;
        RECT 39.600 268.200 40.400 268.400 ;
        RECT 36.400 267.600 38.000 268.200 ;
        RECT 39.600 267.600 42.000 268.200 ;
        RECT 42.800 267.600 43.600 269.200 ;
        RECT 37.200 267.200 38.000 267.600 ;
        RECT 36.600 266.200 40.200 266.600 ;
        RECT 41.400 266.200 42.000 267.600 ;
        RECT 46.000 266.200 46.800 279.800 ;
        RECT 49.800 272.600 50.600 279.800 ;
        RECT 55.600 275.800 56.400 279.800 ;
        RECT 49.800 271.800 51.600 272.600 ;
        RECT 49.200 269.600 50.000 271.200 ;
        RECT 50.800 270.300 51.400 271.800 ;
        RECT 55.800 271.600 56.400 275.800 ;
        RECT 58.800 272.300 59.600 279.800 ;
        RECT 60.400 272.300 61.200 273.200 ;
        RECT 58.800 271.800 61.200 272.300 ;
        RECT 58.900 271.700 61.200 271.800 ;
        RECT 55.800 271.000 58.200 271.600 ;
        RECT 52.400 270.300 53.200 270.400 ;
        RECT 50.800 269.700 53.200 270.300 ;
        RECT 50.800 268.400 51.400 269.700 ;
        RECT 52.400 269.600 53.200 269.700 ;
        RECT 55.600 269.600 56.400 270.400 ;
        RECT 47.600 266.800 48.400 268.400 ;
        RECT 50.800 267.600 51.600 268.400 ;
        RECT 54.000 267.600 54.800 269.200 ;
        RECT 55.800 268.800 56.400 269.600 ;
        RECT 55.800 268.200 56.800 268.800 ;
        RECT 56.000 268.000 56.800 268.200 ;
        RECT 57.600 267.600 58.200 271.000 ;
        RECT 59.000 270.400 59.600 271.700 ;
        RECT 60.400 271.600 61.200 271.700 ;
        RECT 58.800 269.600 59.600 270.400 ;
        RECT 36.400 266.000 40.400 266.200 ;
        RECT 36.400 262.200 37.200 266.000 ;
        RECT 39.600 262.800 40.400 266.000 ;
        RECT 41.200 263.400 42.000 266.200 ;
        RECT 42.800 262.800 43.600 266.200 ;
        RECT 39.600 262.200 43.600 262.800 ;
        RECT 45.000 265.600 46.800 266.200 ;
        RECT 45.000 264.400 45.800 265.600 ;
        RECT 45.000 263.600 46.800 264.400 ;
        RECT 50.800 264.200 51.400 267.600 ;
        RECT 57.600 267.400 58.400 267.600 ;
        RECT 55.400 267.000 58.400 267.400 ;
        RECT 54.200 266.800 58.400 267.000 ;
        RECT 54.200 266.400 56.000 266.800 ;
        RECT 52.400 264.800 53.200 266.400 ;
        RECT 54.200 266.200 54.800 266.400 ;
        RECT 59.000 266.200 59.600 269.600 ;
        RECT 62.000 266.200 62.800 279.800 ;
        RECT 65.200 271.600 66.000 273.200 ;
        RECT 63.600 266.800 64.400 268.400 ;
        RECT 66.800 266.200 67.600 279.800 ;
        RECT 70.800 273.600 71.600 274.400 ;
        RECT 70.800 272.400 71.400 273.600 ;
        RECT 72.200 272.400 73.000 279.800 ;
        RECT 79.000 272.600 79.800 279.800 ;
        RECT 82.800 275.800 83.600 279.800 ;
        RECT 70.000 271.800 71.400 272.400 ;
        RECT 72.000 271.800 73.000 272.400 ;
        RECT 78.000 271.800 79.800 272.600 ;
        RECT 70.000 271.600 70.800 271.800 ;
        RECT 72.000 268.400 72.600 271.800 ;
        RECT 73.200 270.300 74.000 270.400 ;
        RECT 78.200 270.300 78.800 271.800 ;
        RECT 83.000 271.600 83.600 275.800 ;
        RECT 86.000 271.800 86.800 279.800 ;
        RECT 73.200 269.700 78.800 270.300 ;
        RECT 73.200 268.800 74.000 269.700 ;
        RECT 78.200 268.400 78.800 269.700 ;
        RECT 79.600 269.600 80.400 271.200 ;
        RECT 83.000 271.000 85.400 271.600 ;
        RECT 82.800 269.600 83.600 270.400 ;
        RECT 68.400 266.800 69.200 268.400 ;
        RECT 70.000 267.600 72.600 268.400 ;
        RECT 74.800 268.200 75.600 268.400 ;
        RECT 74.000 267.600 75.600 268.200 ;
        RECT 78.000 267.600 78.800 268.400 ;
        RECT 79.700 268.300 80.300 269.600 ;
        RECT 81.200 268.300 82.000 269.200 ;
        RECT 79.700 267.700 82.000 268.300 ;
        RECT 83.000 268.800 83.600 269.600 ;
        RECT 83.000 268.200 84.000 268.800 ;
        RECT 83.200 268.000 84.000 268.200 ;
        RECT 81.200 267.600 82.000 267.700 ;
        RECT 84.800 267.600 85.400 271.000 ;
        RECT 86.200 270.400 86.800 271.800 ;
        RECT 86.000 269.600 86.800 270.400 ;
        RECT 70.200 266.200 70.800 267.600 ;
        RECT 74.000 267.200 74.800 267.600 ;
        RECT 71.800 266.200 75.400 266.600 ;
        RECT 45.000 262.200 45.800 263.600 ;
        RECT 50.800 262.200 51.600 264.200 ;
        RECT 54.000 262.200 54.800 266.200 ;
        RECT 58.200 265.200 59.600 266.200 ;
        RECT 61.000 265.600 62.800 266.200 ;
        RECT 65.800 265.600 67.600 266.200 ;
        RECT 58.200 262.200 59.000 265.200 ;
        RECT 61.000 264.400 61.800 265.600 ;
        RECT 61.000 263.600 62.800 264.400 ;
        RECT 61.000 262.200 61.800 263.600 ;
        RECT 65.800 262.200 66.600 265.600 ;
        RECT 70.000 262.200 70.800 266.200 ;
        RECT 71.600 266.000 75.600 266.200 ;
        RECT 71.600 262.200 72.400 266.000 ;
        RECT 74.800 262.200 75.600 266.000 ;
        RECT 76.400 264.800 77.200 266.400 ;
        RECT 78.200 264.200 78.800 267.600 ;
        RECT 84.800 267.400 85.600 267.600 ;
        RECT 82.600 267.000 85.600 267.400 ;
        RECT 81.400 266.800 85.600 267.000 ;
        RECT 81.400 266.400 83.200 266.800 ;
        RECT 81.400 266.200 82.000 266.400 ;
        RECT 86.200 266.200 86.800 269.600 ;
        RECT 78.000 262.200 78.800 264.200 ;
        RECT 81.200 262.200 82.000 266.200 ;
        RECT 85.400 265.200 86.800 266.200 ;
        RECT 85.400 262.200 86.200 265.200 ;
        RECT 87.600 264.800 88.400 266.400 ;
        RECT 89.200 262.200 90.000 279.800 ;
        RECT 92.400 276.400 93.200 279.800 ;
        RECT 92.200 275.800 93.200 276.400 ;
        RECT 92.200 275.200 92.800 275.800 ;
        RECT 95.600 275.200 96.400 279.800 ;
        RECT 98.800 277.000 99.600 279.800 ;
        RECT 100.400 277.000 101.200 279.800 ;
        RECT 90.800 274.600 92.800 275.200 ;
        RECT 90.800 269.000 91.600 274.600 ;
        RECT 93.400 274.400 97.600 275.200 ;
        RECT 102.000 275.000 102.800 279.800 ;
        RECT 105.200 275.000 106.000 279.800 ;
        RECT 93.400 274.000 94.000 274.400 ;
        RECT 92.400 273.200 94.000 274.000 ;
        RECT 97.000 273.800 102.800 274.400 ;
        RECT 95.000 273.200 96.400 273.800 ;
        RECT 95.000 273.000 101.200 273.200 ;
        RECT 95.800 272.600 101.200 273.000 ;
        RECT 100.400 272.400 101.200 272.600 ;
        RECT 102.200 273.000 102.800 273.800 ;
        RECT 103.400 273.600 106.000 274.400 ;
        RECT 108.400 273.600 109.200 279.800 ;
        RECT 110.000 277.000 110.800 279.800 ;
        RECT 111.600 277.000 112.400 279.800 ;
        RECT 113.200 277.000 114.000 279.800 ;
        RECT 111.600 274.400 115.800 275.200 ;
        RECT 116.400 274.400 117.200 279.800 ;
        RECT 119.600 275.200 120.400 279.800 ;
        RECT 119.600 274.600 122.200 275.200 ;
        RECT 116.400 273.600 119.000 274.400 ;
        RECT 110.000 273.000 110.800 273.200 ;
        RECT 102.200 272.400 110.800 273.000 ;
        RECT 113.200 273.000 114.000 273.200 ;
        RECT 121.600 273.000 122.200 274.600 ;
        RECT 113.200 272.400 122.200 273.000 ;
        RECT 121.600 270.600 122.200 272.400 ;
        RECT 122.800 272.000 123.600 279.800 ;
        RECT 132.400 279.200 136.400 279.800 ;
        RECT 122.800 271.200 123.800 272.000 ;
        RECT 132.400 271.800 133.200 279.200 ;
        RECT 134.000 271.800 134.800 278.600 ;
        RECT 135.600 272.400 136.400 279.200 ;
        RECT 138.800 272.400 139.600 279.800 ;
        RECT 135.600 271.800 139.600 272.400 ;
        RECT 134.200 271.200 134.800 271.800 ;
        RECT 140.400 271.600 141.200 273.200 ;
        RECT 92.200 270.000 115.600 270.600 ;
        RECT 121.600 270.000 122.400 270.600 ;
        RECT 92.200 269.800 93.000 270.000 ;
        RECT 97.200 269.600 98.000 270.000 ;
        RECT 103.600 269.600 104.400 270.000 ;
        RECT 114.800 269.400 115.600 270.000 ;
        RECT 90.800 268.200 99.600 269.000 ;
        RECT 100.200 268.600 102.200 269.400 ;
        RECT 106.000 268.600 109.200 269.400 ;
        RECT 90.800 262.200 91.600 268.200 ;
        RECT 93.200 266.800 96.200 267.600 ;
        RECT 95.400 266.200 96.200 266.800 ;
        RECT 101.400 266.200 102.200 268.600 ;
        RECT 103.600 266.800 104.400 268.400 ;
        RECT 108.800 267.800 109.600 268.000 ;
        RECT 105.200 267.200 109.600 267.800 ;
        RECT 105.200 267.000 106.000 267.200 ;
        RECT 111.600 266.400 112.400 269.200 ;
        RECT 117.400 268.600 121.200 269.400 ;
        RECT 117.400 267.400 118.200 268.600 ;
        RECT 121.800 268.000 122.400 270.000 ;
        RECT 105.200 266.200 106.000 266.400 ;
        RECT 95.400 265.400 98.000 266.200 ;
        RECT 101.400 265.600 106.000 266.200 ;
        RECT 106.800 265.600 108.400 266.400 ;
        RECT 111.400 265.600 112.400 266.400 ;
        RECT 116.400 266.800 118.200 267.400 ;
        RECT 121.200 267.400 122.400 268.000 ;
        RECT 123.000 268.300 123.800 271.200 ;
        RECT 132.400 269.600 133.200 271.200 ;
        RECT 134.200 270.600 136.200 271.200 ;
        RECT 135.600 270.400 136.200 270.600 ;
        RECT 138.000 270.400 138.800 270.800 ;
        RECT 135.600 269.600 136.400 270.400 ;
        RECT 138.000 269.800 139.600 270.400 ;
        RECT 138.800 269.600 139.600 269.800 ;
        RECT 134.200 268.800 135.000 269.600 ;
        RECT 134.200 268.400 134.800 268.800 ;
        RECT 132.400 268.300 133.200 268.400 ;
        RECT 123.000 267.700 133.200 268.300 ;
        RECT 116.400 266.200 117.200 266.800 ;
        RECT 97.200 262.200 98.000 265.400 ;
        RECT 114.800 265.400 117.200 266.200 ;
        RECT 98.800 262.200 99.600 265.000 ;
        RECT 100.400 262.200 101.200 265.000 ;
        RECT 102.000 262.200 102.800 265.000 ;
        RECT 105.200 262.200 106.000 265.000 ;
        RECT 108.400 262.200 109.200 265.000 ;
        RECT 110.000 262.200 110.800 265.000 ;
        RECT 111.600 262.200 112.400 265.000 ;
        RECT 113.200 262.200 114.000 265.000 ;
        RECT 114.800 262.200 115.600 265.400 ;
        RECT 121.200 262.200 122.000 267.400 ;
        RECT 123.000 266.800 123.800 267.700 ;
        RECT 132.400 267.600 133.200 267.700 ;
        RECT 134.000 267.600 134.800 268.400 ;
        RECT 122.800 266.000 123.800 266.800 ;
        RECT 135.600 266.200 136.200 269.600 ;
        RECT 137.200 268.300 138.000 269.200 ;
        RECT 138.800 268.300 139.600 268.400 ;
        RECT 137.200 267.700 139.600 268.300 ;
        RECT 137.200 267.600 138.000 267.700 ;
        RECT 138.800 267.600 139.600 267.700 ;
        RECT 142.000 266.200 142.800 279.800 ;
        RECT 146.000 273.600 146.800 274.400 ;
        RECT 146.000 272.400 146.600 273.600 ;
        RECT 147.400 272.400 148.200 279.800 ;
        RECT 145.200 271.800 146.600 272.400 ;
        RECT 147.200 271.800 148.200 272.400 ;
        RECT 151.600 271.800 152.400 279.800 ;
        RECT 153.200 272.400 154.000 279.800 ;
        RECT 156.400 272.400 157.200 279.800 ;
        RECT 160.600 272.600 161.400 279.800 ;
        RECT 153.200 271.800 157.200 272.400 ;
        RECT 159.600 271.800 161.400 272.600 ;
        RECT 145.200 271.600 146.000 271.800 ;
        RECT 147.200 268.400 147.800 271.800 ;
        RECT 151.800 270.400 152.400 271.800 ;
        RECT 155.600 270.400 156.400 270.800 ;
        RECT 148.400 268.800 149.200 270.400 ;
        RECT 151.600 269.800 154.000 270.400 ;
        RECT 155.600 269.800 157.200 270.400 ;
        RECT 151.600 269.600 152.400 269.800 ;
        RECT 143.600 268.300 144.400 268.400 ;
        RECT 145.200 268.300 147.800 268.400 ;
        RECT 143.600 267.700 147.800 268.300 ;
        RECT 150.000 268.300 150.800 268.400 ;
        RECT 153.400 268.300 154.000 269.800 ;
        RECT 156.400 269.600 157.200 269.800 ;
        RECT 150.000 268.200 154.000 268.300 ;
        RECT 143.600 266.800 144.400 267.700 ;
        RECT 145.200 267.600 147.800 267.700 ;
        RECT 149.200 267.700 154.000 268.200 ;
        RECT 149.200 267.600 150.800 267.700 ;
        RECT 145.400 266.200 146.000 267.600 ;
        RECT 149.200 267.200 150.000 267.600 ;
        RECT 147.000 266.200 150.600 266.600 ;
        RECT 122.800 262.200 123.600 266.000 ;
        RECT 135.000 262.200 136.600 266.200 ;
        RECT 141.000 265.600 142.800 266.200 ;
        RECT 141.000 262.200 141.800 265.600 ;
        RECT 145.200 262.200 146.000 266.200 ;
        RECT 146.800 266.000 150.800 266.200 ;
        RECT 146.800 262.200 147.600 266.000 ;
        RECT 150.000 262.200 150.800 266.000 ;
        RECT 151.600 265.600 152.400 266.400 ;
        RECT 153.400 266.200 154.000 267.700 ;
        RECT 154.800 267.600 155.600 269.200 ;
        RECT 159.800 268.400 160.400 271.800 ;
        RECT 161.200 269.600 162.000 271.200 ;
        RECT 159.600 268.300 160.400 268.400 ;
        RECT 162.800 268.300 163.600 268.400 ;
        RECT 159.600 267.700 163.600 268.300 ;
        RECT 159.600 267.600 160.400 267.700 ;
        RECT 151.800 264.800 152.600 265.600 ;
        RECT 153.200 262.200 154.000 266.200 ;
        RECT 158.000 264.800 158.800 266.400 ;
        RECT 159.800 264.200 160.400 267.600 ;
        RECT 162.800 266.800 163.600 267.700 ;
        RECT 164.400 266.200 165.200 279.800 ;
        RECT 167.600 274.300 168.400 274.400 ;
        RECT 169.200 274.300 170.000 279.800 ;
        RECT 174.000 275.800 174.800 279.800 ;
        RECT 174.200 275.600 174.800 275.800 ;
        RECT 177.200 275.800 178.000 279.800 ;
        RECT 177.200 275.600 177.800 275.800 ;
        RECT 174.200 275.000 177.800 275.600 ;
        RECT 174.000 274.300 174.800 274.400 ;
        RECT 167.600 273.700 170.000 274.300 ;
        RECT 167.600 273.600 168.400 273.700 ;
        RECT 166.000 271.600 166.800 273.200 ;
        RECT 167.600 266.800 168.400 268.400 ;
        RECT 169.200 266.200 170.000 273.700 ;
        RECT 170.800 273.700 174.800 274.300 ;
        RECT 170.800 271.600 171.600 273.700 ;
        RECT 174.000 273.600 174.800 273.700 ;
        RECT 175.600 272.800 176.400 274.400 ;
        RECT 177.200 272.400 177.800 275.000 ;
        RECT 172.400 270.800 173.200 272.400 ;
        RECT 177.200 271.600 178.000 272.400 ;
        RECT 178.800 271.600 179.600 273.200 ;
        RECT 174.000 269.600 175.600 270.400 ;
        RECT 177.200 268.400 177.800 271.600 ;
        RECT 176.200 268.200 177.800 268.400 ;
        RECT 176.000 267.800 177.800 268.200 ;
        RECT 164.400 265.600 166.200 266.200 ;
        RECT 169.200 265.600 171.000 266.200 ;
        RECT 159.600 262.200 160.400 264.200 ;
        RECT 165.400 264.400 166.200 265.600 ;
        RECT 165.400 263.600 166.800 264.400 ;
        RECT 165.400 262.200 166.200 263.600 ;
        RECT 170.200 262.200 171.000 265.600 ;
        RECT 176.000 262.200 176.800 267.800 ;
        RECT 180.400 266.200 181.200 279.800 ;
        RECT 185.800 274.400 186.600 279.800 ;
        RECT 184.400 273.600 185.200 274.400 ;
        RECT 185.800 273.600 187.600 274.400 ;
        RECT 190.800 273.600 191.600 274.400 ;
        RECT 184.400 272.400 185.000 273.600 ;
        RECT 185.800 272.400 186.600 273.600 ;
        RECT 190.800 272.400 191.400 273.600 ;
        RECT 192.200 272.400 193.000 279.800 ;
        RECT 198.000 275.800 198.800 279.800 ;
        RECT 198.200 275.600 198.800 275.800 ;
        RECT 201.200 275.800 202.000 279.800 ;
        RECT 201.200 275.600 201.800 275.800 ;
        RECT 198.200 275.000 201.800 275.600 ;
        RECT 199.600 272.800 200.400 274.400 ;
        RECT 201.200 272.400 201.800 275.000 ;
        RECT 183.600 271.800 185.000 272.400 ;
        RECT 185.600 271.800 186.600 272.400 ;
        RECT 190.000 271.800 191.400 272.400 ;
        RECT 192.000 271.800 193.000 272.400 ;
        RECT 183.600 271.600 184.400 271.800 ;
        RECT 185.600 268.400 186.200 271.800 ;
        RECT 190.000 271.600 190.800 271.800 ;
        RECT 186.800 270.300 187.600 270.400 ;
        RECT 188.400 270.300 189.200 270.400 ;
        RECT 186.800 269.700 189.200 270.300 ;
        RECT 186.800 268.800 187.600 269.700 ;
        RECT 188.400 269.600 189.200 269.700 ;
        RECT 192.000 268.400 192.600 271.800 ;
        RECT 196.400 270.800 197.200 272.400 ;
        RECT 201.200 271.600 202.000 272.400 ;
        RECT 193.200 268.800 194.000 270.400 ;
        RECT 198.000 269.600 199.600 270.400 ;
        RECT 201.200 268.400 201.800 271.600 ;
        RECT 182.000 266.800 182.800 268.400 ;
        RECT 183.600 267.600 186.200 268.400 ;
        RECT 188.400 268.200 189.200 268.400 ;
        RECT 187.600 267.600 189.200 268.200 ;
        RECT 190.000 267.600 192.600 268.400 ;
        RECT 194.800 268.200 195.600 268.400 ;
        RECT 200.200 268.200 201.800 268.400 ;
        RECT 194.000 267.600 195.600 268.200 ;
        RECT 200.000 267.800 201.800 268.200 ;
        RECT 183.800 266.200 184.400 267.600 ;
        RECT 187.600 267.200 188.400 267.600 ;
        RECT 185.400 266.200 189.000 266.600 ;
        RECT 190.200 266.200 190.800 267.600 ;
        RECT 194.000 267.200 194.800 267.600 ;
        RECT 191.800 266.200 195.400 266.600 ;
        RECT 179.400 265.600 181.200 266.200 ;
        RECT 179.400 264.400 180.200 265.600 ;
        RECT 178.800 263.600 180.200 264.400 ;
        RECT 179.400 262.200 180.200 263.600 ;
        RECT 183.600 262.200 184.400 266.200 ;
        RECT 185.200 266.000 189.200 266.200 ;
        RECT 185.200 262.200 186.000 266.000 ;
        RECT 188.400 262.200 189.200 266.000 ;
        RECT 190.000 262.200 190.800 266.200 ;
        RECT 191.600 266.000 195.600 266.200 ;
        RECT 191.600 262.200 192.400 266.000 ;
        RECT 194.800 262.200 195.600 266.000 ;
        RECT 200.000 262.200 200.800 267.800 ;
        RECT 202.800 262.200 203.600 279.800 ;
        RECT 208.600 278.400 209.400 279.800 ;
        RECT 207.600 277.600 209.400 278.400 ;
        RECT 208.600 272.600 209.400 277.600 ;
        RECT 211.400 274.400 212.200 279.800 ;
        RECT 210.800 273.600 212.200 274.400 ;
        RECT 207.600 271.800 209.400 272.600 ;
        RECT 211.400 272.600 212.200 273.600 ;
        RECT 211.400 271.800 213.200 272.600 ;
        RECT 218.200 272.400 219.000 279.800 ;
        RECT 219.600 273.600 220.400 274.400 ;
        RECT 219.800 272.400 220.400 273.600 ;
        RECT 218.200 271.800 219.200 272.400 ;
        RECT 219.800 271.800 221.200 272.400 ;
        RECT 207.800 268.400 208.400 271.800 ;
        RECT 209.200 269.600 210.000 271.200 ;
        RECT 210.800 269.600 211.600 271.200 ;
        RECT 207.600 267.600 208.400 268.400 ;
        RECT 204.400 264.800 205.200 266.400 ;
        RECT 206.000 264.800 206.800 266.400 ;
        RECT 207.800 264.200 208.400 267.600 ;
        RECT 207.600 262.200 208.400 264.200 ;
        RECT 212.400 268.400 213.000 271.800 ;
        RECT 214.000 270.300 214.800 270.400 ;
        RECT 217.200 270.300 218.000 270.400 ;
        RECT 214.000 269.700 218.000 270.300 ;
        RECT 214.000 269.600 214.800 269.700 ;
        RECT 217.200 268.800 218.000 269.700 ;
        RECT 218.600 268.400 219.200 271.800 ;
        RECT 220.400 271.600 221.200 271.800 ;
        RECT 223.600 270.300 224.400 279.800 ;
        RECT 225.200 271.600 226.000 273.200 ;
        RECT 226.800 270.300 227.600 270.400 ;
        RECT 223.600 269.700 227.600 270.300 ;
        RECT 212.400 267.600 213.200 268.400 ;
        RECT 215.600 268.200 216.400 268.400 ;
        RECT 218.600 268.300 221.200 268.400 ;
        RECT 222.000 268.300 222.800 268.400 ;
        RECT 215.600 267.600 217.200 268.200 ;
        RECT 218.600 267.700 222.800 268.300 ;
        RECT 218.600 267.600 221.200 267.700 ;
        RECT 212.400 264.200 213.000 267.600 ;
        RECT 216.400 267.200 217.200 267.600 ;
        RECT 214.000 264.800 214.800 266.400 ;
        RECT 215.800 266.200 219.400 266.600 ;
        RECT 220.400 266.200 221.000 267.600 ;
        RECT 222.000 266.800 222.800 267.700 ;
        RECT 223.600 266.200 224.400 269.700 ;
        RECT 226.800 269.600 227.600 269.700 ;
        RECT 228.400 268.300 229.200 279.800 ;
        RECT 232.600 272.400 233.400 279.800 ;
        RECT 236.400 279.200 240.400 279.800 ;
        RECT 234.000 273.600 234.800 274.400 ;
        RECT 234.200 272.400 234.800 273.600 ;
        RECT 232.600 271.800 233.600 272.400 ;
        RECT 234.200 271.800 235.600 272.400 ;
        RECT 236.400 271.800 237.200 279.200 ;
        RECT 238.000 271.800 238.800 278.600 ;
        RECT 239.600 272.400 240.400 279.200 ;
        RECT 242.800 272.400 243.600 279.800 ;
        RECT 239.600 271.800 243.600 272.400 ;
        RECT 231.600 268.800 232.400 270.400 ;
        RECT 233.000 268.400 233.600 271.800 ;
        RECT 234.800 271.600 235.600 271.800 ;
        RECT 238.200 271.200 238.800 271.800 ;
        RECT 236.400 269.600 237.200 271.200 ;
        RECT 238.200 270.600 240.200 271.200 ;
        RECT 239.600 270.400 240.200 270.600 ;
        RECT 242.000 270.400 242.800 270.800 ;
        RECT 239.600 269.600 240.400 270.400 ;
        RECT 242.000 269.800 243.600 270.400 ;
        RECT 242.800 269.600 243.600 269.800 ;
        RECT 238.200 268.800 239.000 269.600 ;
        RECT 238.200 268.400 238.800 268.800 ;
        RECT 230.000 268.300 230.800 268.400 ;
        RECT 228.400 268.200 230.800 268.300 ;
        RECT 228.400 267.700 231.600 268.200 ;
        RECT 215.600 266.000 219.600 266.200 ;
        RECT 212.400 262.200 213.200 264.200 ;
        RECT 215.600 262.200 216.400 266.000 ;
        RECT 218.800 262.200 219.600 266.000 ;
        RECT 220.400 262.200 221.200 266.200 ;
        RECT 223.600 265.600 225.400 266.200 ;
        RECT 224.600 262.200 225.400 265.600 ;
        RECT 226.800 264.800 227.600 266.400 ;
        RECT 228.400 262.200 229.200 267.700 ;
        RECT 230.000 267.600 231.600 267.700 ;
        RECT 233.000 267.600 235.600 268.400 ;
        RECT 238.000 267.600 238.800 268.400 ;
        RECT 230.800 267.200 231.600 267.600 ;
        RECT 230.200 266.200 233.800 266.600 ;
        RECT 234.800 266.200 235.400 267.600 ;
        RECT 239.600 266.200 240.200 269.600 ;
        RECT 241.200 267.600 242.000 269.200 ;
        RECT 246.000 268.300 246.800 279.800 ;
        RECT 250.200 272.400 251.000 279.800 ;
        RECT 251.600 273.600 252.400 274.400 ;
        RECT 251.800 272.400 252.400 273.600 ;
        RECT 250.200 271.800 251.200 272.400 ;
        RECT 251.800 271.800 253.200 272.400 ;
        RECT 256.600 271.800 258.600 279.800 ;
        RECT 270.000 272.000 270.800 279.800 ;
        RECT 273.200 275.200 274.000 279.800 ;
        RECT 249.200 268.800 250.000 270.400 ;
        RECT 250.600 268.400 251.200 271.800 ;
        RECT 252.400 271.600 253.200 271.800 ;
        RECT 247.600 268.300 248.400 268.400 ;
        RECT 246.000 268.200 248.400 268.300 ;
        RECT 246.000 267.700 249.200 268.200 ;
        RECT 230.000 266.000 234.000 266.200 ;
        RECT 230.000 262.200 230.800 266.000 ;
        RECT 233.200 262.200 234.000 266.000 ;
        RECT 234.800 262.200 235.600 266.200 ;
        RECT 239.000 262.200 240.600 266.200 ;
        RECT 244.400 264.800 245.200 266.400 ;
        RECT 246.000 262.200 246.800 267.700 ;
        RECT 247.600 267.600 249.200 267.700 ;
        RECT 250.600 267.600 253.200 268.400 ;
        RECT 254.000 267.600 254.800 269.200 ;
        RECT 255.600 268.800 256.400 270.400 ;
        RECT 257.400 268.400 258.000 271.800 ;
        RECT 269.800 271.200 270.800 272.000 ;
        RECT 271.400 274.600 274.000 275.200 ;
        RECT 271.400 273.000 272.000 274.600 ;
        RECT 276.400 274.400 277.200 279.800 ;
        RECT 279.600 277.000 280.400 279.800 ;
        RECT 281.200 277.000 282.000 279.800 ;
        RECT 282.800 277.000 283.600 279.800 ;
        RECT 277.800 274.400 282.000 275.200 ;
        RECT 274.600 273.600 277.200 274.400 ;
        RECT 284.400 273.600 285.200 279.800 ;
        RECT 287.600 275.000 288.400 279.800 ;
        RECT 290.800 275.000 291.600 279.800 ;
        RECT 292.400 277.000 293.200 279.800 ;
        RECT 294.000 277.000 294.800 279.800 ;
        RECT 297.200 275.200 298.000 279.800 ;
        RECT 300.400 276.400 301.200 279.800 ;
        RECT 305.200 276.400 306.000 279.800 ;
        RECT 300.400 275.800 301.400 276.400 ;
        RECT 300.800 275.200 301.400 275.800 ;
        RECT 305.000 275.800 306.000 276.400 ;
        RECT 305.000 275.200 305.600 275.800 ;
        RECT 308.400 275.200 309.200 279.800 ;
        RECT 311.600 277.000 312.400 279.800 ;
        RECT 313.200 277.000 314.000 279.800 ;
        RECT 296.000 274.400 300.200 275.200 ;
        RECT 300.800 274.600 302.800 275.200 ;
        RECT 287.600 273.600 290.200 274.400 ;
        RECT 290.800 273.800 296.600 274.400 ;
        RECT 299.600 274.000 300.200 274.400 ;
        RECT 279.600 273.000 280.400 273.200 ;
        RECT 271.400 272.400 280.400 273.000 ;
        RECT 282.800 273.000 283.600 273.200 ;
        RECT 290.800 273.000 291.400 273.800 ;
        RECT 297.200 273.200 298.600 273.800 ;
        RECT 299.600 273.200 301.200 274.000 ;
        RECT 282.800 272.400 291.400 273.000 ;
        RECT 292.400 273.000 298.600 273.200 ;
        RECT 292.400 272.600 297.800 273.000 ;
        RECT 292.400 272.400 293.200 272.600 ;
        RECT 258.800 268.800 259.600 270.400 ;
        RECT 257.200 268.200 258.000 268.400 ;
        RECT 260.400 268.200 261.200 268.400 ;
        RECT 255.600 267.600 258.000 268.200 ;
        RECT 259.600 267.600 261.200 268.200 ;
        RECT 248.400 267.200 249.200 267.600 ;
        RECT 247.800 266.200 251.400 266.600 ;
        RECT 252.400 266.200 253.000 267.600 ;
        RECT 255.600 266.200 256.200 267.600 ;
        RECT 259.600 267.200 260.400 267.600 ;
        RECT 269.800 266.800 270.600 271.200 ;
        RECT 271.400 270.600 272.000 272.400 ;
        RECT 295.400 271.800 296.400 272.000 ;
        RECT 298.800 271.800 299.600 272.400 ;
        RECT 272.600 271.200 299.600 271.800 ;
        RECT 272.600 271.000 273.400 271.200 ;
        RECT 271.200 270.000 272.000 270.600 ;
        RECT 271.200 268.000 271.800 270.000 ;
        RECT 272.400 268.600 276.200 269.400 ;
        RECT 271.200 267.400 272.400 268.000 ;
        RECT 257.400 266.200 261.000 266.600 ;
        RECT 247.600 266.000 251.600 266.200 ;
        RECT 247.600 262.200 248.400 266.000 ;
        RECT 250.800 262.200 251.600 266.000 ;
        RECT 252.400 262.200 253.200 266.200 ;
        RECT 254.000 262.800 254.800 266.200 ;
        RECT 255.600 263.400 256.400 266.200 ;
        RECT 257.200 266.000 261.200 266.200 ;
        RECT 269.800 266.000 270.800 266.800 ;
        RECT 257.200 262.800 258.000 266.000 ;
        RECT 254.000 262.200 258.000 262.800 ;
        RECT 260.400 262.200 261.200 266.000 ;
        RECT 270.000 262.200 270.800 266.000 ;
        RECT 271.600 262.200 272.400 267.400 ;
        RECT 275.400 267.400 276.200 268.600 ;
        RECT 275.400 266.800 277.200 267.400 ;
        RECT 276.400 266.200 277.200 266.800 ;
        RECT 281.200 266.400 282.000 269.200 ;
        RECT 284.400 268.600 287.600 269.400 ;
        RECT 291.400 268.600 293.400 269.400 ;
        RECT 302.000 269.000 302.800 274.600 ;
        RECT 284.000 267.800 284.800 268.000 ;
        RECT 284.000 267.200 288.400 267.800 ;
        RECT 287.600 267.000 288.400 267.200 ;
        RECT 289.200 266.800 290.000 268.400 ;
        RECT 276.400 265.400 278.800 266.200 ;
        RECT 281.200 265.600 282.200 266.400 ;
        RECT 285.200 265.600 286.800 266.400 ;
        RECT 287.600 266.200 288.400 266.400 ;
        RECT 291.400 266.200 292.200 268.600 ;
        RECT 294.000 268.200 302.800 269.000 ;
        RECT 297.400 266.800 300.400 267.600 ;
        RECT 297.400 266.200 298.200 266.800 ;
        RECT 287.600 265.600 292.200 266.200 ;
        RECT 278.000 262.200 278.800 265.400 ;
        RECT 295.600 265.400 298.200 266.200 ;
        RECT 279.600 262.200 280.400 265.000 ;
        RECT 281.200 262.200 282.000 265.000 ;
        RECT 282.800 262.200 283.600 265.000 ;
        RECT 284.400 262.200 285.200 265.000 ;
        RECT 287.600 262.200 288.400 265.000 ;
        RECT 290.800 262.200 291.600 265.000 ;
        RECT 292.400 262.200 293.200 265.000 ;
        RECT 294.000 262.200 294.800 265.000 ;
        RECT 295.600 262.200 296.400 265.400 ;
        RECT 302.000 262.200 302.800 268.200 ;
        RECT 303.600 274.600 305.600 275.200 ;
        RECT 303.600 269.000 304.400 274.600 ;
        RECT 306.200 274.400 310.400 275.200 ;
        RECT 314.800 275.000 315.600 279.800 ;
        RECT 318.000 275.000 318.800 279.800 ;
        RECT 306.200 274.000 306.800 274.400 ;
        RECT 305.200 273.200 306.800 274.000 ;
        RECT 309.800 273.800 315.600 274.400 ;
        RECT 307.800 273.200 309.200 273.800 ;
        RECT 307.800 273.000 314.000 273.200 ;
        RECT 308.600 272.600 314.000 273.000 ;
        RECT 313.200 272.400 314.000 272.600 ;
        RECT 315.000 273.000 315.600 273.800 ;
        RECT 316.200 273.600 318.800 274.400 ;
        RECT 321.200 273.600 322.000 279.800 ;
        RECT 322.800 277.000 323.600 279.800 ;
        RECT 324.400 277.000 325.200 279.800 ;
        RECT 326.000 277.000 326.800 279.800 ;
        RECT 324.400 274.400 328.600 275.200 ;
        RECT 329.200 274.400 330.000 279.800 ;
        RECT 332.400 275.200 333.200 279.800 ;
        RECT 332.400 274.600 335.000 275.200 ;
        RECT 329.200 273.600 331.800 274.400 ;
        RECT 322.800 273.000 323.600 273.200 ;
        RECT 315.000 272.400 323.600 273.000 ;
        RECT 326.000 273.000 326.800 273.200 ;
        RECT 334.400 273.000 335.000 274.600 ;
        RECT 326.000 272.400 335.000 273.000 ;
        RECT 306.800 271.800 307.600 272.400 ;
        RECT 310.200 271.800 311.000 272.000 ;
        RECT 306.800 271.200 333.800 271.800 ;
        RECT 333.000 271.000 333.800 271.200 ;
        RECT 334.400 270.600 335.000 272.400 ;
        RECT 335.600 272.000 336.400 279.800 ;
        RECT 335.600 271.200 336.600 272.000 ;
        RECT 334.400 270.000 335.200 270.600 ;
        RECT 303.600 268.200 312.400 269.000 ;
        RECT 313.000 268.600 315.000 269.400 ;
        RECT 318.800 268.600 322.000 269.400 ;
        RECT 303.600 262.200 304.400 268.200 ;
        RECT 306.000 266.800 309.000 267.600 ;
        RECT 308.200 266.200 309.000 266.800 ;
        RECT 314.200 266.200 315.000 268.600 ;
        RECT 316.400 266.800 317.200 268.400 ;
        RECT 321.600 267.800 322.400 268.000 ;
        RECT 318.000 267.200 322.400 267.800 ;
        RECT 318.000 267.000 318.800 267.200 ;
        RECT 324.400 266.400 325.200 269.200 ;
        RECT 330.200 268.600 334.000 269.400 ;
        RECT 330.200 267.400 331.000 268.600 ;
        RECT 334.600 268.000 335.200 270.000 ;
        RECT 318.000 266.200 318.800 266.400 ;
        RECT 308.200 265.400 310.800 266.200 ;
        RECT 314.200 265.600 318.800 266.200 ;
        RECT 319.600 265.600 321.200 266.400 ;
        RECT 324.200 265.600 325.200 266.400 ;
        RECT 329.200 266.800 331.000 267.400 ;
        RECT 334.000 267.400 335.200 268.000 ;
        RECT 329.200 266.200 330.000 266.800 ;
        RECT 310.000 262.200 310.800 265.400 ;
        RECT 327.600 265.400 330.000 266.200 ;
        RECT 311.600 262.200 312.400 265.000 ;
        RECT 313.200 262.200 314.000 265.000 ;
        RECT 314.800 262.200 315.600 265.000 ;
        RECT 318.000 262.200 318.800 265.000 ;
        RECT 321.200 262.200 322.000 265.000 ;
        RECT 322.800 262.200 323.600 265.000 ;
        RECT 324.400 262.200 325.200 265.000 ;
        RECT 326.000 262.200 326.800 265.000 ;
        RECT 327.600 262.200 328.400 265.400 ;
        RECT 334.000 262.200 334.800 267.400 ;
        RECT 335.800 266.800 336.600 271.200 ;
        RECT 335.600 266.300 336.600 266.800 ;
        RECT 338.800 266.300 339.600 266.400 ;
        RECT 335.600 265.700 339.600 266.300 ;
        RECT 335.600 262.200 336.400 265.700 ;
        RECT 338.800 264.800 339.600 265.700 ;
        RECT 340.400 262.200 341.200 279.800 ;
        RECT 343.600 275.800 344.400 279.800 ;
        RECT 343.800 271.600 344.400 275.800 ;
        RECT 346.800 271.800 347.600 279.800 ;
        RECT 350.000 276.400 350.800 279.800 ;
        RECT 349.800 275.800 350.800 276.400 ;
        RECT 349.800 275.200 350.400 275.800 ;
        RECT 353.200 275.200 354.000 279.800 ;
        RECT 356.400 277.000 357.200 279.800 ;
        RECT 358.000 277.000 358.800 279.800 ;
        RECT 343.800 271.000 346.200 271.600 ;
        RECT 343.600 269.600 344.400 270.400 ;
        RECT 342.000 267.600 342.800 269.200 ;
        RECT 343.800 268.800 344.400 269.600 ;
        RECT 343.800 268.200 344.800 268.800 ;
        RECT 344.000 268.000 344.800 268.200 ;
        RECT 345.600 267.600 346.200 271.000 ;
        RECT 347.000 270.400 347.600 271.800 ;
        RECT 346.800 269.600 347.600 270.400 ;
        RECT 345.600 267.400 346.400 267.600 ;
        RECT 343.400 267.000 346.400 267.400 ;
        RECT 342.200 266.800 346.400 267.000 ;
        RECT 342.200 266.400 344.000 266.800 ;
        RECT 342.200 266.200 342.800 266.400 ;
        RECT 347.000 266.200 347.600 269.600 ;
        RECT 342.000 262.200 342.800 266.200 ;
        RECT 346.200 265.200 347.600 266.200 ;
        RECT 348.400 274.600 350.400 275.200 ;
        RECT 348.400 269.000 349.200 274.600 ;
        RECT 351.000 274.400 355.200 275.200 ;
        RECT 359.600 275.000 360.400 279.800 ;
        RECT 362.800 275.000 363.600 279.800 ;
        RECT 351.000 274.000 351.600 274.400 ;
        RECT 350.000 273.200 351.600 274.000 ;
        RECT 354.600 273.800 360.400 274.400 ;
        RECT 352.600 273.200 354.000 273.800 ;
        RECT 352.600 273.000 358.800 273.200 ;
        RECT 353.400 272.600 358.800 273.000 ;
        RECT 358.000 272.400 358.800 272.600 ;
        RECT 359.800 273.000 360.400 273.800 ;
        RECT 361.000 273.600 363.600 274.400 ;
        RECT 366.000 273.600 366.800 279.800 ;
        RECT 367.600 277.000 368.400 279.800 ;
        RECT 369.200 277.000 370.000 279.800 ;
        RECT 370.800 277.000 371.600 279.800 ;
        RECT 369.200 274.400 373.400 275.200 ;
        RECT 374.000 274.400 374.800 279.800 ;
        RECT 377.200 275.200 378.000 279.800 ;
        RECT 377.200 274.600 379.800 275.200 ;
        RECT 374.000 273.600 376.600 274.400 ;
        RECT 367.600 273.000 368.400 273.200 ;
        RECT 359.800 272.400 368.400 273.000 ;
        RECT 370.800 273.000 371.600 273.200 ;
        RECT 379.200 273.000 379.800 274.600 ;
        RECT 370.800 272.400 379.800 273.000 ;
        RECT 351.600 271.800 352.400 272.400 ;
        RECT 354.800 271.800 355.800 272.000 ;
        RECT 351.600 271.200 378.600 271.800 ;
        RECT 377.800 271.000 378.600 271.200 ;
        RECT 379.200 270.600 379.800 272.400 ;
        RECT 380.400 272.000 381.200 279.800 ;
        RECT 385.200 276.400 386.000 279.800 ;
        RECT 385.000 275.800 386.000 276.400 ;
        RECT 385.000 275.200 385.600 275.800 ;
        RECT 388.400 275.200 389.200 279.800 ;
        RECT 391.600 277.000 392.400 279.800 ;
        RECT 393.200 277.000 394.000 279.800 ;
        RECT 383.600 274.600 385.600 275.200 ;
        RECT 380.400 271.200 381.400 272.000 ;
        RECT 379.200 270.000 380.000 270.600 ;
        RECT 348.400 268.200 357.200 269.000 ;
        RECT 357.800 268.600 359.800 269.400 ;
        RECT 363.600 268.600 366.800 269.400 ;
        RECT 346.200 264.400 347.000 265.200 ;
        RECT 346.200 263.600 347.600 264.400 ;
        RECT 346.200 262.200 347.000 263.600 ;
        RECT 348.400 262.200 349.200 268.200 ;
        RECT 350.800 266.800 353.800 267.600 ;
        RECT 353.000 266.200 353.800 266.800 ;
        RECT 359.000 266.200 359.800 268.600 ;
        RECT 361.200 266.800 362.000 268.400 ;
        RECT 366.400 267.800 367.200 268.000 ;
        RECT 362.800 267.200 367.200 267.800 ;
        RECT 362.800 267.000 363.600 267.200 ;
        RECT 369.200 266.400 370.000 269.200 ;
        RECT 375.000 268.600 378.800 269.400 ;
        RECT 375.000 267.400 375.800 268.600 ;
        RECT 379.400 268.000 380.000 270.000 ;
        RECT 362.800 266.200 363.600 266.400 ;
        RECT 353.000 265.400 355.600 266.200 ;
        RECT 359.000 265.600 363.600 266.200 ;
        RECT 364.400 265.600 366.000 266.400 ;
        RECT 369.000 265.600 370.000 266.400 ;
        RECT 374.000 266.800 375.800 267.400 ;
        RECT 378.800 267.400 380.000 268.000 ;
        RECT 374.000 266.200 374.800 266.800 ;
        RECT 354.800 262.200 355.600 265.400 ;
        RECT 372.400 265.400 374.800 266.200 ;
        RECT 356.400 262.200 357.200 265.000 ;
        RECT 358.000 262.200 358.800 265.000 ;
        RECT 359.600 262.200 360.400 265.000 ;
        RECT 362.800 262.200 363.600 265.000 ;
        RECT 366.000 262.200 366.800 265.000 ;
        RECT 367.600 262.200 368.400 265.000 ;
        RECT 369.200 262.200 370.000 265.000 ;
        RECT 370.800 262.200 371.600 265.000 ;
        RECT 372.400 262.200 373.200 265.400 ;
        RECT 378.800 262.200 379.600 267.400 ;
        RECT 380.600 266.800 381.400 271.200 ;
        RECT 380.400 266.000 381.400 266.800 ;
        RECT 383.600 269.000 384.400 274.600 ;
        RECT 386.200 274.400 390.400 275.200 ;
        RECT 394.800 275.000 395.600 279.800 ;
        RECT 398.000 275.000 398.800 279.800 ;
        RECT 386.200 274.000 386.800 274.400 ;
        RECT 385.200 273.200 386.800 274.000 ;
        RECT 389.800 273.800 395.600 274.400 ;
        RECT 387.800 273.200 389.200 273.800 ;
        RECT 387.800 273.000 394.000 273.200 ;
        RECT 388.600 272.600 394.000 273.000 ;
        RECT 393.200 272.400 394.000 272.600 ;
        RECT 395.000 273.000 395.600 273.800 ;
        RECT 396.200 273.600 398.800 274.400 ;
        RECT 401.200 273.600 402.000 279.800 ;
        RECT 402.800 277.000 403.600 279.800 ;
        RECT 404.400 277.000 405.200 279.800 ;
        RECT 406.000 277.000 406.800 279.800 ;
        RECT 404.400 274.400 408.600 275.200 ;
        RECT 409.200 274.400 410.000 279.800 ;
        RECT 412.400 275.200 413.200 279.800 ;
        RECT 412.400 274.600 415.000 275.200 ;
        RECT 409.200 273.600 411.800 274.400 ;
        RECT 402.800 273.000 403.600 273.200 ;
        RECT 395.000 272.400 403.600 273.000 ;
        RECT 406.000 273.000 406.800 273.200 ;
        RECT 414.400 273.000 415.000 274.600 ;
        RECT 406.000 272.400 415.000 273.000 ;
        RECT 414.400 270.600 415.000 272.400 ;
        RECT 415.600 274.300 416.400 279.800 ;
        RECT 417.200 274.300 418.000 274.400 ;
        RECT 415.600 273.700 418.000 274.300 ;
        RECT 415.600 272.000 416.400 273.700 ;
        RECT 417.200 273.600 418.000 273.700 ;
        RECT 419.400 272.600 420.200 279.800 ;
        RECT 415.600 271.200 416.600 272.000 ;
        RECT 419.400 271.800 421.200 272.600 ;
        RECT 385.000 270.000 408.400 270.600 ;
        RECT 414.400 270.000 415.200 270.600 ;
        RECT 385.000 269.800 385.800 270.000 ;
        RECT 386.800 269.600 387.600 270.000 ;
        RECT 390.000 269.600 390.800 270.000 ;
        RECT 407.600 269.400 408.400 270.000 ;
        RECT 383.600 268.200 392.400 269.000 ;
        RECT 393.000 268.600 395.000 269.400 ;
        RECT 398.800 268.600 402.000 269.400 ;
        RECT 380.400 262.200 381.200 266.000 ;
        RECT 383.600 262.200 384.400 268.200 ;
        RECT 386.000 266.800 389.000 267.600 ;
        RECT 388.200 266.200 389.000 266.800 ;
        RECT 394.200 266.200 395.000 268.600 ;
        RECT 396.400 266.800 397.200 268.400 ;
        RECT 401.600 267.800 402.400 268.000 ;
        RECT 398.000 267.200 402.400 267.800 ;
        RECT 398.000 267.000 398.800 267.200 ;
        RECT 404.400 266.400 405.200 269.200 ;
        RECT 410.200 268.600 414.000 269.400 ;
        RECT 410.200 267.400 411.000 268.600 ;
        RECT 414.600 268.000 415.200 270.000 ;
        RECT 398.000 266.200 398.800 266.400 ;
        RECT 388.200 265.400 390.800 266.200 ;
        RECT 394.200 265.600 398.800 266.200 ;
        RECT 399.600 265.600 401.200 266.400 ;
        RECT 404.200 265.600 405.200 266.400 ;
        RECT 409.200 266.800 411.000 267.400 ;
        RECT 414.000 267.400 415.200 268.000 ;
        RECT 409.200 266.200 410.000 266.800 ;
        RECT 390.000 262.200 390.800 265.400 ;
        RECT 407.600 265.400 410.000 266.200 ;
        RECT 391.600 262.200 392.400 265.000 ;
        RECT 393.200 262.200 394.000 265.000 ;
        RECT 394.800 262.200 395.600 265.000 ;
        RECT 398.000 262.200 398.800 265.000 ;
        RECT 401.200 262.200 402.000 265.000 ;
        RECT 402.800 262.200 403.600 265.000 ;
        RECT 404.400 262.200 405.200 265.000 ;
        RECT 406.000 262.200 406.800 265.000 ;
        RECT 407.600 262.200 408.400 265.400 ;
        RECT 414.000 262.200 414.800 267.400 ;
        RECT 415.800 266.800 416.600 271.200 ;
        RECT 418.800 269.600 419.600 271.200 ;
        RECT 415.600 266.000 416.600 266.800 ;
        RECT 420.400 268.400 421.000 271.800 ;
        RECT 420.400 267.600 421.200 268.400 ;
        RECT 431.600 268.300 432.400 279.800 ;
        RECT 435.800 272.400 436.600 279.800 ;
        RECT 437.200 273.600 438.000 274.400 ;
        RECT 437.400 272.400 438.000 273.600 ;
        RECT 442.200 272.400 443.000 279.800 ;
        RECT 443.600 273.600 444.400 274.400 ;
        RECT 443.800 272.400 444.400 273.600 ;
        RECT 435.800 271.800 436.800 272.400 ;
        RECT 437.400 271.800 438.800 272.400 ;
        RECT 442.200 271.800 443.200 272.400 ;
        RECT 443.800 271.800 445.200 272.400 ;
        RECT 434.800 268.800 435.600 270.400 ;
        RECT 436.200 268.400 436.800 271.800 ;
        RECT 438.000 271.600 438.800 271.800 ;
        RECT 442.600 270.400 443.200 271.800 ;
        RECT 444.400 271.600 445.200 271.800 ;
        RECT 441.200 268.800 442.000 270.400 ;
        RECT 442.600 269.600 443.600 270.400 ;
        RECT 442.600 268.400 443.200 269.600 ;
        RECT 433.200 268.300 434.000 268.400 ;
        RECT 431.600 268.200 434.000 268.300 ;
        RECT 431.600 267.700 434.800 268.200 ;
        RECT 415.600 262.200 416.400 266.000 ;
        RECT 420.400 264.400 421.000 267.600 ;
        RECT 422.000 264.800 422.800 266.400 ;
        RECT 430.000 264.800 430.800 266.400 ;
        RECT 420.400 262.200 421.200 264.400 ;
        RECT 431.600 262.200 432.400 267.700 ;
        RECT 433.200 267.600 434.800 267.700 ;
        RECT 436.200 267.600 438.800 268.400 ;
        RECT 439.600 268.200 440.400 268.400 ;
        RECT 439.600 267.600 441.200 268.200 ;
        RECT 442.600 267.600 445.200 268.400 ;
        RECT 434.000 267.200 434.800 267.600 ;
        RECT 433.400 266.200 437.000 266.600 ;
        RECT 438.000 266.200 438.600 267.600 ;
        RECT 440.400 267.200 441.200 267.600 ;
        RECT 439.800 266.200 443.400 266.600 ;
        RECT 444.400 266.200 445.000 267.600 ;
        RECT 433.200 266.000 437.200 266.200 ;
        RECT 433.200 262.200 434.000 266.000 ;
        RECT 436.400 262.200 437.200 266.000 ;
        RECT 438.000 262.200 438.800 266.200 ;
        RECT 439.600 266.000 443.600 266.200 ;
        RECT 439.600 262.200 440.400 266.000 ;
        RECT 442.800 262.200 443.600 266.000 ;
        RECT 444.400 262.200 445.200 266.200 ;
        RECT 446.000 264.800 446.800 266.400 ;
        RECT 447.600 262.200 448.400 279.800 ;
        RECT 449.200 262.200 450.000 279.800 ;
        RECT 454.000 272.000 454.800 279.800 ;
        RECT 457.200 275.200 458.000 279.800 ;
        RECT 453.800 271.200 454.800 272.000 ;
        RECT 455.400 274.600 458.000 275.200 ;
        RECT 455.400 273.000 456.000 274.600 ;
        RECT 460.400 274.400 461.200 279.800 ;
        RECT 463.600 277.000 464.400 279.800 ;
        RECT 465.200 277.000 466.000 279.800 ;
        RECT 466.800 277.000 467.600 279.800 ;
        RECT 461.800 274.400 466.000 275.200 ;
        RECT 458.600 273.600 461.200 274.400 ;
        RECT 468.400 273.600 469.200 279.800 ;
        RECT 471.600 275.000 472.400 279.800 ;
        RECT 474.800 275.000 475.600 279.800 ;
        RECT 476.400 277.000 477.200 279.800 ;
        RECT 478.000 277.000 478.800 279.800 ;
        RECT 481.200 275.200 482.000 279.800 ;
        RECT 484.400 276.400 485.200 279.800 ;
        RECT 484.400 275.800 485.400 276.400 ;
        RECT 484.800 275.200 485.400 275.800 ;
        RECT 480.000 274.400 484.200 275.200 ;
        RECT 484.800 274.600 486.800 275.200 ;
        RECT 471.600 273.600 474.200 274.400 ;
        RECT 474.800 273.800 480.600 274.400 ;
        RECT 483.600 274.000 484.200 274.400 ;
        RECT 463.600 273.000 464.400 273.200 ;
        RECT 455.400 272.400 464.400 273.000 ;
        RECT 466.800 273.000 467.600 273.200 ;
        RECT 474.800 273.000 475.400 273.800 ;
        RECT 481.200 273.200 482.600 273.800 ;
        RECT 483.600 273.200 485.200 274.000 ;
        RECT 466.800 272.400 475.400 273.000 ;
        RECT 476.400 273.000 482.600 273.200 ;
        RECT 476.400 272.600 481.800 273.000 ;
        RECT 476.400 272.400 477.200 272.600 ;
        RECT 453.800 266.800 454.600 271.200 ;
        RECT 455.400 270.600 456.000 272.400 ;
        RECT 455.200 270.000 456.000 270.600 ;
        RECT 462.000 270.000 485.400 270.600 ;
        RECT 455.200 268.000 455.800 270.000 ;
        RECT 462.000 269.400 462.800 270.000 ;
        RECT 479.600 269.600 480.400 270.000 ;
        RECT 482.800 269.600 483.600 270.000 ;
        RECT 484.600 269.800 485.400 270.000 ;
        RECT 456.400 268.600 460.200 269.400 ;
        RECT 455.200 267.400 456.400 268.000 ;
        RECT 450.800 266.300 451.600 266.400 ;
        RECT 453.800 266.300 454.800 266.800 ;
        RECT 450.800 265.700 454.800 266.300 ;
        RECT 450.800 264.800 451.600 265.700 ;
        RECT 454.000 262.200 454.800 265.700 ;
        RECT 455.600 262.200 456.400 267.400 ;
        RECT 459.400 267.400 460.200 268.600 ;
        RECT 459.400 266.800 461.200 267.400 ;
        RECT 460.400 266.200 461.200 266.800 ;
        RECT 465.200 266.400 466.000 269.200 ;
        RECT 468.400 268.600 471.600 269.400 ;
        RECT 475.400 268.600 477.400 269.400 ;
        RECT 486.000 269.000 486.800 274.600 ;
        RECT 489.200 272.000 490.000 279.800 ;
        RECT 492.400 275.200 493.200 279.800 ;
        RECT 468.000 267.800 468.800 268.000 ;
        RECT 468.000 267.200 472.400 267.800 ;
        RECT 471.600 267.000 472.400 267.200 ;
        RECT 473.200 266.800 474.000 268.400 ;
        RECT 460.400 265.400 462.800 266.200 ;
        RECT 465.200 265.600 466.200 266.400 ;
        RECT 469.200 265.600 470.800 266.400 ;
        RECT 471.600 266.200 472.400 266.400 ;
        RECT 475.400 266.200 476.200 268.600 ;
        RECT 478.000 268.200 486.800 269.000 ;
        RECT 481.400 266.800 484.400 267.600 ;
        RECT 481.400 266.200 482.200 266.800 ;
        RECT 471.600 265.600 476.200 266.200 ;
        RECT 462.000 262.200 462.800 265.400 ;
        RECT 479.600 265.400 482.200 266.200 ;
        RECT 463.600 262.200 464.400 265.000 ;
        RECT 465.200 262.200 466.000 265.000 ;
        RECT 466.800 262.200 467.600 265.000 ;
        RECT 468.400 262.200 469.200 265.000 ;
        RECT 471.600 262.200 472.400 265.000 ;
        RECT 474.800 262.200 475.600 265.000 ;
        RECT 476.400 262.200 477.200 265.000 ;
        RECT 478.000 262.200 478.800 265.000 ;
        RECT 479.600 262.200 480.400 265.400 ;
        RECT 486.000 262.200 486.800 268.200 ;
        RECT 489.000 271.200 490.000 272.000 ;
        RECT 490.600 274.600 493.200 275.200 ;
        RECT 490.600 273.000 491.200 274.600 ;
        RECT 495.600 274.400 496.400 279.800 ;
        RECT 498.800 277.000 499.600 279.800 ;
        RECT 500.400 277.000 501.200 279.800 ;
        RECT 502.000 277.000 502.800 279.800 ;
        RECT 497.000 274.400 501.200 275.200 ;
        RECT 493.800 273.600 496.400 274.400 ;
        RECT 503.600 273.600 504.400 279.800 ;
        RECT 506.800 275.000 507.600 279.800 ;
        RECT 510.000 275.000 510.800 279.800 ;
        RECT 511.600 277.000 512.400 279.800 ;
        RECT 513.200 277.000 514.000 279.800 ;
        RECT 516.400 275.200 517.200 279.800 ;
        RECT 519.600 276.400 520.400 279.800 ;
        RECT 519.600 275.800 520.600 276.400 ;
        RECT 520.000 275.200 520.600 275.800 ;
        RECT 515.200 274.400 519.400 275.200 ;
        RECT 520.000 274.600 522.000 275.200 ;
        RECT 506.800 273.600 509.400 274.400 ;
        RECT 510.000 273.800 515.800 274.400 ;
        RECT 518.800 274.000 519.400 274.400 ;
        RECT 498.800 273.000 499.600 273.200 ;
        RECT 490.600 272.400 499.600 273.000 ;
        RECT 502.000 273.000 502.800 273.200 ;
        RECT 510.000 273.000 510.600 273.800 ;
        RECT 516.400 273.200 517.800 273.800 ;
        RECT 518.800 273.200 520.400 274.000 ;
        RECT 502.000 272.400 510.600 273.000 ;
        RECT 511.600 273.000 517.800 273.200 ;
        RECT 511.600 272.600 517.000 273.000 ;
        RECT 511.600 272.400 512.400 272.600 ;
        RECT 489.000 266.800 489.800 271.200 ;
        RECT 490.600 270.600 491.200 272.400 ;
        RECT 490.400 270.000 491.200 270.600 ;
        RECT 497.200 270.000 520.600 270.600 ;
        RECT 490.400 268.000 491.000 270.000 ;
        RECT 497.200 269.400 498.000 270.000 ;
        RECT 514.800 269.600 515.600 270.000 ;
        RECT 519.600 269.800 520.600 270.000 ;
        RECT 519.600 269.600 520.400 269.800 ;
        RECT 491.600 268.600 495.400 269.400 ;
        RECT 490.400 267.400 491.600 268.000 ;
        RECT 489.000 266.000 490.000 266.800 ;
        RECT 489.200 262.200 490.000 266.000 ;
        RECT 490.800 262.200 491.600 267.400 ;
        RECT 494.600 267.400 495.400 268.600 ;
        RECT 494.600 266.800 496.400 267.400 ;
        RECT 495.600 266.200 496.400 266.800 ;
        RECT 500.400 266.400 501.200 269.200 ;
        RECT 503.600 268.600 506.800 269.400 ;
        RECT 510.600 268.600 512.600 269.400 ;
        RECT 521.200 269.000 522.000 274.600 ;
        RECT 503.200 267.800 504.000 268.000 ;
        RECT 503.200 267.200 507.600 267.800 ;
        RECT 506.800 267.000 507.600 267.200 ;
        RECT 508.400 266.800 509.200 268.400 ;
        RECT 495.600 265.400 498.000 266.200 ;
        RECT 500.400 265.600 501.400 266.400 ;
        RECT 504.400 265.600 506.000 266.400 ;
        RECT 506.800 266.200 507.600 266.400 ;
        RECT 510.600 266.200 511.400 268.600 ;
        RECT 513.200 268.200 522.000 269.000 ;
        RECT 516.600 266.800 519.600 267.600 ;
        RECT 516.600 266.200 517.400 266.800 ;
        RECT 506.800 265.600 511.400 266.200 ;
        RECT 497.200 262.200 498.000 265.400 ;
        RECT 514.800 265.400 517.400 266.200 ;
        RECT 498.800 262.200 499.600 265.000 ;
        RECT 500.400 262.200 501.200 265.000 ;
        RECT 502.000 262.200 502.800 265.000 ;
        RECT 503.600 262.200 504.400 265.000 ;
        RECT 506.800 262.200 507.600 265.000 ;
        RECT 510.000 262.200 510.800 265.000 ;
        RECT 511.600 262.200 512.400 265.000 ;
        RECT 513.200 262.200 514.000 265.000 ;
        RECT 514.800 262.200 515.600 265.400 ;
        RECT 521.200 262.200 522.000 268.200 ;
        RECT 522.800 262.200 523.600 279.800 ;
        RECT 526.000 271.400 526.800 279.800 ;
        RECT 530.400 276.400 531.200 279.800 ;
        RECT 529.200 275.800 531.200 276.400 ;
        RECT 534.800 275.800 535.600 279.800 ;
        RECT 539.000 275.800 540.200 279.800 ;
        RECT 529.200 275.000 530.000 275.800 ;
        RECT 534.800 275.200 535.400 275.800 ;
        RECT 532.600 274.600 536.200 275.200 ;
        RECT 538.800 275.000 539.600 275.800 ;
        RECT 532.600 274.400 533.400 274.600 ;
        RECT 535.400 274.400 536.200 274.600 ;
        RECT 529.200 273.000 530.000 273.200 ;
        RECT 533.800 273.000 534.600 273.200 ;
        RECT 529.200 272.400 534.600 273.000 ;
        RECT 535.200 273.000 537.400 273.600 ;
        RECT 535.200 271.800 535.800 273.000 ;
        RECT 536.600 272.800 537.400 273.000 ;
        RECT 539.000 273.200 540.400 274.000 ;
        RECT 539.000 272.200 539.600 273.200 ;
        RECT 531.000 271.400 535.800 271.800 ;
        RECT 526.000 271.200 535.800 271.400 ;
        RECT 537.200 271.600 539.600 272.200 ;
        RECT 526.000 271.000 531.800 271.200 ;
        RECT 526.000 270.800 531.600 271.000 ;
        RECT 532.400 270.200 533.200 270.400 ;
        RECT 528.200 269.600 533.200 270.200 ;
        RECT 528.200 269.400 529.000 269.600 ;
        RECT 530.800 269.400 531.600 269.600 ;
        RECT 529.800 268.400 530.600 268.600 ;
        RECT 537.200 268.400 537.800 271.600 ;
        RECT 543.600 271.200 544.400 279.800 ;
        RECT 545.200 272.400 546.000 279.800 ;
        RECT 545.200 271.800 547.400 272.400 ;
        RECT 540.200 270.600 544.400 271.200 ;
        RECT 540.200 270.400 541.000 270.600 ;
        RECT 543.600 270.300 544.400 270.600 ;
        RECT 546.800 271.200 547.400 271.800 ;
        RECT 546.800 270.400 548.000 271.200 ;
        RECT 545.200 270.300 546.000 270.400 ;
        RECT 541.800 269.800 542.600 270.000 ;
        RECT 538.800 269.200 542.600 269.800 ;
        RECT 543.600 269.700 546.000 270.300 ;
        RECT 538.800 269.000 539.600 269.200 ;
        RECT 526.800 267.800 537.800 268.400 ;
        RECT 526.800 267.600 528.400 267.800 ;
        RECT 524.400 264.800 525.200 266.400 ;
        RECT 526.000 262.200 526.800 267.000 ;
        RECT 531.000 265.600 531.600 267.800 ;
        RECT 535.600 267.600 537.400 267.800 ;
        RECT 543.600 267.200 544.400 269.700 ;
        RECT 545.200 268.800 546.000 269.700 ;
        RECT 546.800 267.400 547.400 270.400 ;
        RECT 540.600 266.600 544.400 267.200 ;
        RECT 540.600 266.400 541.400 266.600 ;
        RECT 529.200 264.200 530.000 265.000 ;
        RECT 530.800 264.800 531.600 265.600 ;
        RECT 532.600 265.400 533.400 265.600 ;
        RECT 532.600 264.800 535.400 265.400 ;
        RECT 534.800 264.200 535.400 264.800 ;
        RECT 538.800 264.200 539.600 265.000 ;
        RECT 529.200 263.600 531.200 264.200 ;
        RECT 530.400 262.200 531.200 263.600 ;
        RECT 534.800 262.200 535.600 264.200 ;
        RECT 538.800 263.600 540.200 264.200 ;
        RECT 539.000 262.200 540.200 263.600 ;
        RECT 543.600 262.200 544.400 266.600 ;
        RECT 545.200 266.800 547.400 267.400 ;
        RECT 545.200 262.200 546.000 266.800 ;
        RECT 1.200 255.600 2.000 257.200 ;
        RECT 2.800 252.300 3.600 259.800 ;
        RECT 6.000 257.800 6.800 259.800 ;
        RECT 4.400 255.600 5.200 257.200 ;
        RECT 6.200 254.400 6.800 257.800 ;
        RECT 11.800 256.400 12.600 259.800 ;
        RECT 10.800 255.800 12.600 256.400 ;
        RECT 14.000 255.800 14.800 259.800 ;
        RECT 18.200 256.800 19.000 259.800 ;
        RECT 22.000 257.800 22.800 259.800 ;
        RECT 18.200 255.800 19.600 256.800 ;
        RECT 6.000 253.600 6.800 254.400 ;
        RECT 9.200 253.600 10.000 255.200 ;
        RECT 4.400 252.300 5.200 252.400 ;
        RECT 2.800 251.700 5.200 252.300 ;
        RECT 2.800 242.200 3.600 251.700 ;
        RECT 4.400 251.600 5.200 251.700 ;
        RECT 6.200 250.200 6.800 253.600 ;
        RECT 7.600 250.800 8.400 252.400 ;
        RECT 6.000 249.400 7.800 250.200 ;
        RECT 7.000 244.400 7.800 249.400 ;
        RECT 7.000 243.600 8.400 244.400 ;
        RECT 7.000 242.200 7.800 243.600 ;
        RECT 10.800 242.200 11.600 255.800 ;
        RECT 14.200 255.600 14.800 255.800 ;
        RECT 14.200 255.200 16.000 255.600 ;
        RECT 14.200 255.000 18.400 255.200 ;
        RECT 15.400 254.600 18.400 255.000 ;
        RECT 17.600 254.400 18.400 254.600 ;
        RECT 14.000 252.800 14.800 254.400 ;
        RECT 16.000 253.800 16.800 254.000 ;
        RECT 15.800 253.200 16.800 253.800 ;
        RECT 15.800 252.400 16.400 253.200 ;
        RECT 15.600 251.600 16.400 252.400 ;
        RECT 17.600 251.000 18.200 254.400 ;
        RECT 19.000 252.400 19.600 255.800 ;
        RECT 22.000 254.400 22.600 257.800 ;
        RECT 23.600 255.600 24.400 257.200 ;
        RECT 25.200 255.800 26.000 259.800 ;
        RECT 29.400 258.400 30.200 259.800 ;
        RECT 29.400 257.600 30.800 258.400 ;
        RECT 29.400 256.800 30.200 257.600 ;
        RECT 29.400 255.800 30.800 256.800 ;
        RECT 31.600 256.000 32.400 259.800 ;
        RECT 34.800 256.000 35.600 259.800 ;
        RECT 31.600 255.800 35.600 256.000 ;
        RECT 36.400 255.800 37.200 259.800 ;
        RECT 39.600 257.800 40.400 259.800 ;
        RECT 25.400 255.600 26.000 255.800 ;
        RECT 25.400 255.200 27.200 255.600 ;
        RECT 25.400 255.000 29.600 255.200 ;
        RECT 26.600 254.600 29.600 255.000 ;
        RECT 28.800 254.400 29.600 254.600 ;
        RECT 22.000 253.600 22.800 254.400 ;
        RECT 18.800 251.600 19.600 252.400 ;
        RECT 15.800 250.400 18.200 251.000 ;
        RECT 12.400 248.800 13.200 250.400 ;
        RECT 15.800 246.200 16.400 250.400 ;
        RECT 19.000 250.200 19.600 251.600 ;
        RECT 20.400 250.800 21.200 252.400 ;
        RECT 22.000 252.300 22.600 253.600 ;
        RECT 25.200 252.800 26.000 254.400 ;
        RECT 27.200 253.800 28.000 254.000 ;
        RECT 27.000 253.200 28.000 253.800 ;
        RECT 27.000 252.400 27.600 253.200 ;
        RECT 23.600 252.300 24.400 252.400 ;
        RECT 22.000 251.700 24.400 252.300 ;
        RECT 22.000 250.200 22.600 251.700 ;
        RECT 23.600 251.600 24.400 251.700 ;
        RECT 26.800 251.600 27.600 252.400 ;
        RECT 28.800 251.000 29.400 254.400 ;
        RECT 30.200 252.400 30.800 255.800 ;
        RECT 31.800 255.400 35.400 255.800 ;
        RECT 32.400 254.400 33.200 254.800 ;
        RECT 36.400 254.400 37.000 255.800 ;
        RECT 39.600 254.400 40.200 257.800 ;
        RECT 41.200 255.600 42.000 257.200 ;
        RECT 45.400 256.400 46.200 259.800 ;
        RECT 44.400 255.800 46.200 256.400 ;
        RECT 31.600 253.800 33.200 254.400 ;
        RECT 31.600 253.600 32.400 253.800 ;
        RECT 34.600 253.600 37.200 254.400 ;
        RECT 39.600 253.600 40.400 254.400 ;
        RECT 42.800 253.600 43.600 255.200 ;
        RECT 30.000 251.600 30.800 252.400 ;
        RECT 31.600 252.300 32.400 252.400 ;
        RECT 33.200 252.300 34.000 253.200 ;
        RECT 31.600 251.700 34.000 252.300 ;
        RECT 31.600 251.600 32.400 251.700 ;
        RECT 33.200 251.600 34.000 251.700 ;
        RECT 34.600 252.400 35.200 253.600 ;
        RECT 34.600 251.600 35.600 252.400 ;
        RECT 27.000 250.400 29.400 251.000 ;
        RECT 15.600 242.200 16.400 246.200 ;
        RECT 18.800 242.200 19.600 250.200 ;
        RECT 21.000 249.400 22.800 250.200 ;
        RECT 21.000 242.200 21.800 249.400 ;
        RECT 27.000 246.200 27.600 250.400 ;
        RECT 30.200 250.200 30.800 251.600 ;
        RECT 34.600 250.200 35.200 251.600 ;
        RECT 38.000 250.800 38.800 252.400 ;
        RECT 36.400 250.200 37.200 250.400 ;
        RECT 39.600 250.200 40.200 253.600 ;
        RECT 26.800 242.200 27.600 246.200 ;
        RECT 30.000 242.200 30.800 250.200 ;
        RECT 34.200 249.600 35.200 250.200 ;
        RECT 35.800 249.600 37.200 250.200 ;
        RECT 34.200 242.200 35.000 249.600 ;
        RECT 35.800 248.400 36.400 249.600 ;
        RECT 35.600 247.600 36.400 248.400 ;
        RECT 38.600 249.400 40.400 250.200 ;
        RECT 38.600 244.400 39.400 249.400 ;
        RECT 38.600 243.600 40.400 244.400 ;
        RECT 38.600 242.200 39.400 243.600 ;
        RECT 44.400 242.200 45.200 255.800 ;
        RECT 51.200 254.200 52.000 259.800 ;
        RECT 56.600 258.400 57.400 259.800 ;
        RECT 56.600 257.600 58.000 258.400 ;
        RECT 56.600 256.400 57.400 257.600 ;
        RECT 55.600 255.800 57.400 256.400 ;
        RECT 59.400 256.400 60.200 259.800 ;
        RECT 65.200 257.800 66.000 259.800 ;
        RECT 59.400 255.800 61.200 256.400 ;
        RECT 51.200 253.800 53.000 254.200 ;
        RECT 51.400 253.600 53.000 253.800 ;
        RECT 54.000 253.600 54.800 255.200 ;
        RECT 49.200 251.600 50.800 252.400 ;
        RECT 46.000 248.800 46.800 250.400 ;
        RECT 47.600 249.600 48.400 251.200 ;
        RECT 52.400 250.400 53.000 253.600 ;
        RECT 52.400 249.600 53.200 250.400 ;
        RECT 50.800 247.600 51.600 249.200 ;
        RECT 52.400 247.000 53.000 249.600 ;
        RECT 49.400 246.400 53.000 247.000 ;
        RECT 49.400 246.200 50.000 246.400 ;
        RECT 49.200 242.200 50.000 246.200 ;
        RECT 52.400 246.200 53.000 246.400 ;
        RECT 52.400 242.200 53.200 246.200 ;
        RECT 55.600 242.200 56.400 255.800 ;
        RECT 60.400 252.300 61.200 255.800 ;
        RECT 63.600 255.600 64.400 257.200 ;
        RECT 62.000 254.300 62.800 255.200 ;
        RECT 63.700 254.300 64.300 255.600 ;
        RECT 65.400 254.400 66.000 257.800 ;
        RECT 68.400 255.800 69.200 259.800 ;
        RECT 70.000 256.000 70.800 259.800 ;
        RECT 73.200 256.000 74.000 259.800 ;
        RECT 76.400 257.800 77.200 259.800 ;
        RECT 70.000 255.800 74.000 256.000 ;
        RECT 68.600 254.400 69.200 255.800 ;
        RECT 70.200 255.400 73.800 255.800 ;
        RECT 74.800 255.600 75.600 257.200 ;
        RECT 72.400 254.400 73.200 254.800 ;
        RECT 76.600 254.400 77.200 257.800 ;
        RECT 81.200 256.000 82.000 259.800 ;
        RECT 62.000 253.700 64.300 254.300 ;
        RECT 62.000 253.600 62.800 253.700 ;
        RECT 65.200 253.600 66.000 254.400 ;
        RECT 68.400 253.600 71.000 254.400 ;
        RECT 72.400 253.800 74.000 254.400 ;
        RECT 73.200 253.600 74.000 253.800 ;
        RECT 76.400 253.600 77.200 254.400 ;
        RECT 63.600 252.300 64.400 252.400 ;
        RECT 60.400 251.700 64.400 252.300 ;
        RECT 57.200 248.800 58.000 250.400 ;
        RECT 58.800 248.800 59.600 250.400 ;
        RECT 60.400 242.200 61.200 251.700 ;
        RECT 63.600 251.600 64.400 251.700 ;
        RECT 65.400 250.200 66.000 253.600 ;
        RECT 70.400 252.400 71.000 253.600 ;
        RECT 66.800 252.300 67.600 252.400 ;
        RECT 68.400 252.300 69.200 252.400 ;
        RECT 66.800 251.700 69.200 252.300 ;
        RECT 66.800 250.800 67.600 251.700 ;
        RECT 68.400 251.600 69.200 251.700 ;
        RECT 70.000 251.600 71.000 252.400 ;
        RECT 71.600 251.600 72.400 253.200 ;
        RECT 68.400 250.200 69.200 250.400 ;
        RECT 70.400 250.200 71.000 251.600 ;
        RECT 76.600 250.200 77.200 253.600 ;
        RECT 81.000 255.200 82.000 256.000 ;
        RECT 78.000 252.300 78.800 252.400 ;
        RECT 79.600 252.300 80.400 252.400 ;
        RECT 78.000 251.700 80.400 252.300 ;
        RECT 78.000 250.800 78.800 251.700 ;
        RECT 79.600 251.600 80.400 251.700 ;
        RECT 81.000 250.800 81.800 255.200 ;
        RECT 82.800 254.600 83.600 259.800 ;
        RECT 89.200 256.600 90.000 259.800 ;
        RECT 90.800 257.000 91.600 259.800 ;
        RECT 92.400 257.000 93.200 259.800 ;
        RECT 94.000 257.000 94.800 259.800 ;
        RECT 95.600 257.000 96.400 259.800 ;
        RECT 98.800 257.000 99.600 259.800 ;
        RECT 102.000 257.000 102.800 259.800 ;
        RECT 103.600 257.000 104.400 259.800 ;
        RECT 105.200 257.000 106.000 259.800 ;
        RECT 87.600 255.800 90.000 256.600 ;
        RECT 106.800 256.600 107.600 259.800 ;
        RECT 87.600 255.200 88.400 255.800 ;
        RECT 82.400 254.000 83.600 254.600 ;
        RECT 86.600 254.600 88.400 255.200 ;
        RECT 92.400 255.600 93.400 256.400 ;
        RECT 96.400 255.600 98.000 256.400 ;
        RECT 98.800 255.800 103.400 256.400 ;
        RECT 106.800 255.800 109.400 256.600 ;
        RECT 98.800 255.600 99.600 255.800 ;
        RECT 82.400 252.000 83.000 254.000 ;
        RECT 86.600 253.400 87.400 254.600 ;
        RECT 83.600 252.600 87.400 253.400 ;
        RECT 92.400 252.800 93.200 255.600 ;
        RECT 98.800 254.800 99.600 255.000 ;
        RECT 95.200 254.200 99.600 254.800 ;
        RECT 95.200 254.000 96.000 254.200 ;
        RECT 100.400 253.600 101.200 255.200 ;
        RECT 102.600 253.400 103.400 255.800 ;
        RECT 108.600 255.200 109.400 255.800 ;
        RECT 108.600 254.400 111.600 255.200 ;
        RECT 113.200 253.800 114.000 259.800 ;
        RECT 119.600 257.800 120.400 259.800 ;
        RECT 122.800 258.400 123.600 259.800 ;
        RECT 95.600 252.600 98.800 253.400 ;
        RECT 102.600 252.600 104.600 253.400 ;
        RECT 105.200 253.000 114.000 253.800 ;
        RECT 89.200 252.000 90.000 252.600 ;
        RECT 106.800 252.000 107.600 252.400 ;
        RECT 110.000 252.000 110.800 252.400 ;
        RECT 111.800 252.000 112.600 252.200 ;
        RECT 82.400 251.400 83.200 252.000 ;
        RECT 89.200 251.400 112.600 252.000 ;
        RECT 65.200 249.400 67.000 250.200 ;
        RECT 68.400 249.600 69.800 250.200 ;
        RECT 70.400 249.600 71.400 250.200 ;
        RECT 66.200 244.400 67.000 249.400 ;
        RECT 69.200 248.400 69.800 249.600 ;
        RECT 69.200 247.600 70.000 248.400 ;
        RECT 65.200 243.600 67.000 244.400 ;
        RECT 66.200 242.200 67.000 243.600 ;
        RECT 70.600 242.200 71.400 249.600 ;
        RECT 76.400 249.400 78.200 250.200 ;
        RECT 81.000 250.000 82.000 250.800 ;
        RECT 77.400 246.400 78.200 249.400 ;
        RECT 76.400 245.600 78.200 246.400 ;
        RECT 77.400 242.200 78.200 245.600 ;
        RECT 81.200 242.200 82.000 250.000 ;
        RECT 82.600 249.600 83.200 251.400 ;
        RECT 82.600 249.000 91.600 249.600 ;
        RECT 82.600 247.400 83.200 249.000 ;
        RECT 90.800 248.800 91.600 249.000 ;
        RECT 94.000 249.000 102.600 249.600 ;
        RECT 94.000 248.800 94.800 249.000 ;
        RECT 85.800 247.600 88.400 248.400 ;
        RECT 82.600 246.800 85.200 247.400 ;
        RECT 84.400 242.200 85.200 246.800 ;
        RECT 87.600 242.200 88.400 247.600 ;
        RECT 89.000 246.800 93.200 247.600 ;
        RECT 90.800 242.200 91.600 245.000 ;
        RECT 92.400 242.200 93.200 245.000 ;
        RECT 94.000 242.200 94.800 245.000 ;
        RECT 95.600 242.200 96.400 248.400 ;
        RECT 98.800 247.600 101.400 248.400 ;
        RECT 102.000 248.200 102.600 249.000 ;
        RECT 103.600 249.400 104.400 249.600 ;
        RECT 103.600 249.000 109.000 249.400 ;
        RECT 103.600 248.800 109.800 249.000 ;
        RECT 108.400 248.200 109.800 248.800 ;
        RECT 102.000 247.600 107.800 248.200 ;
        RECT 110.800 248.000 112.400 248.800 ;
        RECT 110.800 247.600 111.400 248.000 ;
        RECT 98.800 242.200 99.600 247.000 ;
        RECT 102.000 242.200 102.800 247.000 ;
        RECT 107.200 246.800 111.400 247.600 ;
        RECT 113.200 247.400 114.000 253.000 ;
        RECT 119.200 257.600 120.400 257.800 ;
        RECT 122.600 257.600 123.600 258.400 ;
        RECT 119.200 257.000 123.200 257.600 ;
        RECT 119.200 250.400 119.800 257.000 ;
        RECT 123.400 256.300 125.200 256.400 ;
        RECT 132.400 256.300 133.200 256.400 ;
        RECT 123.400 255.700 133.200 256.300 ;
        RECT 136.600 255.800 138.200 259.800 ;
        RECT 123.400 255.600 125.200 255.700 ;
        RECT 132.400 255.600 133.200 255.700 ;
        RECT 122.000 253.600 123.600 254.400 ;
        RECT 135.600 253.600 136.400 254.400 ;
        RECT 135.800 253.200 136.400 253.600 ;
        RECT 135.800 252.400 136.600 253.200 ;
        RECT 137.200 252.400 137.800 255.800 ;
        RECT 138.800 252.800 139.600 254.400 ;
        RECT 120.400 251.600 122.000 252.400 ;
        RECT 132.400 252.300 133.200 252.400 ;
        RECT 134.000 252.300 134.800 252.400 ;
        RECT 132.400 251.700 134.800 252.300 ;
        RECT 132.400 251.600 133.200 251.700 ;
        RECT 134.000 250.800 134.800 251.700 ;
        RECT 137.200 251.600 138.000 252.400 ;
        RECT 140.400 252.200 141.200 252.400 ;
        RECT 139.600 251.600 141.200 252.200 ;
        RECT 137.200 251.400 137.800 251.600 ;
        RECT 135.800 250.800 137.800 251.400 ;
        RECT 139.600 251.200 140.400 251.600 ;
        RECT 116.400 249.800 119.800 250.400 ;
        RECT 135.800 250.200 136.400 250.800 ;
        RECT 116.400 249.600 117.200 249.800 ;
        RECT 116.600 249.000 117.200 249.600 ;
        RECT 118.200 249.000 121.800 249.200 ;
        RECT 112.000 246.800 114.000 247.400 ;
        RECT 103.600 242.200 104.400 245.000 ;
        RECT 105.200 242.200 106.000 245.000 ;
        RECT 108.400 242.200 109.200 246.800 ;
        RECT 112.000 246.200 112.600 246.800 ;
        RECT 111.600 245.600 112.600 246.200 ;
        RECT 111.600 242.200 112.400 245.600 ;
        RECT 114.800 243.000 115.600 249.000 ;
        RECT 116.400 243.400 117.200 249.000 ;
        RECT 118.000 248.600 121.800 249.000 ;
        RECT 115.000 242.800 115.600 243.000 ;
        RECT 118.000 243.000 118.800 248.600 ;
        RECT 121.200 248.200 121.800 248.600 ;
        RECT 123.000 248.800 126.600 249.400 ;
        RECT 123.000 248.200 123.600 248.800 ;
        RECT 118.000 242.800 118.600 243.000 ;
        RECT 115.000 242.200 118.600 242.800 ;
        RECT 119.600 242.800 120.400 248.000 ;
        RECT 121.200 243.400 122.000 248.200 ;
        RECT 122.800 242.800 123.600 248.200 ;
        RECT 119.600 242.200 123.600 242.800 ;
        RECT 126.000 248.200 126.600 248.800 ;
        RECT 126.000 242.200 126.800 248.200 ;
        RECT 134.000 242.800 134.800 250.200 ;
        RECT 135.600 243.400 136.400 250.200 ;
        RECT 137.200 249.600 141.200 250.200 ;
        RECT 137.200 242.800 138.000 249.600 ;
        RECT 134.000 242.200 138.000 242.800 ;
        RECT 140.400 242.200 141.200 249.600 ;
        RECT 142.000 242.200 142.800 259.800 ;
        RECT 143.600 255.600 144.400 257.200 ;
        RECT 145.200 253.800 146.000 259.800 ;
        RECT 151.600 256.600 152.400 259.800 ;
        RECT 153.200 257.000 154.000 259.800 ;
        RECT 154.800 257.000 155.600 259.800 ;
        RECT 156.400 257.000 157.200 259.800 ;
        RECT 159.600 257.000 160.400 259.800 ;
        RECT 162.800 257.000 163.600 259.800 ;
        RECT 164.400 257.000 165.200 259.800 ;
        RECT 166.000 257.000 166.800 259.800 ;
        RECT 167.600 257.000 168.400 259.800 ;
        RECT 149.800 255.800 152.400 256.600 ;
        RECT 169.200 256.600 170.000 259.800 ;
        RECT 155.800 255.800 160.400 256.400 ;
        RECT 149.800 255.200 150.600 255.800 ;
        RECT 147.600 254.400 150.600 255.200 ;
        RECT 145.200 253.000 154.000 253.800 ;
        RECT 155.800 253.400 156.600 255.800 ;
        RECT 159.600 255.600 160.400 255.800 ;
        RECT 161.200 255.600 162.800 256.400 ;
        RECT 165.800 255.600 166.800 256.400 ;
        RECT 169.200 255.800 171.600 256.600 ;
        RECT 158.000 253.600 158.800 255.200 ;
        RECT 159.600 254.800 160.400 255.000 ;
        RECT 159.600 254.200 164.000 254.800 ;
        RECT 163.200 254.000 164.000 254.200 ;
        RECT 145.200 247.400 146.000 253.000 ;
        RECT 154.600 252.600 156.600 253.400 ;
        RECT 160.400 252.600 163.600 253.400 ;
        RECT 166.000 252.800 166.800 255.600 ;
        RECT 170.800 255.200 171.600 255.800 ;
        RECT 170.800 254.600 172.600 255.200 ;
        RECT 171.800 253.400 172.600 254.600 ;
        RECT 175.600 254.600 176.400 259.800 ;
        RECT 177.200 256.000 178.000 259.800 ;
        RECT 177.200 255.200 178.200 256.000 ;
        RECT 175.600 254.000 176.800 254.600 ;
        RECT 171.800 252.600 175.600 253.400 ;
        RECT 146.600 252.000 147.400 252.200 ;
        RECT 151.600 252.000 152.400 252.400 ;
        RECT 158.000 252.000 158.800 252.400 ;
        RECT 169.200 252.000 170.000 252.600 ;
        RECT 176.200 252.000 176.800 254.000 ;
        RECT 146.600 251.400 170.000 252.000 ;
        RECT 176.000 251.400 176.800 252.000 ;
        RECT 176.000 249.600 176.600 251.400 ;
        RECT 177.400 250.800 178.200 255.200 ;
        RECT 154.800 249.400 155.600 249.600 ;
        RECT 150.200 249.000 155.600 249.400 ;
        RECT 149.400 248.800 155.600 249.000 ;
        RECT 156.600 249.000 165.200 249.600 ;
        RECT 146.800 248.000 148.400 248.800 ;
        RECT 149.400 248.200 150.800 248.800 ;
        RECT 156.600 248.200 157.200 249.000 ;
        RECT 164.400 248.800 165.200 249.000 ;
        RECT 167.600 249.000 176.600 249.600 ;
        RECT 167.600 248.800 168.400 249.000 ;
        RECT 147.800 247.600 148.400 248.000 ;
        RECT 151.400 247.600 157.200 248.200 ;
        RECT 157.800 247.600 160.400 248.400 ;
        RECT 145.200 246.800 147.200 247.400 ;
        RECT 147.800 246.800 152.000 247.600 ;
        RECT 146.600 246.200 147.200 246.800 ;
        RECT 146.600 245.600 147.600 246.200 ;
        RECT 146.800 242.200 147.600 245.600 ;
        RECT 150.000 242.200 150.800 246.800 ;
        RECT 153.200 242.200 154.000 245.000 ;
        RECT 154.800 242.200 155.600 245.000 ;
        RECT 156.400 242.200 157.200 247.000 ;
        RECT 159.600 242.200 160.400 247.000 ;
        RECT 162.800 242.200 163.600 248.400 ;
        RECT 170.800 247.600 173.400 248.400 ;
        RECT 166.000 246.800 170.200 247.600 ;
        RECT 164.400 242.200 165.200 245.000 ;
        RECT 166.000 242.200 166.800 245.000 ;
        RECT 167.600 242.200 168.400 245.000 ;
        RECT 170.800 242.200 171.600 247.600 ;
        RECT 176.000 247.400 176.600 249.000 ;
        RECT 174.000 246.800 176.600 247.400 ;
        RECT 177.200 250.000 178.200 250.800 ;
        RECT 174.000 242.200 174.800 246.800 ;
        RECT 177.200 242.200 178.000 250.000 ;
        RECT 182.000 242.200 182.800 259.800 ;
        RECT 187.800 258.400 188.600 259.800 ;
        RECT 187.800 257.600 189.200 258.400 ;
        RECT 187.800 256.400 188.600 257.600 ;
        RECT 186.800 255.800 188.600 256.400 ;
        RECT 183.600 253.600 184.400 255.200 ;
        RECT 185.200 253.600 186.000 255.200 ;
        RECT 183.700 252.300 184.300 253.600 ;
        RECT 186.800 252.300 187.600 255.800 ;
        RECT 183.700 251.700 187.600 252.300 ;
        RECT 186.800 242.200 187.600 251.700 ;
        RECT 188.400 248.800 189.200 250.400 ;
        RECT 190.000 242.200 190.800 259.800 ;
        RECT 191.600 256.300 192.400 257.200 ;
        RECT 193.200 256.300 194.000 259.800 ;
        RECT 191.600 255.700 194.000 256.300 ;
        RECT 194.800 256.000 195.600 259.800 ;
        RECT 198.000 256.000 198.800 259.800 ;
        RECT 201.200 257.800 202.000 259.800 ;
        RECT 194.800 255.800 198.800 256.000 ;
        RECT 191.600 255.600 192.400 255.700 ;
        RECT 193.400 254.400 194.000 255.700 ;
        RECT 195.000 255.400 198.600 255.800 ;
        RECT 199.600 255.600 200.400 257.200 ;
        RECT 201.400 255.600 202.000 257.800 ;
        RECT 204.400 256.300 205.200 259.800 ;
        RECT 206.000 256.300 206.800 256.400 ;
        RECT 204.400 255.800 206.800 256.300 ;
        RECT 207.600 256.000 208.400 259.800 ;
        RECT 204.500 255.700 206.800 255.800 ;
        RECT 201.400 255.000 203.800 255.600 ;
        RECT 197.200 254.400 198.000 254.800 ;
        RECT 193.200 253.600 195.800 254.400 ;
        RECT 197.200 254.300 198.800 254.400 ;
        RECT 201.200 254.300 202.200 254.400 ;
        RECT 197.200 253.800 202.200 254.300 ;
        RECT 198.000 253.700 202.200 253.800 ;
        RECT 198.000 253.600 198.800 253.700 ;
        RECT 201.200 253.600 202.200 253.700 ;
        RECT 193.200 250.200 194.000 250.400 ;
        RECT 195.200 250.200 195.800 253.600 ;
        RECT 196.400 252.300 197.200 253.200 ;
        RECT 201.600 252.800 202.400 253.600 ;
        RECT 198.000 252.300 198.800 252.400 ;
        RECT 196.400 251.700 198.800 252.300 ;
        RECT 203.200 252.000 203.800 255.000 ;
        RECT 204.600 252.400 205.200 255.700 ;
        RECT 206.000 255.600 206.800 255.700 ;
        RECT 196.400 251.600 197.200 251.700 ;
        RECT 198.000 251.600 198.800 251.700 ;
        RECT 203.000 251.400 203.800 252.000 ;
        RECT 204.400 251.600 205.200 252.400 ;
        RECT 199.600 251.200 203.800 251.400 ;
        RECT 199.600 250.800 203.600 251.200 ;
        RECT 193.200 249.600 194.600 250.200 ;
        RECT 195.200 249.600 196.200 250.200 ;
        RECT 194.000 248.400 194.600 249.600 ;
        RECT 194.000 247.600 194.800 248.400 ;
        RECT 195.400 242.200 196.200 249.600 ;
        RECT 199.600 242.200 200.400 250.800 ;
        RECT 204.600 250.200 205.200 251.600 ;
        RECT 203.800 249.600 205.200 250.200 ;
        RECT 207.400 255.200 208.400 256.000 ;
        RECT 207.400 250.800 208.200 255.200 ;
        RECT 209.200 254.600 210.000 259.800 ;
        RECT 215.600 256.600 216.400 259.800 ;
        RECT 217.200 257.000 218.000 259.800 ;
        RECT 218.800 257.000 219.600 259.800 ;
        RECT 220.400 257.000 221.200 259.800 ;
        RECT 222.000 257.000 222.800 259.800 ;
        RECT 225.200 257.000 226.000 259.800 ;
        RECT 228.400 257.000 229.200 259.800 ;
        RECT 230.000 257.000 230.800 259.800 ;
        RECT 231.600 257.000 232.400 259.800 ;
        RECT 214.000 255.800 216.400 256.600 ;
        RECT 233.200 256.600 234.000 259.800 ;
        RECT 214.000 255.200 214.800 255.800 ;
        RECT 208.800 254.000 210.000 254.600 ;
        RECT 213.000 254.600 214.800 255.200 ;
        RECT 218.800 255.600 219.800 256.400 ;
        RECT 222.800 255.600 224.400 256.400 ;
        RECT 225.200 255.800 229.800 256.400 ;
        RECT 233.200 255.800 235.800 256.600 ;
        RECT 225.200 255.600 226.000 255.800 ;
        RECT 208.800 252.000 209.400 254.000 ;
        RECT 213.000 253.400 213.800 254.600 ;
        RECT 210.000 252.600 213.800 253.400 ;
        RECT 218.800 252.800 219.600 255.600 ;
        RECT 225.200 254.800 226.000 255.000 ;
        RECT 221.600 254.200 226.000 254.800 ;
        RECT 221.600 254.000 222.400 254.200 ;
        RECT 226.800 253.600 227.600 255.200 ;
        RECT 229.000 253.400 229.800 255.800 ;
        RECT 235.000 255.200 235.800 255.800 ;
        RECT 235.000 254.400 238.000 255.200 ;
        RECT 239.600 253.800 240.400 259.800 ;
        RECT 241.800 258.400 242.600 259.800 ;
        RECT 241.800 257.600 243.600 258.400 ;
        RECT 241.800 256.400 242.600 257.600 ;
        RECT 241.800 255.800 243.600 256.400 ;
        RECT 247.600 256.000 248.400 259.800 ;
        RECT 222.000 252.600 225.200 253.400 ;
        RECT 229.000 252.600 231.000 253.400 ;
        RECT 231.600 253.000 240.400 253.800 ;
        RECT 215.600 252.000 216.400 252.600 ;
        RECT 233.200 252.000 234.000 252.400 ;
        RECT 238.200 252.000 239.000 252.200 ;
        RECT 208.800 251.400 209.600 252.000 ;
        RECT 215.600 251.400 239.000 252.000 ;
        RECT 207.400 250.000 208.400 250.800 ;
        RECT 203.800 242.200 204.600 249.600 ;
        RECT 207.600 242.200 208.400 250.000 ;
        RECT 209.000 249.600 209.600 251.400 ;
        RECT 209.000 249.000 218.000 249.600 ;
        RECT 209.000 247.400 209.600 249.000 ;
        RECT 217.200 248.800 218.000 249.000 ;
        RECT 220.400 249.000 229.000 249.600 ;
        RECT 220.400 248.800 221.200 249.000 ;
        RECT 212.200 247.600 214.800 248.400 ;
        RECT 209.000 246.800 211.600 247.400 ;
        RECT 210.800 242.200 211.600 246.800 ;
        RECT 214.000 242.200 214.800 247.600 ;
        RECT 215.400 246.800 219.600 247.600 ;
        RECT 217.200 242.200 218.000 245.000 ;
        RECT 218.800 242.200 219.600 245.000 ;
        RECT 220.400 242.200 221.200 245.000 ;
        RECT 222.000 242.200 222.800 248.400 ;
        RECT 225.200 247.600 227.800 248.400 ;
        RECT 228.400 248.200 229.000 249.000 ;
        RECT 230.000 249.400 230.800 249.600 ;
        RECT 230.000 249.000 235.400 249.400 ;
        RECT 230.000 248.800 236.200 249.000 ;
        RECT 234.800 248.200 236.200 248.800 ;
        RECT 228.400 247.600 234.200 248.200 ;
        RECT 237.200 248.000 238.800 248.800 ;
        RECT 237.200 247.600 237.800 248.000 ;
        RECT 225.200 242.200 226.000 247.000 ;
        RECT 228.400 242.200 229.200 247.000 ;
        RECT 233.600 246.800 237.800 247.600 ;
        RECT 239.600 247.400 240.400 253.000 ;
        RECT 241.200 248.800 242.000 250.400 ;
        RECT 238.400 246.800 240.400 247.400 ;
        RECT 230.000 242.200 230.800 245.000 ;
        RECT 231.600 242.200 232.400 245.000 ;
        RECT 234.800 242.200 235.600 246.800 ;
        RECT 238.400 246.200 239.000 246.800 ;
        RECT 238.000 245.600 239.000 246.200 ;
        RECT 238.000 242.200 238.800 245.600 ;
        RECT 242.800 242.200 243.600 255.800 ;
        RECT 247.400 255.200 248.400 256.000 ;
        RECT 244.400 254.300 245.200 255.200 ;
        RECT 247.400 254.300 248.200 255.200 ;
        RECT 249.200 254.600 250.000 259.800 ;
        RECT 255.600 256.600 256.400 259.800 ;
        RECT 257.200 257.000 258.000 259.800 ;
        RECT 258.800 257.000 259.600 259.800 ;
        RECT 260.400 257.000 261.200 259.800 ;
        RECT 262.000 257.000 262.800 259.800 ;
        RECT 265.200 257.000 266.000 259.800 ;
        RECT 268.400 257.000 269.200 259.800 ;
        RECT 270.000 257.000 270.800 259.800 ;
        RECT 271.600 257.000 272.400 259.800 ;
        RECT 254.000 255.800 256.400 256.600 ;
        RECT 273.200 256.600 274.000 259.800 ;
        RECT 254.000 255.200 254.800 255.800 ;
        RECT 244.400 253.700 248.200 254.300 ;
        RECT 244.400 253.600 245.200 253.700 ;
        RECT 247.400 250.800 248.200 253.700 ;
        RECT 248.800 254.000 250.000 254.600 ;
        RECT 253.000 254.600 254.800 255.200 ;
        RECT 258.800 255.600 259.800 256.400 ;
        RECT 262.800 255.600 264.400 256.400 ;
        RECT 265.200 255.800 269.800 256.400 ;
        RECT 273.200 255.800 275.800 256.600 ;
        RECT 265.200 255.600 266.000 255.800 ;
        RECT 248.800 252.000 249.400 254.000 ;
        RECT 253.000 253.400 253.800 254.600 ;
        RECT 250.000 252.600 253.800 253.400 ;
        RECT 258.800 252.800 259.600 255.600 ;
        RECT 265.200 254.800 266.000 255.000 ;
        RECT 261.600 254.200 266.000 254.800 ;
        RECT 261.600 254.000 262.400 254.200 ;
        RECT 266.800 253.600 267.600 255.200 ;
        RECT 269.000 253.400 269.800 255.800 ;
        RECT 275.000 255.200 275.800 255.800 ;
        RECT 275.000 254.400 278.000 255.200 ;
        RECT 279.600 253.800 280.400 259.800 ;
        RECT 289.200 256.000 290.000 259.800 ;
        RECT 262.000 252.600 265.200 253.400 ;
        RECT 269.000 252.600 271.000 253.400 ;
        RECT 271.600 253.000 280.400 253.800 ;
        RECT 248.800 251.400 249.600 252.000 ;
        RECT 247.400 250.000 248.400 250.800 ;
        RECT 247.600 242.200 248.400 250.000 ;
        RECT 249.000 249.600 249.600 251.400 ;
        RECT 250.200 250.800 251.000 251.000 ;
        RECT 250.200 250.200 277.200 250.800 ;
        RECT 273.000 250.000 273.800 250.200 ;
        RECT 276.400 249.600 277.200 250.200 ;
        RECT 249.000 249.000 258.000 249.600 ;
        RECT 249.000 247.400 249.600 249.000 ;
        RECT 257.200 248.800 258.000 249.000 ;
        RECT 260.400 249.000 269.000 249.600 ;
        RECT 260.400 248.800 261.200 249.000 ;
        RECT 252.200 247.600 254.800 248.400 ;
        RECT 249.000 246.800 251.600 247.400 ;
        RECT 250.800 242.200 251.600 246.800 ;
        RECT 254.000 242.200 254.800 247.600 ;
        RECT 255.400 246.800 259.600 247.600 ;
        RECT 257.200 242.200 258.000 245.000 ;
        RECT 258.800 242.200 259.600 245.000 ;
        RECT 260.400 242.200 261.200 245.000 ;
        RECT 262.000 242.200 262.800 248.400 ;
        RECT 265.200 247.600 267.800 248.400 ;
        RECT 268.400 248.200 269.000 249.000 ;
        RECT 270.000 249.400 270.800 249.600 ;
        RECT 270.000 249.000 275.400 249.400 ;
        RECT 270.000 248.800 276.200 249.000 ;
        RECT 274.800 248.200 276.200 248.800 ;
        RECT 268.400 247.600 274.200 248.200 ;
        RECT 277.200 248.000 278.800 248.800 ;
        RECT 277.200 247.600 277.800 248.000 ;
        RECT 265.200 242.200 266.000 247.000 ;
        RECT 268.400 242.200 269.200 247.000 ;
        RECT 273.600 246.800 277.800 247.600 ;
        RECT 279.600 247.400 280.400 253.000 ;
        RECT 289.000 255.200 290.000 256.000 ;
        RECT 289.000 250.800 289.800 255.200 ;
        RECT 290.800 254.600 291.600 259.800 ;
        RECT 297.200 256.600 298.000 259.800 ;
        RECT 298.800 257.000 299.600 259.800 ;
        RECT 300.400 257.000 301.200 259.800 ;
        RECT 302.000 257.000 302.800 259.800 ;
        RECT 303.600 257.000 304.400 259.800 ;
        RECT 306.800 257.000 307.600 259.800 ;
        RECT 310.000 257.000 310.800 259.800 ;
        RECT 311.600 257.000 312.400 259.800 ;
        RECT 313.200 257.000 314.000 259.800 ;
        RECT 295.600 255.800 298.000 256.600 ;
        RECT 314.800 256.600 315.600 259.800 ;
        RECT 295.600 255.200 296.400 255.800 ;
        RECT 290.400 254.000 291.600 254.600 ;
        RECT 294.600 254.600 296.400 255.200 ;
        RECT 300.400 255.600 301.400 256.400 ;
        RECT 304.400 255.600 306.000 256.400 ;
        RECT 306.800 255.800 311.400 256.400 ;
        RECT 314.800 255.800 317.400 256.600 ;
        RECT 306.800 255.600 307.600 255.800 ;
        RECT 290.400 252.000 291.000 254.000 ;
        RECT 294.600 253.400 295.400 254.600 ;
        RECT 291.600 252.600 295.400 253.400 ;
        RECT 300.400 252.800 301.200 255.600 ;
        RECT 306.800 254.800 307.600 255.000 ;
        RECT 303.200 254.200 307.600 254.800 ;
        RECT 303.200 254.000 304.000 254.200 ;
        RECT 308.400 253.600 309.200 255.200 ;
        RECT 310.600 253.400 311.400 255.800 ;
        RECT 316.600 255.200 317.400 255.800 ;
        RECT 316.600 254.400 319.600 255.200 ;
        RECT 321.200 253.800 322.000 259.800 ;
        RECT 322.800 255.800 323.600 259.800 ;
        RECT 324.400 256.000 325.200 259.800 ;
        RECT 327.600 256.000 328.400 259.800 ;
        RECT 324.400 255.800 328.400 256.000 ;
        RECT 329.200 255.800 330.000 259.800 ;
        RECT 330.800 256.000 331.600 259.800 ;
        RECT 334.000 256.000 334.800 259.800 ;
        RECT 330.800 255.800 334.800 256.000 ;
        RECT 323.000 254.400 323.600 255.800 ;
        RECT 324.600 255.400 328.200 255.800 ;
        RECT 326.800 254.400 327.600 254.800 ;
        RECT 329.400 254.400 330.000 255.800 ;
        RECT 331.000 255.400 334.600 255.800 ;
        RECT 333.200 254.400 334.000 254.800 ;
        RECT 303.600 252.600 306.800 253.400 ;
        RECT 310.600 252.600 312.600 253.400 ;
        RECT 313.200 253.000 322.000 253.800 ;
        RECT 322.800 253.600 325.400 254.400 ;
        RECT 326.800 253.800 328.400 254.400 ;
        RECT 327.600 253.600 328.400 253.800 ;
        RECT 329.200 253.600 331.800 254.400 ;
        RECT 333.200 253.800 334.800 254.400 ;
        RECT 334.000 253.600 334.800 253.800 ;
        RECT 290.400 251.400 291.200 252.000 ;
        RECT 289.000 250.000 290.000 250.800 ;
        RECT 278.400 246.800 280.400 247.400 ;
        RECT 270.000 242.200 270.800 245.000 ;
        RECT 271.600 242.200 272.400 245.000 ;
        RECT 274.800 242.200 275.600 246.800 ;
        RECT 278.400 246.200 279.000 246.800 ;
        RECT 278.000 245.600 279.000 246.200 ;
        RECT 278.000 242.200 278.800 245.600 ;
        RECT 289.200 242.200 290.000 250.000 ;
        RECT 290.600 249.600 291.200 251.400 ;
        RECT 291.800 250.800 292.600 251.000 ;
        RECT 291.800 250.200 318.800 250.800 ;
        RECT 314.600 250.000 315.400 250.200 ;
        RECT 318.000 249.600 318.800 250.200 ;
        RECT 290.600 249.000 299.600 249.600 ;
        RECT 290.600 247.400 291.200 249.000 ;
        RECT 298.800 248.800 299.600 249.000 ;
        RECT 302.000 249.000 310.600 249.600 ;
        RECT 302.000 248.800 302.800 249.000 ;
        RECT 293.800 247.600 296.400 248.400 ;
        RECT 290.600 246.800 293.200 247.400 ;
        RECT 292.400 242.200 293.200 246.800 ;
        RECT 295.600 242.200 296.400 247.600 ;
        RECT 297.000 246.800 301.200 247.600 ;
        RECT 298.800 242.200 299.600 245.000 ;
        RECT 300.400 242.200 301.200 245.000 ;
        RECT 302.000 242.200 302.800 245.000 ;
        RECT 303.600 242.200 304.400 248.400 ;
        RECT 306.800 247.600 309.400 248.400 ;
        RECT 310.000 248.200 310.600 249.000 ;
        RECT 311.600 249.400 312.400 249.600 ;
        RECT 311.600 249.000 317.000 249.400 ;
        RECT 311.600 248.800 317.800 249.000 ;
        RECT 316.400 248.200 317.800 248.800 ;
        RECT 310.000 247.600 315.800 248.200 ;
        RECT 318.800 248.000 320.400 248.800 ;
        RECT 318.800 247.600 319.400 248.000 ;
        RECT 306.800 242.200 307.600 247.000 ;
        RECT 310.000 242.200 310.800 247.000 ;
        RECT 315.200 246.800 319.400 247.600 ;
        RECT 321.200 247.400 322.000 253.000 ;
        RECT 322.800 250.200 323.600 250.400 ;
        RECT 324.800 250.200 325.400 253.600 ;
        RECT 326.000 252.300 326.800 253.200 ;
        RECT 326.000 251.700 329.900 252.300 ;
        RECT 326.000 251.600 326.800 251.700 ;
        RECT 329.300 250.400 329.900 251.700 ;
        RECT 329.200 250.200 330.000 250.400 ;
        RECT 331.200 250.200 331.800 253.600 ;
        RECT 322.800 249.600 324.200 250.200 ;
        RECT 324.800 249.600 325.800 250.200 ;
        RECT 329.200 249.600 330.600 250.200 ;
        RECT 331.200 249.600 332.200 250.200 ;
        RECT 323.600 248.400 324.200 249.600 ;
        RECT 323.600 247.600 324.400 248.400 ;
        RECT 320.000 246.800 322.000 247.400 ;
        RECT 311.600 242.200 312.400 245.000 ;
        RECT 313.200 242.200 314.000 245.000 ;
        RECT 316.400 242.200 317.200 246.800 ;
        RECT 320.000 246.200 320.600 246.800 ;
        RECT 319.600 245.600 320.600 246.200 ;
        RECT 319.600 242.200 320.400 245.600 ;
        RECT 325.000 242.200 325.800 249.600 ;
        RECT 330.000 248.400 330.600 249.600 ;
        RECT 330.000 247.600 330.800 248.400 ;
        RECT 331.400 242.200 332.200 249.600 ;
        RECT 337.200 242.200 338.000 259.800 ;
        RECT 340.400 255.600 341.200 257.200 ;
        RECT 338.800 253.600 339.600 255.200 ;
        RECT 342.000 254.300 342.800 259.800 ;
        RECT 343.600 256.000 344.400 259.800 ;
        RECT 346.800 256.000 347.600 259.800 ;
        RECT 343.600 255.800 347.600 256.000 ;
        RECT 348.400 255.800 349.200 259.800 ;
        RECT 343.800 255.400 347.400 255.800 ;
        RECT 344.400 254.400 345.200 254.800 ;
        RECT 348.400 254.400 349.000 255.800 ;
        RECT 343.600 254.300 345.200 254.400 ;
        RECT 342.000 253.800 345.200 254.300 ;
        RECT 342.000 253.700 344.400 253.800 ;
        RECT 342.000 242.200 342.800 253.700 ;
        RECT 343.600 253.600 344.400 253.700 ;
        RECT 346.600 253.600 349.200 254.400 ;
        RECT 350.000 253.800 350.800 259.800 ;
        RECT 356.400 256.600 357.200 259.800 ;
        RECT 358.000 257.000 358.800 259.800 ;
        RECT 359.600 257.000 360.400 259.800 ;
        RECT 361.200 257.000 362.000 259.800 ;
        RECT 364.400 257.000 365.200 259.800 ;
        RECT 367.600 257.000 368.400 259.800 ;
        RECT 369.200 257.000 370.000 259.800 ;
        RECT 370.800 257.000 371.600 259.800 ;
        RECT 372.400 257.000 373.200 259.800 ;
        RECT 354.600 255.800 357.200 256.600 ;
        RECT 374.000 256.600 374.800 259.800 ;
        RECT 360.600 255.800 365.200 256.400 ;
        RECT 354.600 255.200 355.400 255.800 ;
        RECT 352.400 254.400 355.400 255.200 ;
        RECT 345.200 251.600 346.000 253.200 ;
        RECT 346.600 250.200 347.200 253.600 ;
        RECT 350.000 253.000 358.800 253.800 ;
        RECT 360.600 253.400 361.400 255.800 ;
        RECT 364.400 255.600 365.200 255.800 ;
        RECT 366.000 255.600 367.600 256.400 ;
        RECT 370.600 255.600 371.600 256.400 ;
        RECT 374.000 255.800 376.400 256.600 ;
        RECT 362.800 253.600 363.600 255.200 ;
        RECT 364.400 254.800 365.200 255.000 ;
        RECT 364.400 254.200 368.800 254.800 ;
        RECT 368.000 254.000 368.800 254.200 ;
        RECT 348.400 250.200 349.200 250.400 ;
        RECT 346.200 249.600 347.200 250.200 ;
        RECT 347.800 249.600 349.200 250.200 ;
        RECT 346.200 242.200 347.000 249.600 ;
        RECT 347.800 248.400 348.400 249.600 ;
        RECT 347.600 247.600 348.400 248.400 ;
        RECT 350.000 247.400 350.800 253.000 ;
        RECT 359.400 252.600 361.400 253.400 ;
        RECT 365.200 252.600 368.400 253.400 ;
        RECT 370.800 252.800 371.600 255.600 ;
        RECT 375.600 255.200 376.400 255.800 ;
        RECT 375.600 254.600 377.400 255.200 ;
        RECT 376.600 253.400 377.400 254.600 ;
        RECT 380.400 254.600 381.200 259.800 ;
        RECT 382.000 256.000 382.800 259.800 ;
        RECT 382.000 255.200 383.000 256.000 ;
        RECT 380.400 254.000 381.600 254.600 ;
        RECT 376.600 252.600 380.400 253.400 ;
        RECT 351.400 252.000 352.200 252.200 ;
        RECT 354.800 252.000 355.600 252.400 ;
        RECT 356.400 252.000 357.200 252.400 ;
        RECT 362.800 252.000 363.600 252.400 ;
        RECT 374.000 252.000 374.800 252.600 ;
        RECT 381.000 252.000 381.600 254.000 ;
        RECT 351.400 251.400 374.800 252.000 ;
        RECT 380.800 251.400 381.600 252.000 ;
        RECT 380.800 249.600 381.400 251.400 ;
        RECT 382.200 250.800 383.000 255.200 ;
        RECT 359.600 249.400 360.400 249.600 ;
        RECT 355.000 249.000 360.400 249.400 ;
        RECT 354.200 248.800 360.400 249.000 ;
        RECT 361.400 249.000 370.000 249.600 ;
        RECT 351.600 248.000 353.200 248.800 ;
        RECT 354.200 248.200 355.600 248.800 ;
        RECT 361.400 248.200 362.000 249.000 ;
        RECT 369.200 248.800 370.000 249.000 ;
        RECT 372.400 249.000 381.400 249.600 ;
        RECT 372.400 248.800 373.200 249.000 ;
        RECT 352.600 247.600 353.200 248.000 ;
        RECT 356.200 247.600 362.000 248.200 ;
        RECT 362.600 247.600 365.200 248.400 ;
        RECT 350.000 246.800 352.000 247.400 ;
        RECT 352.600 246.800 356.800 247.600 ;
        RECT 351.400 246.200 352.000 246.800 ;
        RECT 351.400 245.600 352.400 246.200 ;
        RECT 351.600 242.200 352.400 245.600 ;
        RECT 354.800 242.200 355.600 246.800 ;
        RECT 358.000 242.200 358.800 245.000 ;
        RECT 359.600 242.200 360.400 245.000 ;
        RECT 361.200 242.200 362.000 247.000 ;
        RECT 364.400 242.200 365.200 247.000 ;
        RECT 367.600 242.200 368.400 248.400 ;
        RECT 375.600 247.600 378.200 248.400 ;
        RECT 370.800 246.800 375.000 247.600 ;
        RECT 369.200 242.200 370.000 245.000 ;
        RECT 370.800 242.200 371.600 245.000 ;
        RECT 372.400 242.200 373.200 245.000 ;
        RECT 375.600 242.200 376.400 247.600 ;
        RECT 380.800 247.400 381.400 249.000 ;
        RECT 378.800 246.800 381.400 247.400 ;
        RECT 382.000 250.000 383.000 250.800 ;
        RECT 382.000 248.300 382.800 250.000 ;
        RECT 383.600 248.300 384.400 248.400 ;
        RECT 382.000 247.700 384.400 248.300 ;
        RECT 378.800 242.200 379.600 246.800 ;
        RECT 382.000 242.200 382.800 247.700 ;
        RECT 383.600 247.600 384.400 247.700 ;
        RECT 385.200 242.200 386.000 259.800 ;
        RECT 386.800 256.300 387.600 257.200 ;
        RECT 388.400 256.300 389.200 256.400 ;
        RECT 390.000 256.300 390.800 259.800 ;
        RECT 386.800 255.700 390.800 256.300 ;
        RECT 386.800 255.600 387.600 255.700 ;
        RECT 388.400 255.600 389.200 255.700 ;
        RECT 389.800 255.200 390.800 255.700 ;
        RECT 389.800 250.800 390.600 255.200 ;
        RECT 391.600 254.600 392.400 259.800 ;
        RECT 398.000 256.600 398.800 259.800 ;
        RECT 399.600 257.000 400.400 259.800 ;
        RECT 401.200 257.000 402.000 259.800 ;
        RECT 402.800 257.000 403.600 259.800 ;
        RECT 404.400 257.000 405.200 259.800 ;
        RECT 407.600 257.000 408.400 259.800 ;
        RECT 410.800 257.000 411.600 259.800 ;
        RECT 412.400 257.000 413.200 259.800 ;
        RECT 414.000 257.000 414.800 259.800 ;
        RECT 396.400 255.800 398.800 256.600 ;
        RECT 415.600 256.600 416.400 259.800 ;
        RECT 396.400 255.200 397.200 255.800 ;
        RECT 391.200 254.000 392.400 254.600 ;
        RECT 395.400 254.600 397.200 255.200 ;
        RECT 401.200 255.600 402.200 256.400 ;
        RECT 405.200 255.600 406.800 256.400 ;
        RECT 407.600 255.800 412.200 256.400 ;
        RECT 415.600 255.800 418.200 256.600 ;
        RECT 407.600 255.600 408.400 255.800 ;
        RECT 391.200 252.000 391.800 254.000 ;
        RECT 395.400 253.400 396.200 254.600 ;
        RECT 392.400 252.600 396.200 253.400 ;
        RECT 401.200 252.800 402.000 255.600 ;
        RECT 407.600 254.800 408.400 255.000 ;
        RECT 404.000 254.200 408.400 254.800 ;
        RECT 404.000 254.000 404.800 254.200 ;
        RECT 409.200 253.600 410.000 255.200 ;
        RECT 411.400 253.400 412.200 255.800 ;
        RECT 417.400 255.200 418.200 255.800 ;
        RECT 417.400 254.400 420.400 255.200 ;
        RECT 422.000 253.800 422.800 259.800 ;
        RECT 430.000 255.600 430.800 257.200 ;
        RECT 404.400 252.600 407.600 253.400 ;
        RECT 411.400 252.600 413.400 253.400 ;
        RECT 414.000 253.000 422.800 253.800 ;
        RECT 398.000 252.000 398.800 252.600 ;
        RECT 415.600 252.000 416.400 252.400 ;
        RECT 418.800 252.000 419.600 252.400 ;
        RECT 420.600 252.000 421.400 252.200 ;
        RECT 391.200 251.400 392.000 252.000 ;
        RECT 398.000 251.400 421.400 252.000 ;
        RECT 389.800 250.000 390.800 250.800 ;
        RECT 390.000 242.200 390.800 250.000 ;
        RECT 391.400 249.600 392.000 251.400 ;
        RECT 391.400 249.000 400.400 249.600 ;
        RECT 391.400 247.400 392.000 249.000 ;
        RECT 399.600 248.800 400.400 249.000 ;
        RECT 402.800 249.000 411.400 249.600 ;
        RECT 402.800 248.800 403.600 249.000 ;
        RECT 394.600 247.600 397.200 248.400 ;
        RECT 391.400 246.800 394.000 247.400 ;
        RECT 393.200 242.200 394.000 246.800 ;
        RECT 396.400 242.200 397.200 247.600 ;
        RECT 397.800 246.800 402.000 247.600 ;
        RECT 399.600 242.200 400.400 245.000 ;
        RECT 401.200 242.200 402.000 245.000 ;
        RECT 402.800 242.200 403.600 245.000 ;
        RECT 404.400 242.200 405.200 248.400 ;
        RECT 407.600 247.600 410.200 248.400 ;
        RECT 410.800 248.200 411.400 249.000 ;
        RECT 412.400 249.400 413.200 249.600 ;
        RECT 412.400 249.000 417.800 249.400 ;
        RECT 412.400 248.800 418.600 249.000 ;
        RECT 417.200 248.200 418.600 248.800 ;
        RECT 410.800 247.600 416.600 248.200 ;
        RECT 419.600 248.000 421.200 248.800 ;
        RECT 419.600 247.600 420.200 248.000 ;
        RECT 407.600 242.200 408.400 247.000 ;
        RECT 410.800 242.200 411.600 247.000 ;
        RECT 416.000 246.800 420.200 247.600 ;
        RECT 422.000 247.400 422.800 253.000 ;
        RECT 420.800 246.800 422.800 247.400 ;
        RECT 412.400 242.200 413.200 245.000 ;
        RECT 414.000 242.200 414.800 245.000 ;
        RECT 417.200 242.200 418.000 246.800 ;
        RECT 420.800 246.200 421.400 246.800 ;
        RECT 420.400 245.600 421.400 246.200 ;
        RECT 420.400 242.200 421.200 245.600 ;
        RECT 431.600 242.200 432.400 259.800 ;
        RECT 434.800 256.000 435.600 259.800 ;
        RECT 434.600 255.200 435.600 256.000 ;
        RECT 434.600 250.800 435.400 255.200 ;
        RECT 436.400 254.600 437.200 259.800 ;
        RECT 442.800 256.600 443.600 259.800 ;
        RECT 444.400 257.000 445.200 259.800 ;
        RECT 446.000 257.000 446.800 259.800 ;
        RECT 447.600 257.000 448.400 259.800 ;
        RECT 449.200 257.000 450.000 259.800 ;
        RECT 452.400 257.000 453.200 259.800 ;
        RECT 455.600 257.000 456.400 259.800 ;
        RECT 457.200 257.000 458.000 259.800 ;
        RECT 458.800 257.000 459.600 259.800 ;
        RECT 441.200 255.800 443.600 256.600 ;
        RECT 460.400 256.600 461.200 259.800 ;
        RECT 441.200 255.200 442.000 255.800 ;
        RECT 436.000 254.000 437.200 254.600 ;
        RECT 440.200 254.600 442.000 255.200 ;
        RECT 446.000 255.600 447.000 256.400 ;
        RECT 450.000 255.600 451.600 256.400 ;
        RECT 452.400 255.800 457.000 256.400 ;
        RECT 460.400 255.800 463.000 256.600 ;
        RECT 452.400 255.600 453.200 255.800 ;
        RECT 436.000 252.000 436.600 254.000 ;
        RECT 440.200 253.400 441.000 254.600 ;
        RECT 437.200 252.600 441.000 253.400 ;
        RECT 446.000 252.800 446.800 255.600 ;
        RECT 452.400 254.800 453.200 255.000 ;
        RECT 448.800 254.200 453.200 254.800 ;
        RECT 448.800 254.000 449.600 254.200 ;
        RECT 454.000 253.600 454.800 255.200 ;
        RECT 456.200 253.400 457.000 255.800 ;
        RECT 462.200 255.200 463.000 255.800 ;
        RECT 462.200 254.400 465.200 255.200 ;
        RECT 466.800 253.800 467.600 259.800 ;
        RECT 468.600 256.400 469.400 257.200 ;
        RECT 468.400 255.600 469.200 256.400 ;
        RECT 470.000 255.800 470.800 259.800 ;
        RECT 449.200 252.600 452.400 253.400 ;
        RECT 456.200 252.600 458.200 253.400 ;
        RECT 458.800 253.000 467.600 253.800 ;
        RECT 442.800 252.000 443.600 252.600 ;
        RECT 460.400 252.000 461.200 252.400 ;
        RECT 462.000 252.000 462.800 252.400 ;
        RECT 465.400 252.000 466.200 252.200 ;
        RECT 436.000 251.400 436.800 252.000 ;
        RECT 442.800 251.400 466.200 252.000 ;
        RECT 434.600 250.000 435.600 250.800 ;
        RECT 434.800 242.200 435.600 250.000 ;
        RECT 436.200 249.600 436.800 251.400 ;
        RECT 436.200 249.000 445.200 249.600 ;
        RECT 436.200 247.400 436.800 249.000 ;
        RECT 444.400 248.800 445.200 249.000 ;
        RECT 447.600 249.000 456.200 249.600 ;
        RECT 447.600 248.800 448.400 249.000 ;
        RECT 439.400 247.600 442.000 248.400 ;
        RECT 436.200 246.800 438.800 247.400 ;
        RECT 438.000 242.200 438.800 246.800 ;
        RECT 441.200 242.200 442.000 247.600 ;
        RECT 442.600 246.800 446.800 247.600 ;
        RECT 444.400 242.200 445.200 245.000 ;
        RECT 446.000 242.200 446.800 245.000 ;
        RECT 447.600 242.200 448.400 245.000 ;
        RECT 449.200 242.200 450.000 248.400 ;
        RECT 452.400 247.600 455.000 248.400 ;
        RECT 455.600 248.200 456.200 249.000 ;
        RECT 457.200 249.400 458.000 249.600 ;
        RECT 457.200 249.000 462.600 249.400 ;
        RECT 457.200 248.800 463.400 249.000 ;
        RECT 462.000 248.200 463.400 248.800 ;
        RECT 455.600 247.600 461.400 248.200 ;
        RECT 464.400 248.000 466.000 248.800 ;
        RECT 464.400 247.600 465.000 248.000 ;
        RECT 452.400 242.200 453.200 247.000 ;
        RECT 455.600 242.200 456.400 247.000 ;
        RECT 460.800 246.800 465.000 247.600 ;
        RECT 466.800 247.400 467.600 253.000 ;
        RECT 470.200 252.400 470.800 255.800 ;
        RECT 476.400 257.800 477.200 259.800 ;
        RECT 476.400 254.400 477.000 257.800 ;
        RECT 478.000 255.600 478.800 257.200 ;
        RECT 471.600 252.800 472.400 254.400 ;
        RECT 476.400 253.600 477.200 254.400 ;
        RECT 479.600 253.800 480.400 259.800 ;
        RECT 486.000 256.600 486.800 259.800 ;
        RECT 487.600 257.000 488.400 259.800 ;
        RECT 489.200 257.000 490.000 259.800 ;
        RECT 490.800 257.000 491.600 259.800 ;
        RECT 494.000 257.000 494.800 259.800 ;
        RECT 497.200 257.000 498.000 259.800 ;
        RECT 498.800 257.000 499.600 259.800 ;
        RECT 500.400 257.000 501.200 259.800 ;
        RECT 502.000 257.000 502.800 259.800 ;
        RECT 484.200 255.800 486.800 256.600 ;
        RECT 503.600 256.600 504.400 259.800 ;
        RECT 490.200 255.800 494.800 256.400 ;
        RECT 484.200 255.200 485.000 255.800 ;
        RECT 482.000 254.400 485.000 255.200 ;
        RECT 468.400 252.200 469.200 252.400 ;
        RECT 470.000 252.200 470.800 252.400 ;
        RECT 473.200 252.200 474.000 252.400 ;
        RECT 468.400 251.600 470.800 252.200 ;
        RECT 472.400 251.600 474.000 252.200 ;
        RECT 468.600 250.200 469.200 251.600 ;
        RECT 472.400 251.200 473.200 251.600 ;
        RECT 474.800 250.800 475.600 252.400 ;
        RECT 476.400 250.200 477.000 253.600 ;
        RECT 479.600 253.000 488.400 253.800 ;
        RECT 490.200 253.400 491.000 255.800 ;
        RECT 494.000 255.600 494.800 255.800 ;
        RECT 495.600 255.600 497.200 256.400 ;
        RECT 500.200 255.600 501.200 256.400 ;
        RECT 503.600 255.800 506.000 256.600 ;
        RECT 492.400 253.600 493.200 255.200 ;
        RECT 494.000 254.800 494.800 255.000 ;
        RECT 494.000 254.200 498.400 254.800 ;
        RECT 497.600 254.000 498.400 254.200 ;
        RECT 465.600 246.800 467.600 247.400 ;
        RECT 457.200 242.200 458.000 245.000 ;
        RECT 458.800 242.200 459.600 245.000 ;
        RECT 462.000 242.200 462.800 246.800 ;
        RECT 465.600 246.200 466.200 246.800 ;
        RECT 465.200 245.600 466.200 246.200 ;
        RECT 465.200 242.200 466.000 245.600 ;
        RECT 468.400 242.200 469.200 250.200 ;
        RECT 470.000 249.600 474.000 250.200 ;
        RECT 470.000 242.200 470.800 249.600 ;
        RECT 473.200 242.200 474.000 249.600 ;
        RECT 475.400 249.400 477.200 250.200 ;
        RECT 475.400 242.200 476.200 249.400 ;
        RECT 479.600 247.400 480.400 253.000 ;
        RECT 489.000 252.600 491.000 253.400 ;
        RECT 494.800 252.600 498.000 253.400 ;
        RECT 500.400 252.800 501.200 255.600 ;
        RECT 505.200 255.200 506.000 255.800 ;
        RECT 505.200 254.600 507.000 255.200 ;
        RECT 506.200 253.400 507.000 254.600 ;
        RECT 510.000 254.600 510.800 259.800 ;
        RECT 511.600 256.000 512.400 259.800 ;
        RECT 511.600 255.200 512.600 256.000 ;
        RECT 510.000 254.000 511.200 254.600 ;
        RECT 506.200 252.600 510.000 253.400 ;
        RECT 481.000 252.000 481.800 252.200 ;
        RECT 482.800 252.000 483.600 252.400 ;
        RECT 486.000 252.000 486.800 252.400 ;
        RECT 503.600 252.000 504.400 252.600 ;
        RECT 510.600 252.000 511.200 254.000 ;
        RECT 481.000 251.400 504.400 252.000 ;
        RECT 510.400 251.400 511.200 252.000 ;
        RECT 510.400 249.600 511.000 251.400 ;
        RECT 511.800 250.800 512.600 255.200 ;
        RECT 516.400 255.200 517.200 259.800 ;
        RECT 519.600 255.200 520.400 259.800 ;
        RECT 522.800 255.200 523.600 259.800 ;
        RECT 526.000 255.200 526.800 259.800 ;
        RECT 529.200 255.400 530.000 259.800 ;
        RECT 533.400 258.400 534.600 259.800 ;
        RECT 533.400 257.800 534.800 258.400 ;
        RECT 538.000 257.800 538.800 259.800 ;
        RECT 542.400 258.400 543.200 259.800 ;
        RECT 542.400 257.800 544.400 258.400 ;
        RECT 534.000 257.000 534.800 257.800 ;
        RECT 538.200 257.200 538.800 257.800 ;
        RECT 538.200 256.600 541.000 257.200 ;
        RECT 540.200 256.400 541.000 256.600 ;
        RECT 542.000 256.400 542.800 257.200 ;
        RECT 543.600 257.000 544.400 257.800 ;
        RECT 532.200 255.400 533.000 255.600 ;
        RECT 516.400 254.400 518.200 255.200 ;
        RECT 519.600 254.400 521.800 255.200 ;
        RECT 522.800 254.400 525.000 255.200 ;
        RECT 526.000 254.400 528.400 255.200 ;
        RECT 517.400 253.800 518.200 254.400 ;
        RECT 521.000 253.800 521.800 254.400 ;
        RECT 524.200 253.800 525.000 254.400 ;
        RECT 517.400 253.000 520.000 253.800 ;
        RECT 521.000 253.000 523.400 253.800 ;
        RECT 524.200 253.000 526.800 253.800 ;
        RECT 517.400 251.600 518.200 253.000 ;
        RECT 521.000 251.600 521.800 253.000 ;
        RECT 524.200 251.600 525.000 253.000 ;
        RECT 527.600 251.600 528.400 254.400 ;
        RECT 489.200 249.400 490.000 249.600 ;
        RECT 484.600 249.000 490.000 249.400 ;
        RECT 483.800 248.800 490.000 249.000 ;
        RECT 491.000 249.000 499.600 249.600 ;
        RECT 481.200 248.000 482.800 248.800 ;
        RECT 483.800 248.200 485.200 248.800 ;
        RECT 491.000 248.200 491.600 249.000 ;
        RECT 498.800 248.800 499.600 249.000 ;
        RECT 502.000 249.000 511.000 249.600 ;
        RECT 502.000 248.800 502.800 249.000 ;
        RECT 482.200 247.600 482.800 248.000 ;
        RECT 485.800 247.600 491.600 248.200 ;
        RECT 492.200 247.600 494.800 248.400 ;
        RECT 479.600 246.800 481.600 247.400 ;
        RECT 482.200 246.800 486.400 247.600 ;
        RECT 481.000 246.200 481.600 246.800 ;
        RECT 481.000 245.600 482.000 246.200 ;
        RECT 481.200 242.200 482.000 245.600 ;
        RECT 484.400 242.200 485.200 246.800 ;
        RECT 487.600 242.200 488.400 245.000 ;
        RECT 489.200 242.200 490.000 245.000 ;
        RECT 490.800 242.200 491.600 247.000 ;
        RECT 494.000 242.200 494.800 247.000 ;
        RECT 497.200 242.200 498.000 248.400 ;
        RECT 505.200 247.600 507.800 248.400 ;
        RECT 500.400 246.800 504.600 247.600 ;
        RECT 498.800 242.200 499.600 245.000 ;
        RECT 500.400 242.200 501.200 245.000 ;
        RECT 502.000 242.200 502.800 245.000 ;
        RECT 505.200 242.200 506.000 247.600 ;
        RECT 510.400 247.400 511.000 249.000 ;
        RECT 508.400 246.800 511.000 247.400 ;
        RECT 511.600 250.000 512.600 250.800 ;
        RECT 516.400 250.800 518.200 251.600 ;
        RECT 519.600 250.800 521.800 251.600 ;
        RECT 522.800 250.800 525.000 251.600 ;
        RECT 526.000 250.800 528.400 251.600 ;
        RECT 529.200 254.800 533.000 255.400 ;
        RECT 529.200 251.400 530.000 254.800 ;
        RECT 536.200 254.200 537.000 254.400 ;
        RECT 542.000 254.200 542.600 256.400 ;
        RECT 546.800 255.000 547.600 259.800 ;
        RECT 545.200 254.200 546.800 254.400 ;
        RECT 535.800 253.600 546.800 254.200 ;
        RECT 534.000 252.800 534.800 253.000 ;
        RECT 531.000 252.200 534.800 252.800 ;
        RECT 535.800 252.400 536.400 253.600 ;
        RECT 543.000 253.400 543.800 253.600 ;
        RECT 542.000 252.400 542.800 252.600 ;
        RECT 544.600 252.400 545.400 252.600 ;
        RECT 531.000 252.000 531.800 252.200 ;
        RECT 535.600 251.600 536.400 252.400 ;
        RECT 540.400 251.800 545.400 252.400 ;
        RECT 540.400 251.600 541.200 251.800 ;
        RECT 532.600 251.400 533.400 251.600 ;
        RECT 529.200 250.800 533.400 251.400 ;
        RECT 508.400 242.200 509.200 246.800 ;
        RECT 511.600 242.200 512.400 250.000 ;
        RECT 516.400 242.200 517.200 250.800 ;
        RECT 519.600 242.200 520.400 250.800 ;
        RECT 522.800 242.200 523.600 250.800 ;
        RECT 526.000 242.200 526.800 250.800 ;
        RECT 529.200 242.200 530.000 250.800 ;
        RECT 532.400 249.600 533.200 250.800 ;
        RECT 535.800 250.400 536.400 251.600 ;
        RECT 542.000 251.000 547.600 251.200 ;
        RECT 541.800 250.800 547.600 251.000 ;
        RECT 534.000 249.800 536.400 250.400 ;
        RECT 537.800 250.600 547.600 250.800 ;
        RECT 537.800 250.200 542.600 250.600 ;
        RECT 534.000 248.800 534.600 249.800 ;
        RECT 533.200 248.000 534.600 248.800 ;
        RECT 536.200 249.000 537.000 249.200 ;
        RECT 537.800 249.000 538.400 250.200 ;
        RECT 536.200 248.400 538.400 249.000 ;
        RECT 539.000 249.000 544.400 249.600 ;
        RECT 539.000 248.800 539.800 249.000 ;
        RECT 543.600 248.800 544.400 249.000 ;
        RECT 537.400 247.400 538.200 247.600 ;
        RECT 540.200 247.400 541.000 247.600 ;
        RECT 534.000 246.200 534.800 247.000 ;
        RECT 537.400 246.800 541.000 247.400 ;
        RECT 538.200 246.200 538.800 246.800 ;
        RECT 543.600 246.200 544.400 247.000 ;
        RECT 533.400 242.200 534.600 246.200 ;
        RECT 538.000 242.200 538.800 246.200 ;
        RECT 542.400 245.600 544.400 246.200 ;
        RECT 542.400 242.200 543.200 245.600 ;
        RECT 546.800 242.200 547.600 250.600 ;
        RECT 2.800 232.000 3.600 239.800 ;
        RECT 6.000 235.200 6.800 239.800 ;
        RECT 2.600 231.200 3.600 232.000 ;
        RECT 4.200 234.600 6.800 235.200 ;
        RECT 4.200 233.000 4.800 234.600 ;
        RECT 9.200 234.400 10.000 239.800 ;
        RECT 12.400 237.000 13.200 239.800 ;
        RECT 14.000 237.000 14.800 239.800 ;
        RECT 15.600 237.000 16.400 239.800 ;
        RECT 10.600 234.400 14.800 235.200 ;
        RECT 7.400 233.600 10.000 234.400 ;
        RECT 17.200 233.600 18.000 239.800 ;
        RECT 20.400 235.000 21.200 239.800 ;
        RECT 23.600 235.000 24.400 239.800 ;
        RECT 25.200 237.000 26.000 239.800 ;
        RECT 26.800 237.000 27.600 239.800 ;
        RECT 30.000 235.200 30.800 239.800 ;
        RECT 33.200 236.400 34.000 239.800 ;
        RECT 33.200 235.800 34.200 236.400 ;
        RECT 38.000 235.800 38.800 239.800 ;
        RECT 33.600 235.200 34.200 235.800 ;
        RECT 38.200 235.600 38.800 235.800 ;
        RECT 41.200 235.800 42.000 239.800 ;
        RECT 41.200 235.600 41.800 235.800 ;
        RECT 28.800 234.400 33.000 235.200 ;
        RECT 33.600 234.600 35.600 235.200 ;
        RECT 38.200 235.000 41.800 235.600 ;
        RECT 20.400 233.600 23.000 234.400 ;
        RECT 23.600 233.800 29.400 234.400 ;
        RECT 32.400 234.000 33.000 234.400 ;
        RECT 12.400 233.000 13.200 233.200 ;
        RECT 4.200 232.400 13.200 233.000 ;
        RECT 15.600 233.000 16.400 233.200 ;
        RECT 23.600 233.000 24.200 233.800 ;
        RECT 30.000 233.200 31.400 233.800 ;
        RECT 32.400 233.200 34.000 234.000 ;
        RECT 15.600 232.400 24.200 233.000 ;
        RECT 25.200 233.000 31.400 233.200 ;
        RECT 25.200 232.600 30.600 233.000 ;
        RECT 25.200 232.400 26.000 232.600 ;
        RECT 2.600 226.800 3.400 231.200 ;
        RECT 4.200 230.600 4.800 232.400 ;
        RECT 4.000 230.000 4.800 230.600 ;
        RECT 10.800 230.000 34.200 230.600 ;
        RECT 4.000 228.000 4.600 230.000 ;
        RECT 10.800 229.400 11.600 230.000 ;
        RECT 28.400 229.600 29.200 230.000 ;
        RECT 33.400 229.800 34.200 230.000 ;
        RECT 5.200 228.600 9.000 229.400 ;
        RECT 4.000 227.400 5.200 228.000 ;
        RECT 2.600 226.000 3.600 226.800 ;
        RECT 2.800 222.200 3.600 226.000 ;
        RECT 4.400 222.200 5.200 227.400 ;
        RECT 8.200 227.400 9.000 228.600 ;
        RECT 8.200 226.800 10.000 227.400 ;
        RECT 9.200 226.200 10.000 226.800 ;
        RECT 14.000 226.400 14.800 229.200 ;
        RECT 17.200 228.600 20.400 229.400 ;
        RECT 24.200 228.600 26.200 229.400 ;
        RECT 34.800 229.000 35.600 234.600 ;
        RECT 39.600 232.800 40.400 234.400 ;
        RECT 41.200 232.400 41.800 235.000 ;
        RECT 45.400 232.400 47.400 239.800 ;
        RECT 36.400 230.800 37.200 232.400 ;
        RECT 41.200 231.600 42.000 232.400 ;
        RECT 44.400 231.800 47.400 232.400 ;
        RECT 51.400 232.600 52.200 239.800 ;
        RECT 51.400 231.800 53.200 232.600 ;
        RECT 55.600 231.800 56.400 239.800 ;
        RECT 58.800 235.800 59.600 239.800 ;
        RECT 44.400 231.600 46.600 231.800 ;
        RECT 38.000 229.600 39.600 230.400 ;
        RECT 16.800 227.800 17.600 228.000 ;
        RECT 16.800 227.200 21.200 227.800 ;
        RECT 20.400 227.000 21.200 227.200 ;
        RECT 22.000 226.800 22.800 228.400 ;
        RECT 9.200 225.400 11.600 226.200 ;
        RECT 14.000 225.600 15.000 226.400 ;
        RECT 18.000 225.600 19.600 226.400 ;
        RECT 20.400 226.200 21.200 226.400 ;
        RECT 24.200 226.200 25.000 228.600 ;
        RECT 26.800 228.200 35.600 229.000 ;
        RECT 41.200 228.400 41.800 231.600 ;
        RECT 44.400 228.800 45.200 230.400 ;
        RECT 46.000 228.400 46.600 231.600 ;
        RECT 47.600 228.800 48.400 230.400 ;
        RECT 50.800 229.600 51.600 231.200 ;
        RECT 40.200 228.200 41.800 228.400 ;
        RECT 30.200 226.800 33.200 227.600 ;
        RECT 30.200 226.200 31.000 226.800 ;
        RECT 20.400 225.600 25.000 226.200 ;
        RECT 10.800 222.200 11.600 225.400 ;
        RECT 28.400 225.400 31.000 226.200 ;
        RECT 12.400 222.200 13.200 225.000 ;
        RECT 14.000 222.200 14.800 225.000 ;
        RECT 15.600 222.200 16.400 225.000 ;
        RECT 17.200 222.200 18.000 225.000 ;
        RECT 20.400 222.200 21.200 225.000 ;
        RECT 23.600 222.200 24.400 225.000 ;
        RECT 25.200 222.200 26.000 225.000 ;
        RECT 26.800 222.200 27.600 225.000 ;
        RECT 28.400 222.200 29.200 225.400 ;
        RECT 34.800 222.200 35.600 228.200 ;
        RECT 40.000 227.800 41.800 228.200 ;
        RECT 42.800 228.200 43.600 228.400 ;
        RECT 46.000 228.200 46.800 228.400 ;
        RECT 40.000 224.400 40.800 227.800 ;
        RECT 42.800 227.600 44.400 228.200 ;
        RECT 46.000 227.600 48.400 228.200 ;
        RECT 49.200 227.600 50.000 229.200 ;
        RECT 52.400 228.400 53.000 231.800 ;
        RECT 55.600 230.400 56.200 231.800 ;
        RECT 58.800 231.600 59.400 235.800 ;
        RECT 62.000 231.600 62.800 233.200 ;
        RECT 57.000 231.000 59.400 231.600 ;
        RECT 55.600 229.600 56.400 230.400 ;
        RECT 50.800 228.300 51.600 228.400 ;
        RECT 52.400 228.300 53.200 228.400 ;
        RECT 50.800 227.700 53.200 228.300 ;
        RECT 50.800 227.600 51.600 227.700 ;
        RECT 52.400 227.600 53.200 227.700 ;
        RECT 43.600 227.200 44.400 227.600 ;
        RECT 43.000 226.200 46.600 226.600 ;
        RECT 47.800 226.200 48.400 227.600 ;
        RECT 39.600 223.600 40.800 224.400 ;
        RECT 40.000 222.200 40.800 223.600 ;
        RECT 42.800 226.000 46.800 226.200 ;
        RECT 42.800 222.200 43.600 226.000 ;
        RECT 46.000 222.800 46.800 226.000 ;
        RECT 47.600 223.400 48.400 226.200 ;
        RECT 49.200 222.800 50.000 226.200 ;
        RECT 46.000 222.200 50.000 222.800 ;
        RECT 52.400 224.200 53.000 227.600 ;
        RECT 54.000 224.800 54.800 226.400 ;
        RECT 55.600 226.200 56.200 229.600 ;
        RECT 57.000 227.600 57.600 231.000 ;
        RECT 58.800 229.600 59.600 230.400 ;
        RECT 58.800 228.800 59.400 229.600 ;
        RECT 58.400 228.200 59.400 228.800 ;
        RECT 58.400 228.000 59.200 228.200 ;
        RECT 60.400 227.600 61.200 229.200 ;
        RECT 56.800 227.400 57.600 227.600 ;
        RECT 56.800 227.000 59.800 227.400 ;
        RECT 56.800 226.800 61.000 227.000 ;
        RECT 59.200 226.400 61.000 226.800 ;
        RECT 63.600 226.400 64.400 239.800 ;
        RECT 66.800 235.800 67.600 239.800 ;
        RECT 67.000 235.600 67.600 235.800 ;
        RECT 70.000 235.800 70.800 239.800 ;
        RECT 74.800 235.800 75.600 239.800 ;
        RECT 70.000 235.600 70.700 235.800 ;
        RECT 67.000 235.000 70.700 235.600 ;
        RECT 67.000 232.400 67.600 235.000 ;
        RECT 68.400 232.800 69.200 234.400 ;
        RECT 70.100 234.300 70.700 235.000 ;
        RECT 71.600 234.300 72.400 234.400 ;
        RECT 70.100 233.700 72.400 234.300 ;
        RECT 71.600 233.600 72.400 233.700 ;
        RECT 66.800 231.600 67.600 232.400 ;
        RECT 67.000 228.400 67.600 231.600 ;
        RECT 71.600 230.800 72.400 232.400 ;
        RECT 75.000 231.600 75.600 235.800 ;
        RECT 78.000 231.800 78.800 239.800 ;
        RECT 79.600 231.800 80.400 239.800 ;
        RECT 81.200 232.400 82.000 239.800 ;
        RECT 84.400 232.400 85.200 239.800 ;
        RECT 88.600 232.600 89.400 239.800 ;
        RECT 92.400 235.800 93.200 239.800 ;
        RECT 81.200 231.800 85.200 232.400 ;
        RECT 87.600 231.800 89.400 232.600 ;
        RECT 75.000 231.000 77.400 231.600 ;
        RECT 69.200 229.600 70.800 230.400 ;
        RECT 74.800 229.600 75.600 230.400 ;
        RECT 65.200 226.800 66.000 228.400 ;
        RECT 67.000 228.200 68.600 228.400 ;
        RECT 67.000 227.800 68.800 228.200 ;
        RECT 60.400 226.200 61.000 226.400 ;
        RECT 55.600 225.200 57.000 226.200 ;
        RECT 56.200 224.400 57.000 225.200 ;
        RECT 52.400 222.200 53.200 224.200 ;
        RECT 55.600 223.600 57.000 224.400 ;
        RECT 56.200 222.200 57.000 223.600 ;
        RECT 60.400 222.200 61.200 226.200 ;
        RECT 62.000 225.600 64.400 226.400 ;
        RECT 62.600 222.200 63.400 225.600 ;
        RECT 68.000 224.400 68.800 227.800 ;
        RECT 73.200 227.600 74.000 229.200 ;
        RECT 75.000 228.800 75.600 229.600 ;
        RECT 75.000 228.200 76.000 228.800 ;
        RECT 75.200 228.000 76.000 228.200 ;
        RECT 76.800 227.600 77.400 231.000 ;
        RECT 78.200 230.400 78.800 231.800 ;
        RECT 79.800 230.400 80.400 231.800 ;
        RECT 83.600 230.400 84.400 230.800 ;
        RECT 78.000 229.600 78.800 230.400 ;
        RECT 79.600 229.800 82.000 230.400 ;
        RECT 83.600 229.800 85.200 230.400 ;
        RECT 79.600 229.600 80.400 229.800 ;
        RECT 76.800 227.400 77.600 227.600 ;
        RECT 74.600 227.000 77.600 227.400 ;
        RECT 73.400 226.800 77.600 227.000 ;
        RECT 73.400 226.400 75.200 226.800 ;
        RECT 73.400 226.200 74.000 226.400 ;
        RECT 78.200 226.200 78.800 229.600 ;
        RECT 66.800 223.600 68.800 224.400 ;
        RECT 68.000 222.200 68.800 223.600 ;
        RECT 73.200 222.200 74.000 226.200 ;
        RECT 77.400 225.200 78.800 226.200 ;
        RECT 79.600 225.600 80.400 226.400 ;
        RECT 81.400 226.200 82.000 229.800 ;
        RECT 84.400 229.600 85.200 229.800 ;
        RECT 82.800 228.300 83.600 229.200 ;
        RECT 87.800 228.400 88.400 231.800 ;
        RECT 92.600 231.600 93.200 235.800 ;
        RECT 95.600 231.800 96.400 239.800 ;
        RECT 97.200 231.800 98.000 239.800 ;
        RECT 98.800 232.400 99.600 239.800 ;
        RECT 102.000 232.400 102.800 239.800 ;
        RECT 98.800 231.800 102.800 232.400 ;
        RECT 105.200 232.000 106.000 239.800 ;
        RECT 108.400 235.200 109.200 239.800 ;
        RECT 89.200 229.600 90.000 231.200 ;
        RECT 92.600 231.000 95.000 231.600 ;
        RECT 92.400 229.600 93.200 230.400 ;
        RECT 87.600 228.300 88.400 228.400 ;
        RECT 82.800 227.700 88.400 228.300 ;
        RECT 89.300 228.300 89.900 229.600 ;
        RECT 90.800 228.300 91.600 229.200 ;
        RECT 89.300 227.700 91.600 228.300 ;
        RECT 92.600 228.800 93.200 229.600 ;
        RECT 92.600 228.200 93.600 228.800 ;
        RECT 92.800 228.000 93.600 228.200 ;
        RECT 82.800 227.600 83.600 227.700 ;
        RECT 87.600 227.600 88.400 227.700 ;
        RECT 90.800 227.600 91.600 227.700 ;
        RECT 94.400 227.600 95.000 231.000 ;
        RECT 95.800 230.400 96.400 231.800 ;
        RECT 97.400 230.400 98.000 231.800 ;
        RECT 105.000 231.200 106.000 232.000 ;
        RECT 106.600 234.600 109.200 235.200 ;
        RECT 106.600 233.000 107.200 234.600 ;
        RECT 111.600 234.400 112.400 239.800 ;
        RECT 114.800 237.000 115.600 239.800 ;
        RECT 116.400 237.000 117.200 239.800 ;
        RECT 118.000 237.000 118.800 239.800 ;
        RECT 113.000 234.400 117.200 235.200 ;
        RECT 109.800 233.600 112.400 234.400 ;
        RECT 119.600 233.600 120.400 239.800 ;
        RECT 122.800 235.000 123.600 239.800 ;
        RECT 126.000 235.000 126.800 239.800 ;
        RECT 127.600 237.000 128.400 239.800 ;
        RECT 129.200 237.000 130.000 239.800 ;
        RECT 132.400 235.200 133.200 239.800 ;
        RECT 135.600 236.400 136.400 239.800 ;
        RECT 135.600 235.800 136.600 236.400 ;
        RECT 136.000 235.200 136.600 235.800 ;
        RECT 131.200 234.400 135.400 235.200 ;
        RECT 136.000 234.600 138.000 235.200 ;
        RECT 122.800 233.600 125.400 234.400 ;
        RECT 126.000 233.800 131.800 234.400 ;
        RECT 134.800 234.000 135.400 234.400 ;
        RECT 114.800 233.000 115.600 233.200 ;
        RECT 106.600 232.400 115.600 233.000 ;
        RECT 118.000 233.000 118.800 233.200 ;
        RECT 126.000 233.000 126.600 233.800 ;
        RECT 132.400 233.200 133.800 233.800 ;
        RECT 134.800 233.200 136.400 234.000 ;
        RECT 118.000 232.400 126.600 233.000 ;
        RECT 127.600 233.000 133.800 233.200 ;
        RECT 127.600 232.600 133.000 233.000 ;
        RECT 127.600 232.400 128.400 232.600 ;
        RECT 101.200 230.400 102.000 230.800 ;
        RECT 95.600 229.600 96.400 230.400 ;
        RECT 97.200 229.800 99.600 230.400 ;
        RECT 101.200 229.800 102.800 230.400 ;
        RECT 97.200 229.600 98.000 229.800 ;
        RECT 77.400 222.200 78.200 225.200 ;
        RECT 79.800 224.800 80.600 225.600 ;
        RECT 81.200 222.200 82.000 226.200 ;
        RECT 86.000 224.800 86.800 226.400 ;
        RECT 87.800 224.200 88.400 227.600 ;
        RECT 94.400 227.400 95.200 227.600 ;
        RECT 92.200 227.000 95.200 227.400 ;
        RECT 91.000 226.800 95.200 227.000 ;
        RECT 91.000 226.400 92.800 226.800 ;
        RECT 91.000 226.200 91.600 226.400 ;
        RECT 95.800 226.200 96.400 229.600 ;
        RECT 87.600 222.200 88.400 224.200 ;
        RECT 90.800 222.200 91.600 226.200 ;
        RECT 95.000 225.200 96.400 226.200 ;
        RECT 97.200 225.600 98.000 226.400 ;
        RECT 99.000 226.200 99.600 229.800 ;
        RECT 102.000 229.600 102.800 229.800 ;
        RECT 100.400 227.600 101.200 229.200 ;
        RECT 95.000 224.400 95.800 225.200 ;
        RECT 97.400 224.800 98.200 225.600 ;
        RECT 95.000 223.600 96.400 224.400 ;
        RECT 95.000 222.200 95.800 223.600 ;
        RECT 98.800 222.200 99.600 226.200 ;
        RECT 105.000 226.800 105.800 231.200 ;
        RECT 106.600 230.600 107.200 232.400 ;
        RECT 106.400 230.000 107.200 230.600 ;
        RECT 113.200 230.000 136.600 230.600 ;
        RECT 106.400 228.000 107.000 230.000 ;
        RECT 113.200 229.400 114.000 230.000 ;
        RECT 130.800 229.600 131.600 230.000 ;
        RECT 134.000 229.600 134.800 230.000 ;
        RECT 135.800 229.800 136.600 230.000 ;
        RECT 107.600 228.600 111.400 229.400 ;
        RECT 106.400 227.400 107.600 228.000 ;
        RECT 105.000 226.000 106.000 226.800 ;
        RECT 105.200 222.200 106.000 226.000 ;
        RECT 106.800 222.200 107.600 227.400 ;
        RECT 110.600 227.400 111.400 228.600 ;
        RECT 110.600 226.800 112.400 227.400 ;
        RECT 111.600 226.200 112.400 226.800 ;
        RECT 116.400 226.400 117.200 229.200 ;
        RECT 119.600 228.600 122.800 229.400 ;
        RECT 126.600 228.600 128.600 229.400 ;
        RECT 137.200 229.000 138.000 234.600 ;
        RECT 119.200 227.800 120.000 228.000 ;
        RECT 119.200 227.200 123.600 227.800 ;
        RECT 122.800 227.000 123.600 227.200 ;
        RECT 124.400 226.800 125.200 228.400 ;
        RECT 111.600 225.400 114.000 226.200 ;
        RECT 116.400 225.600 117.400 226.400 ;
        RECT 120.400 225.600 122.000 226.400 ;
        RECT 122.800 226.200 123.600 226.400 ;
        RECT 126.600 226.200 127.400 228.600 ;
        RECT 129.200 228.200 138.000 229.000 ;
        RECT 132.600 226.800 135.600 227.600 ;
        RECT 132.600 226.200 133.400 226.800 ;
        RECT 122.800 225.600 127.400 226.200 ;
        RECT 113.200 222.200 114.000 225.400 ;
        RECT 130.800 225.400 133.400 226.200 ;
        RECT 114.800 222.200 115.600 225.000 ;
        RECT 116.400 222.200 117.200 225.000 ;
        RECT 118.000 222.200 118.800 225.000 ;
        RECT 119.600 222.200 120.400 225.000 ;
        RECT 122.800 222.200 123.600 225.000 ;
        RECT 126.000 222.200 126.800 225.000 ;
        RECT 127.600 222.200 128.400 225.000 ;
        RECT 129.200 222.200 130.000 225.000 ;
        RECT 130.800 222.200 131.600 225.400 ;
        RECT 137.200 222.200 138.000 228.200 ;
        RECT 145.200 226.800 146.000 228.400 ;
        RECT 146.800 222.200 147.600 239.800 ;
        RECT 150.000 222.200 150.800 239.800 ;
        RECT 154.000 233.600 154.800 234.400 ;
        RECT 154.000 232.400 154.600 233.600 ;
        RECT 155.400 232.400 156.200 239.800 ;
        RECT 162.200 232.400 163.000 239.800 ;
        RECT 163.600 233.600 164.400 234.400 ;
        RECT 163.800 232.400 164.400 233.600 ;
        RECT 167.600 234.300 168.400 239.800 ;
        RECT 172.400 235.800 173.200 239.800 ;
        RECT 170.800 234.300 171.600 234.400 ;
        RECT 167.600 233.700 171.600 234.300 ;
        RECT 153.200 231.800 154.600 232.400 ;
        RECT 153.200 231.600 154.000 231.800 ;
        RECT 155.200 231.600 157.200 232.400 ;
        RECT 162.200 231.800 163.200 232.400 ;
        RECT 163.800 231.800 165.200 232.400 ;
        RECT 155.200 228.400 155.800 231.600 ;
        RECT 162.600 230.400 163.200 231.800 ;
        RECT 164.400 231.600 165.200 231.800 ;
        RECT 166.000 231.600 166.800 233.200 ;
        RECT 156.400 230.300 157.200 230.400 ;
        RECT 158.000 230.300 158.800 230.400 ;
        RECT 156.400 229.700 158.800 230.300 ;
        RECT 156.400 228.800 157.200 229.700 ;
        RECT 158.000 229.600 158.800 229.700 ;
        RECT 161.200 228.800 162.000 230.400 ;
        RECT 162.600 229.600 163.600 230.400 ;
        RECT 162.600 228.400 163.200 229.600 ;
        RECT 153.200 227.600 155.800 228.400 ;
        RECT 158.000 228.200 158.800 228.400 ;
        RECT 157.200 227.600 158.800 228.200 ;
        RECT 159.600 228.200 160.400 228.400 ;
        RECT 159.600 227.600 161.200 228.200 ;
        RECT 162.600 227.600 165.200 228.400 ;
        RECT 166.000 228.300 166.800 228.400 ;
        RECT 167.600 228.300 168.400 233.700 ;
        RECT 170.800 233.600 171.600 233.700 ;
        RECT 172.600 231.600 173.200 235.800 ;
        RECT 175.600 234.300 176.400 239.800 ;
        RECT 177.200 234.300 178.000 234.400 ;
        RECT 175.600 233.700 178.000 234.300 ;
        RECT 175.600 231.800 176.400 233.700 ;
        RECT 177.200 233.600 178.000 233.700 ;
        RECT 172.600 231.000 175.000 231.600 ;
        RECT 172.400 229.600 173.200 230.400 ;
        RECT 166.000 227.700 168.400 228.300 ;
        RECT 166.000 227.600 166.800 227.700 ;
        RECT 151.600 224.800 152.400 226.400 ;
        RECT 153.400 226.200 154.000 227.600 ;
        RECT 157.200 227.200 158.000 227.600 ;
        RECT 160.400 227.200 161.200 227.600 ;
        RECT 155.000 226.200 158.600 226.600 ;
        RECT 159.800 226.200 163.400 226.600 ;
        RECT 164.400 226.200 165.000 227.600 ;
        RECT 167.600 226.200 168.400 227.700 ;
        RECT 169.200 226.800 170.000 228.400 ;
        RECT 170.800 227.600 171.600 229.200 ;
        RECT 172.600 228.800 173.200 229.600 ;
        RECT 172.400 228.000 173.600 228.800 ;
        RECT 174.400 227.600 175.000 231.000 ;
        RECT 175.800 230.400 176.400 231.800 ;
        RECT 175.600 229.600 176.400 230.400 ;
        RECT 174.400 227.400 175.200 227.600 ;
        RECT 172.200 227.000 175.200 227.400 ;
        RECT 171.000 226.800 175.200 227.000 ;
        RECT 171.000 226.400 172.800 226.800 ;
        RECT 171.000 226.200 171.600 226.400 ;
        RECT 175.800 226.200 176.400 229.600 ;
        RECT 177.200 226.800 178.000 228.400 ;
        RECT 153.200 222.200 154.000 226.200 ;
        RECT 154.800 226.000 158.800 226.200 ;
        RECT 154.800 222.200 155.600 226.000 ;
        RECT 158.000 222.200 158.800 226.000 ;
        RECT 159.600 226.000 163.600 226.200 ;
        RECT 159.600 222.200 160.400 226.000 ;
        RECT 162.800 222.200 163.600 226.000 ;
        RECT 164.400 222.200 165.200 226.200 ;
        RECT 166.600 225.600 168.400 226.200 ;
        RECT 166.600 222.200 167.400 225.600 ;
        RECT 170.800 222.200 171.600 226.200 ;
        RECT 175.000 225.200 176.400 226.200 ;
        RECT 178.800 226.200 179.600 239.800 ;
        RECT 180.400 231.600 181.200 233.200 ;
        RECT 182.000 231.800 182.800 239.800 ;
        RECT 185.200 232.400 186.000 239.800 ;
        RECT 183.800 231.800 186.000 232.400 ;
        RECT 182.000 229.600 182.600 231.800 ;
        RECT 183.800 231.200 184.400 231.800 ;
        RECT 183.200 230.400 184.400 231.200 ;
        RECT 178.800 225.600 180.600 226.200 ;
        RECT 175.000 222.200 175.800 225.200 ;
        RECT 179.800 222.200 180.600 225.600 ;
        RECT 182.000 222.200 182.800 229.600 ;
        RECT 183.800 227.400 184.400 230.400 ;
        RECT 188.400 230.300 189.200 239.800 ;
        RECT 193.800 238.400 194.600 239.800 ;
        RECT 193.800 237.600 195.600 238.400 ;
        RECT 192.400 233.600 193.200 234.400 ;
        RECT 190.000 231.600 190.800 233.200 ;
        RECT 192.400 232.400 193.000 233.600 ;
        RECT 193.800 232.400 194.600 237.600 ;
        RECT 191.600 231.800 193.000 232.400 ;
        RECT 193.600 231.800 194.600 232.400 ;
        RECT 200.600 232.400 201.400 239.800 ;
        RECT 202.000 233.600 202.800 234.400 ;
        RECT 204.400 234.300 205.200 234.400 ;
        RECT 206.000 234.300 206.800 239.800 ;
        RECT 209.200 235.200 210.000 239.800 ;
        RECT 204.400 233.700 206.800 234.300 ;
        RECT 204.400 233.600 205.200 233.700 ;
        RECT 202.200 232.400 202.800 233.600 ;
        RECT 200.600 231.800 201.600 232.400 ;
        RECT 202.200 231.800 203.600 232.400 ;
        RECT 206.000 232.000 206.800 233.700 ;
        RECT 191.600 231.600 192.400 231.800 ;
        RECT 191.600 230.300 192.400 230.400 ;
        RECT 188.400 229.700 192.400 230.300 ;
        RECT 183.800 226.800 186.000 227.400 ;
        RECT 186.800 226.800 187.600 228.400 ;
        RECT 185.200 222.200 186.000 226.800 ;
        RECT 188.400 226.200 189.200 229.700 ;
        RECT 191.600 229.600 192.400 229.700 ;
        RECT 193.600 228.400 194.200 231.800 ;
        RECT 194.800 228.800 195.600 230.400 ;
        RECT 199.600 228.800 200.400 230.400 ;
        RECT 201.000 228.400 201.600 231.800 ;
        RECT 202.800 231.600 203.600 231.800 ;
        RECT 205.800 231.200 206.800 232.000 ;
        RECT 207.400 234.600 210.000 235.200 ;
        RECT 207.400 233.000 208.000 234.600 ;
        RECT 212.400 234.400 213.200 239.800 ;
        RECT 215.600 237.000 216.400 239.800 ;
        RECT 217.200 237.000 218.000 239.800 ;
        RECT 218.800 237.000 219.600 239.800 ;
        RECT 213.800 234.400 218.000 235.200 ;
        RECT 210.600 233.600 213.200 234.400 ;
        RECT 220.400 233.600 221.200 239.800 ;
        RECT 223.600 235.000 224.400 239.800 ;
        RECT 226.800 235.000 227.600 239.800 ;
        RECT 228.400 237.000 229.200 239.800 ;
        RECT 230.000 237.000 230.800 239.800 ;
        RECT 233.200 235.200 234.000 239.800 ;
        RECT 236.400 236.400 237.200 239.800 ;
        RECT 236.400 235.800 237.400 236.400 ;
        RECT 236.800 235.200 237.400 235.800 ;
        RECT 232.000 234.400 236.200 235.200 ;
        RECT 236.800 234.600 238.800 235.200 ;
        RECT 223.600 233.600 226.200 234.400 ;
        RECT 226.800 233.800 232.600 234.400 ;
        RECT 235.600 234.000 236.200 234.400 ;
        RECT 215.600 233.000 216.400 233.200 ;
        RECT 207.400 232.400 216.400 233.000 ;
        RECT 218.800 233.000 219.600 233.200 ;
        RECT 226.800 233.000 227.400 233.800 ;
        RECT 233.200 233.200 234.600 233.800 ;
        RECT 235.600 233.200 237.200 234.000 ;
        RECT 218.800 232.400 227.400 233.000 ;
        RECT 228.400 233.000 234.600 233.200 ;
        RECT 228.400 232.600 233.800 233.000 ;
        RECT 228.400 232.400 229.200 232.600 ;
        RECT 191.600 227.600 194.200 228.400 ;
        RECT 196.400 228.200 197.200 228.400 ;
        RECT 195.600 227.600 197.200 228.200 ;
        RECT 198.000 228.200 198.800 228.400 ;
        RECT 198.000 227.600 199.600 228.200 ;
        RECT 201.000 227.600 203.600 228.400 ;
        RECT 191.800 226.200 192.400 227.600 ;
        RECT 195.600 227.200 196.400 227.600 ;
        RECT 198.800 227.200 199.600 227.600 ;
        RECT 193.400 226.200 197.000 226.600 ;
        RECT 198.200 226.200 201.800 226.600 ;
        RECT 202.800 226.300 203.400 227.600 ;
        RECT 205.800 226.800 206.600 231.200 ;
        RECT 207.400 230.600 208.000 232.400 ;
        RECT 207.200 230.000 208.000 230.600 ;
        RECT 214.000 230.000 237.400 230.600 ;
        RECT 207.200 228.000 207.800 230.000 ;
        RECT 214.000 229.400 214.800 230.000 ;
        RECT 231.600 229.600 232.400 230.000 ;
        RECT 233.200 229.600 234.000 230.000 ;
        RECT 234.800 229.600 235.600 230.000 ;
        RECT 236.600 229.800 237.400 230.000 ;
        RECT 208.400 228.600 212.200 229.400 ;
        RECT 207.200 227.400 208.400 228.000 ;
        RECT 204.400 226.300 205.200 226.400 ;
        RECT 188.400 225.600 190.200 226.200 ;
        RECT 189.400 222.200 190.200 225.600 ;
        RECT 191.600 222.200 192.400 226.200 ;
        RECT 193.200 226.000 197.200 226.200 ;
        RECT 193.200 222.200 194.000 226.000 ;
        RECT 196.400 222.200 197.200 226.000 ;
        RECT 198.000 226.000 202.000 226.200 ;
        RECT 198.000 222.200 198.800 226.000 ;
        RECT 201.200 222.200 202.000 226.000 ;
        RECT 202.800 225.700 205.200 226.300 ;
        RECT 205.800 226.000 206.800 226.800 ;
        RECT 202.800 222.200 203.600 225.700 ;
        RECT 204.400 225.600 205.200 225.700 ;
        RECT 206.000 222.200 206.800 226.000 ;
        RECT 207.600 222.200 208.400 227.400 ;
        RECT 211.400 227.400 212.200 228.600 ;
        RECT 211.400 226.800 213.200 227.400 ;
        RECT 212.400 226.200 213.200 226.800 ;
        RECT 217.200 226.400 218.000 229.200 ;
        RECT 220.400 228.600 223.600 229.400 ;
        RECT 227.400 228.600 229.400 229.400 ;
        RECT 238.000 229.000 238.800 234.600 ;
        RECT 241.200 232.000 242.000 239.800 ;
        RECT 244.400 235.200 245.200 239.800 ;
        RECT 220.000 227.800 220.800 228.000 ;
        RECT 220.000 227.200 224.400 227.800 ;
        RECT 223.600 227.000 224.400 227.200 ;
        RECT 225.200 226.800 226.000 228.400 ;
        RECT 212.400 225.400 214.800 226.200 ;
        RECT 217.200 225.600 218.200 226.400 ;
        RECT 221.200 225.600 222.800 226.400 ;
        RECT 223.600 226.200 224.400 226.400 ;
        RECT 227.400 226.200 228.200 228.600 ;
        RECT 230.000 228.200 238.800 229.000 ;
        RECT 233.400 226.800 236.400 227.600 ;
        RECT 233.400 226.200 234.200 226.800 ;
        RECT 223.600 225.600 228.200 226.200 ;
        RECT 214.000 222.200 214.800 225.400 ;
        RECT 231.600 225.400 234.200 226.200 ;
        RECT 215.600 222.200 216.400 225.000 ;
        RECT 217.200 222.200 218.000 225.000 ;
        RECT 218.800 222.200 219.600 225.000 ;
        RECT 220.400 222.200 221.200 225.000 ;
        RECT 223.600 222.200 224.400 225.000 ;
        RECT 226.800 222.200 227.600 225.000 ;
        RECT 228.400 222.200 229.200 225.000 ;
        RECT 230.000 222.200 230.800 225.000 ;
        RECT 231.600 222.200 232.400 225.400 ;
        RECT 238.000 222.200 238.800 228.200 ;
        RECT 241.000 231.200 242.000 232.000 ;
        RECT 242.600 234.600 245.200 235.200 ;
        RECT 242.600 233.000 243.200 234.600 ;
        RECT 247.600 234.400 248.400 239.800 ;
        RECT 250.800 237.000 251.600 239.800 ;
        RECT 252.400 237.000 253.200 239.800 ;
        RECT 254.000 237.000 254.800 239.800 ;
        RECT 249.000 234.400 253.200 235.200 ;
        RECT 245.800 233.600 248.400 234.400 ;
        RECT 255.600 233.600 256.400 239.800 ;
        RECT 258.800 235.000 259.600 239.800 ;
        RECT 262.000 235.000 262.800 239.800 ;
        RECT 263.600 237.000 264.400 239.800 ;
        RECT 265.200 237.000 266.000 239.800 ;
        RECT 268.400 235.200 269.200 239.800 ;
        RECT 271.600 236.400 272.400 239.800 ;
        RECT 271.600 235.800 272.600 236.400 ;
        RECT 272.000 235.200 272.600 235.800 ;
        RECT 267.200 234.400 271.400 235.200 ;
        RECT 272.000 234.600 274.000 235.200 ;
        RECT 258.800 233.600 261.400 234.400 ;
        RECT 262.000 233.800 267.800 234.400 ;
        RECT 270.800 234.000 271.400 234.400 ;
        RECT 250.800 233.000 251.600 233.200 ;
        RECT 242.600 232.400 251.600 233.000 ;
        RECT 254.000 233.000 254.800 233.200 ;
        RECT 262.000 233.000 262.600 233.800 ;
        RECT 268.400 233.200 269.800 233.800 ;
        RECT 270.800 233.200 272.400 234.000 ;
        RECT 254.000 232.400 262.600 233.000 ;
        RECT 263.600 233.000 269.800 233.200 ;
        RECT 263.600 232.600 269.000 233.000 ;
        RECT 263.600 232.400 264.400 232.600 ;
        RECT 241.000 226.800 241.800 231.200 ;
        RECT 242.600 230.600 243.200 232.400 ;
        RECT 242.400 230.000 243.200 230.600 ;
        RECT 249.200 230.000 272.600 230.600 ;
        RECT 242.400 228.000 243.000 230.000 ;
        RECT 249.200 229.400 250.000 230.000 ;
        RECT 266.800 229.600 267.600 230.000 ;
        RECT 270.000 229.600 270.800 230.000 ;
        RECT 271.800 229.800 272.600 230.000 ;
        RECT 243.600 228.600 247.400 229.400 ;
        RECT 242.400 227.400 243.600 228.000 ;
        RECT 239.600 226.300 240.400 226.400 ;
        RECT 241.000 226.300 242.000 226.800 ;
        RECT 239.600 225.700 242.000 226.300 ;
        RECT 239.600 225.600 240.400 225.700 ;
        RECT 241.200 222.200 242.000 225.700 ;
        RECT 242.800 222.200 243.600 227.400 ;
        RECT 246.600 227.400 247.400 228.600 ;
        RECT 246.600 226.800 248.400 227.400 ;
        RECT 247.600 226.200 248.400 226.800 ;
        RECT 252.400 226.400 253.200 229.200 ;
        RECT 255.600 228.600 258.800 229.400 ;
        RECT 262.600 228.600 264.600 229.400 ;
        RECT 273.200 229.000 274.000 234.600 ;
        RECT 255.200 227.800 256.000 228.000 ;
        RECT 255.200 227.200 259.600 227.800 ;
        RECT 258.800 227.000 259.600 227.200 ;
        RECT 260.400 226.800 261.200 228.400 ;
        RECT 247.600 225.400 250.000 226.200 ;
        RECT 252.400 225.600 253.400 226.400 ;
        RECT 256.400 225.600 258.000 226.400 ;
        RECT 258.800 226.200 259.600 226.400 ;
        RECT 262.600 226.200 263.400 228.600 ;
        RECT 265.200 228.200 274.000 229.000 ;
        RECT 268.600 226.800 271.600 227.600 ;
        RECT 268.600 226.200 269.400 226.800 ;
        RECT 258.800 225.600 263.400 226.200 ;
        RECT 249.200 222.200 250.000 225.400 ;
        RECT 266.800 225.400 269.400 226.200 ;
        RECT 250.800 222.200 251.600 225.000 ;
        RECT 252.400 222.200 253.200 225.000 ;
        RECT 254.000 222.200 254.800 225.000 ;
        RECT 255.600 222.200 256.400 225.000 ;
        RECT 258.800 222.200 259.600 225.000 ;
        RECT 262.000 222.200 262.800 225.000 ;
        RECT 263.600 222.200 264.400 225.000 ;
        RECT 265.200 222.200 266.000 225.000 ;
        RECT 266.800 222.200 267.600 225.400 ;
        RECT 273.200 222.200 274.000 228.200 ;
        RECT 276.400 226.300 277.200 226.400 ;
        RECT 281.200 226.300 282.000 226.400 ;
        RECT 276.400 225.700 282.000 226.300 ;
        RECT 276.400 225.600 277.200 225.700 ;
        RECT 281.200 224.800 282.000 225.700 ;
        RECT 282.800 222.200 283.600 239.800 ;
        RECT 286.000 232.000 286.800 239.800 ;
        RECT 289.200 235.200 290.000 239.800 ;
        RECT 285.800 231.200 286.800 232.000 ;
        RECT 287.400 234.600 290.000 235.200 ;
        RECT 287.400 233.000 288.000 234.600 ;
        RECT 292.400 234.400 293.200 239.800 ;
        RECT 295.600 237.000 296.400 239.800 ;
        RECT 297.200 237.000 298.000 239.800 ;
        RECT 298.800 237.000 299.600 239.800 ;
        RECT 293.800 234.400 298.000 235.200 ;
        RECT 290.600 233.600 293.200 234.400 ;
        RECT 300.400 233.600 301.200 239.800 ;
        RECT 303.600 235.000 304.400 239.800 ;
        RECT 306.800 235.000 307.600 239.800 ;
        RECT 308.400 237.000 309.200 239.800 ;
        RECT 310.000 237.000 310.800 239.800 ;
        RECT 313.200 235.200 314.000 239.800 ;
        RECT 316.400 236.400 317.200 239.800 ;
        RECT 322.200 238.400 323.000 239.800 ;
        RECT 321.200 237.600 323.000 238.400 ;
        RECT 316.400 235.800 317.400 236.400 ;
        RECT 316.800 235.200 317.400 235.800 ;
        RECT 312.000 234.400 316.200 235.200 ;
        RECT 316.800 234.600 318.800 235.200 ;
        RECT 303.600 233.600 306.200 234.400 ;
        RECT 306.800 233.800 312.600 234.400 ;
        RECT 315.600 234.000 316.200 234.400 ;
        RECT 295.600 233.000 296.400 233.200 ;
        RECT 287.400 232.400 296.400 233.000 ;
        RECT 298.800 233.000 299.600 233.200 ;
        RECT 306.800 233.000 307.400 233.800 ;
        RECT 313.200 233.200 314.600 233.800 ;
        RECT 315.600 233.200 317.200 234.000 ;
        RECT 298.800 232.400 307.400 233.000 ;
        RECT 308.400 233.000 314.600 233.200 ;
        RECT 308.400 232.600 313.800 233.000 ;
        RECT 308.400 232.400 309.200 232.600 ;
        RECT 285.800 226.800 286.600 231.200 ;
        RECT 287.400 230.600 288.000 232.400 ;
        RECT 311.400 231.800 312.400 232.000 ;
        RECT 314.800 231.800 315.600 232.400 ;
        RECT 288.600 231.200 315.600 231.800 ;
        RECT 288.600 231.000 289.400 231.200 ;
        RECT 287.200 230.000 288.000 230.600 ;
        RECT 287.200 228.000 287.800 230.000 ;
        RECT 288.400 228.600 292.200 229.400 ;
        RECT 287.200 227.400 288.400 228.000 ;
        RECT 285.800 226.000 286.800 226.800 ;
        RECT 286.000 222.200 286.800 226.000 ;
        RECT 287.600 222.200 288.400 227.400 ;
        RECT 291.400 227.400 292.200 228.600 ;
        RECT 291.400 226.800 293.200 227.400 ;
        RECT 292.400 226.200 293.200 226.800 ;
        RECT 297.200 226.400 298.000 229.200 ;
        RECT 300.400 228.600 303.600 229.400 ;
        RECT 307.400 228.600 309.400 229.400 ;
        RECT 318.000 229.000 318.800 234.600 ;
        RECT 322.200 232.400 323.000 237.600 ;
        RECT 323.600 233.600 324.400 234.400 ;
        RECT 323.800 232.400 324.400 233.600 ;
        RECT 328.600 232.400 329.400 239.800 ;
        RECT 330.000 233.600 330.800 234.400 ;
        RECT 330.200 232.400 330.800 233.600 ;
        RECT 333.200 233.600 334.000 234.400 ;
        RECT 333.200 232.400 333.800 233.600 ;
        RECT 334.600 232.400 335.400 239.800 ;
        RECT 339.600 233.600 340.400 234.400 ;
        RECT 339.600 232.400 340.200 233.600 ;
        RECT 341.000 232.400 341.800 239.800 ;
        RECT 322.200 231.800 323.200 232.400 ;
        RECT 323.800 231.800 325.200 232.400 ;
        RECT 328.600 231.800 329.600 232.400 ;
        RECT 330.200 231.800 331.600 232.400 ;
        RECT 300.000 227.800 300.800 228.000 ;
        RECT 300.000 227.200 304.400 227.800 ;
        RECT 303.600 227.000 304.400 227.200 ;
        RECT 305.200 226.800 306.000 228.400 ;
        RECT 292.400 225.400 294.800 226.200 ;
        RECT 297.200 225.600 298.200 226.400 ;
        RECT 301.200 225.600 302.800 226.400 ;
        RECT 303.600 226.200 304.400 226.400 ;
        RECT 307.400 226.200 308.200 228.600 ;
        RECT 310.000 228.200 318.800 229.000 ;
        RECT 321.200 228.800 322.000 230.400 ;
        RECT 322.600 228.400 323.200 231.800 ;
        RECT 324.400 231.600 325.200 231.800 ;
        RECT 327.600 228.800 328.400 230.400 ;
        RECT 329.000 228.400 329.600 231.800 ;
        RECT 330.800 231.600 331.600 231.800 ;
        RECT 332.400 231.800 333.800 232.400 ;
        RECT 334.400 231.800 335.400 232.400 ;
        RECT 338.800 231.800 340.200 232.400 ;
        RECT 340.800 231.800 341.800 232.400 ;
        RECT 345.200 231.800 346.000 239.800 ;
        RECT 348.400 232.400 349.200 239.800 ;
        RECT 347.000 231.800 349.200 232.400 ;
        RECT 350.000 232.400 350.800 239.800 ;
        RECT 350.000 231.800 352.200 232.400 ;
        RECT 353.200 231.800 354.000 239.800 ;
        RECT 357.400 238.400 358.200 239.800 ;
        RECT 356.400 237.600 358.200 238.400 ;
        RECT 357.400 232.400 358.200 237.600 ;
        RECT 358.800 233.600 359.600 234.400 ;
        RECT 359.000 232.400 359.600 233.600 ;
        RECT 357.400 231.800 358.400 232.400 ;
        RECT 359.000 231.800 360.400 232.400 ;
        RECT 332.400 231.600 333.200 231.800 ;
        RECT 334.400 228.400 335.000 231.800 ;
        RECT 338.800 231.600 339.600 231.800 ;
        RECT 337.200 230.300 338.000 230.400 ;
        RECT 340.800 230.300 341.400 231.800 ;
        RECT 337.200 229.700 341.400 230.300 ;
        RECT 337.200 229.600 338.000 229.700 ;
        RECT 340.800 228.400 341.400 229.700 ;
        RECT 345.200 229.600 345.800 231.800 ;
        RECT 347.000 231.200 347.600 231.800 ;
        RECT 346.400 230.400 347.600 231.200 ;
        RECT 313.400 226.800 316.400 227.600 ;
        RECT 313.400 226.200 314.200 226.800 ;
        RECT 303.600 225.600 308.200 226.200 ;
        RECT 294.000 222.200 294.800 225.400 ;
        RECT 311.600 225.400 314.200 226.200 ;
        RECT 295.600 222.200 296.400 225.000 ;
        RECT 297.200 222.200 298.000 225.000 ;
        RECT 298.800 222.200 299.600 225.000 ;
        RECT 300.400 222.200 301.200 225.000 ;
        RECT 303.600 222.200 304.400 225.000 ;
        RECT 306.800 222.200 307.600 225.000 ;
        RECT 308.400 222.200 309.200 225.000 ;
        RECT 310.000 222.200 310.800 225.000 ;
        RECT 311.600 222.200 312.400 225.400 ;
        RECT 318.000 222.200 318.800 228.200 ;
        RECT 319.600 228.200 320.400 228.400 ;
        RECT 319.600 227.600 321.200 228.200 ;
        RECT 322.600 227.600 325.200 228.400 ;
        RECT 326.000 228.200 326.800 228.400 ;
        RECT 326.000 227.600 327.600 228.200 ;
        RECT 329.000 227.600 331.600 228.400 ;
        RECT 332.400 227.600 335.000 228.400 ;
        RECT 337.200 228.200 338.000 228.400 ;
        RECT 336.400 227.600 338.000 228.200 ;
        RECT 338.800 227.600 341.400 228.400 ;
        RECT 343.600 228.300 344.400 228.400 ;
        RECT 345.200 228.300 346.000 229.600 ;
        RECT 343.600 228.200 346.000 228.300 ;
        RECT 342.800 227.700 346.000 228.200 ;
        RECT 342.800 227.600 344.400 227.700 ;
        RECT 320.400 227.200 321.200 227.600 ;
        RECT 319.800 226.200 323.400 226.600 ;
        RECT 324.400 226.200 325.000 227.600 ;
        RECT 326.800 227.200 327.600 227.600 ;
        RECT 326.200 226.200 329.800 226.600 ;
        RECT 330.800 226.200 331.400 227.600 ;
        RECT 332.600 226.200 333.200 227.600 ;
        RECT 336.400 227.200 337.200 227.600 ;
        RECT 334.200 226.200 337.800 226.600 ;
        RECT 339.000 226.200 339.600 227.600 ;
        RECT 342.800 227.200 343.600 227.600 ;
        RECT 340.600 226.200 344.200 226.600 ;
        RECT 319.600 226.000 323.600 226.200 ;
        RECT 319.600 222.200 320.400 226.000 ;
        RECT 322.800 222.200 323.600 226.000 ;
        RECT 324.400 222.200 325.200 226.200 ;
        RECT 326.000 226.000 330.000 226.200 ;
        RECT 326.000 222.200 326.800 226.000 ;
        RECT 329.200 222.200 330.000 226.000 ;
        RECT 330.800 222.200 331.600 226.200 ;
        RECT 332.400 222.200 333.200 226.200 ;
        RECT 334.000 226.000 338.000 226.200 ;
        RECT 334.000 222.200 334.800 226.000 ;
        RECT 337.200 222.200 338.000 226.000 ;
        RECT 338.800 222.200 339.600 226.200 ;
        RECT 340.400 226.000 344.400 226.200 ;
        RECT 340.400 222.200 341.200 226.000 ;
        RECT 343.600 222.200 344.400 226.000 ;
        RECT 345.200 222.200 346.000 227.700 ;
        RECT 347.000 227.400 347.600 230.400 ;
        RECT 351.600 231.200 352.200 231.800 ;
        RECT 351.600 230.400 352.800 231.200 ;
        RECT 351.600 227.400 352.200 230.400 ;
        RECT 353.400 229.600 354.000 231.800 ;
        RECT 347.000 226.800 349.200 227.400 ;
        RECT 348.400 222.200 349.200 226.800 ;
        RECT 350.000 226.800 352.200 227.400 ;
        RECT 350.000 222.200 350.800 226.800 ;
        RECT 353.200 222.200 354.000 229.600 ;
        RECT 356.400 228.800 357.200 230.400 ;
        RECT 357.800 228.400 358.400 231.800 ;
        RECT 359.600 231.600 360.400 231.800 ;
        RECT 361.200 231.800 362.000 239.800 ;
        RECT 364.400 232.400 365.200 239.800 ;
        RECT 366.800 233.600 367.600 234.400 ;
        RECT 366.800 232.400 367.400 233.600 ;
        RECT 368.200 232.400 369.000 239.800 ;
        RECT 363.000 231.800 365.200 232.400 ;
        RECT 366.000 231.800 367.400 232.400 ;
        RECT 368.000 231.800 369.000 232.400 ;
        RECT 361.200 229.600 361.800 231.800 ;
        RECT 363.000 231.200 363.600 231.800 ;
        RECT 366.000 231.600 366.800 231.800 ;
        RECT 362.400 230.400 363.600 231.200 ;
        RECT 368.000 230.400 368.600 231.800 ;
        RECT 354.800 228.200 355.600 228.400 ;
        RECT 354.800 227.600 356.400 228.200 ;
        RECT 357.800 227.600 360.400 228.400 ;
        RECT 355.600 227.200 356.400 227.600 ;
        RECT 355.000 226.200 358.600 226.600 ;
        RECT 359.600 226.200 360.200 227.600 ;
        RECT 354.800 226.000 358.800 226.200 ;
        RECT 354.800 222.200 355.600 226.000 ;
        RECT 358.000 222.200 358.800 226.000 ;
        RECT 359.600 222.200 360.400 226.200 ;
        RECT 361.200 222.200 362.000 229.600 ;
        RECT 363.000 227.400 363.600 230.400 ;
        RECT 367.600 229.600 368.600 230.400 ;
        RECT 368.000 228.400 368.600 229.600 ;
        RECT 374.000 230.300 374.800 239.800 ;
        RECT 375.600 231.600 376.400 233.200 ;
        RECT 378.800 232.000 379.600 239.800 ;
        RECT 382.000 235.200 382.800 239.800 ;
        RECT 378.600 231.200 379.600 232.000 ;
        RECT 380.200 234.600 382.800 235.200 ;
        RECT 380.200 233.000 380.800 234.600 ;
        RECT 385.200 234.400 386.000 239.800 ;
        RECT 388.400 237.000 389.200 239.800 ;
        RECT 390.000 237.000 390.800 239.800 ;
        RECT 391.600 237.000 392.400 239.800 ;
        RECT 386.600 234.400 390.800 235.200 ;
        RECT 383.400 233.600 386.000 234.400 ;
        RECT 393.200 233.600 394.000 239.800 ;
        RECT 396.400 235.000 397.200 239.800 ;
        RECT 399.600 235.000 400.400 239.800 ;
        RECT 401.200 237.000 402.000 239.800 ;
        RECT 402.800 237.000 403.600 239.800 ;
        RECT 406.000 235.200 406.800 239.800 ;
        RECT 409.200 236.400 410.000 239.800 ;
        RECT 409.200 235.800 410.200 236.400 ;
        RECT 409.600 235.200 410.200 235.800 ;
        RECT 404.800 234.400 409.000 235.200 ;
        RECT 409.600 234.600 411.600 235.200 ;
        RECT 396.400 233.600 399.000 234.400 ;
        RECT 399.600 233.800 405.400 234.400 ;
        RECT 408.400 234.000 409.000 234.400 ;
        RECT 388.400 233.000 389.200 233.200 ;
        RECT 380.200 232.400 389.200 233.000 ;
        RECT 391.600 233.000 392.400 233.200 ;
        RECT 399.600 233.000 400.200 233.800 ;
        RECT 406.000 233.200 407.400 233.800 ;
        RECT 408.400 233.200 410.000 234.000 ;
        RECT 391.600 232.400 400.200 233.000 ;
        RECT 401.200 233.000 407.400 233.200 ;
        RECT 401.200 232.600 406.600 233.000 ;
        RECT 401.200 232.400 402.000 232.600 ;
        RECT 377.200 230.300 378.000 230.400 ;
        RECT 374.000 229.700 378.000 230.300 ;
        RECT 366.000 227.600 368.600 228.400 ;
        RECT 370.800 228.200 371.600 228.400 ;
        RECT 370.000 227.600 371.600 228.200 ;
        RECT 363.000 226.800 365.200 227.400 ;
        RECT 364.400 222.200 365.200 226.800 ;
        RECT 366.200 226.200 366.800 227.600 ;
        RECT 370.000 227.200 370.800 227.600 ;
        RECT 367.800 226.200 371.400 226.600 ;
        RECT 374.000 226.200 374.800 229.700 ;
        RECT 377.200 229.600 378.000 229.700 ;
        RECT 378.600 226.800 379.400 231.200 ;
        RECT 380.200 230.600 380.800 232.400 ;
        RECT 380.000 230.000 380.800 230.600 ;
        RECT 386.800 230.000 410.200 230.600 ;
        RECT 380.000 228.000 380.600 230.000 ;
        RECT 386.800 229.400 387.600 230.000 ;
        RECT 404.400 229.600 405.200 230.000 ;
        RECT 409.400 229.800 410.200 230.000 ;
        RECT 381.200 228.600 385.000 229.400 ;
        RECT 380.000 227.400 381.200 228.000 ;
        RECT 366.000 222.200 366.800 226.200 ;
        RECT 367.600 226.000 371.600 226.200 ;
        RECT 367.600 222.200 368.400 226.000 ;
        RECT 370.800 222.200 371.600 226.000 ;
        RECT 374.000 225.600 375.800 226.200 ;
        RECT 378.600 226.000 379.600 226.800 ;
        RECT 375.000 222.200 375.800 225.600 ;
        RECT 378.800 222.200 379.600 226.000 ;
        RECT 380.400 222.200 381.200 227.400 ;
        RECT 384.200 227.400 385.000 228.600 ;
        RECT 384.200 226.800 386.000 227.400 ;
        RECT 385.200 226.200 386.000 226.800 ;
        RECT 390.000 226.400 390.800 229.200 ;
        RECT 393.200 228.600 396.400 229.400 ;
        RECT 400.200 228.600 402.200 229.400 ;
        RECT 410.800 229.000 411.600 234.600 ;
        RECT 392.800 227.800 393.600 228.000 ;
        RECT 392.800 227.200 397.200 227.800 ;
        RECT 396.400 227.000 397.200 227.200 ;
        RECT 398.000 226.800 398.800 228.400 ;
        RECT 385.200 225.400 387.600 226.200 ;
        RECT 390.000 225.600 391.000 226.400 ;
        RECT 394.000 225.600 395.600 226.400 ;
        RECT 396.400 226.200 397.200 226.400 ;
        RECT 400.200 226.200 401.000 228.600 ;
        RECT 402.800 228.200 411.600 229.000 ;
        RECT 406.200 226.800 409.200 227.600 ;
        RECT 406.200 226.200 407.000 226.800 ;
        RECT 396.400 225.600 401.000 226.200 ;
        RECT 386.800 222.200 387.600 225.400 ;
        RECT 404.400 225.400 407.000 226.200 ;
        RECT 388.400 222.200 389.200 225.000 ;
        RECT 390.000 222.200 390.800 225.000 ;
        RECT 391.600 222.200 392.400 225.000 ;
        RECT 393.200 222.200 394.000 225.000 ;
        RECT 396.400 222.200 397.200 225.000 ;
        RECT 399.600 222.200 400.400 225.000 ;
        RECT 401.200 222.200 402.000 225.000 ;
        RECT 402.800 222.200 403.600 225.000 ;
        RECT 404.400 222.200 405.200 225.400 ;
        RECT 410.800 222.200 411.600 228.200 ;
        RECT 414.000 228.300 414.800 239.800 ;
        RECT 418.200 232.400 419.000 239.800 ;
        RECT 430.000 235.600 430.800 239.800 ;
        RECT 433.200 235.800 434.000 239.800 ;
        RECT 433.200 235.600 433.800 235.800 ;
        RECT 430.200 235.000 433.800 235.600 ;
        RECT 419.600 233.600 420.400 234.400 ;
        RECT 422.000 234.300 422.800 234.400 ;
        RECT 431.600 234.300 432.400 234.400 ;
        RECT 422.000 233.700 432.400 234.300 ;
        RECT 422.000 233.600 422.800 233.700 ;
        RECT 419.800 232.400 420.400 233.600 ;
        RECT 431.600 232.800 432.400 233.700 ;
        RECT 433.200 232.400 433.800 235.000 ;
        RECT 435.400 232.600 436.200 239.800 ;
        RECT 441.200 235.800 442.000 239.800 ;
        RECT 441.400 235.600 442.000 235.800 ;
        RECT 444.400 235.800 445.200 239.800 ;
        RECT 444.400 235.600 445.000 235.800 ;
        RECT 441.400 235.000 445.000 235.600 ;
        RECT 439.600 234.300 440.400 234.400 ;
        RECT 442.800 234.300 443.600 234.400 ;
        RECT 439.600 233.700 443.600 234.300 ;
        RECT 439.600 233.600 440.400 233.700 ;
        RECT 442.800 232.800 443.600 233.700 ;
        RECT 418.200 231.800 419.200 232.400 ;
        RECT 419.800 232.300 421.200 232.400 ;
        RECT 426.800 232.300 427.600 232.400 ;
        RECT 419.800 231.800 427.600 232.300 ;
        RECT 417.200 228.800 418.000 230.400 ;
        RECT 418.600 228.400 419.200 231.800 ;
        RECT 420.400 231.700 427.600 231.800 ;
        RECT 420.400 231.600 421.200 231.700 ;
        RECT 426.800 231.600 427.600 231.700 ;
        RECT 428.400 230.800 429.200 232.400 ;
        RECT 433.200 231.600 434.000 232.400 ;
        RECT 435.400 231.800 437.200 232.600 ;
        RECT 444.400 232.400 445.000 235.000 ;
        RECT 439.600 232.300 440.400 232.400 ;
        RECT 441.200 232.300 442.000 232.400 ;
        RECT 430.000 229.600 431.600 230.400 ;
        RECT 433.200 228.400 433.800 231.600 ;
        RECT 434.800 229.600 435.600 231.200 ;
        RECT 436.400 230.400 437.000 231.800 ;
        RECT 439.600 231.700 442.000 232.300 ;
        RECT 439.600 230.800 440.400 231.700 ;
        RECT 441.200 231.600 442.000 231.700 ;
        RECT 444.400 231.600 445.200 232.400 ;
        RECT 446.000 232.300 446.800 232.400 ;
        RECT 447.600 232.300 448.400 239.800 ;
        RECT 446.000 231.700 448.400 232.300 ;
        RECT 446.000 231.600 446.800 231.700 ;
        RECT 436.400 229.600 437.200 230.400 ;
        RECT 441.200 229.600 442.800 230.400 ;
        RECT 415.600 228.300 416.400 228.400 ;
        RECT 414.000 228.200 416.400 228.300 ;
        RECT 414.000 227.700 417.200 228.200 ;
        RECT 412.400 224.800 413.200 226.400 ;
        RECT 414.000 222.200 414.800 227.700 ;
        RECT 415.600 227.600 417.200 227.700 ;
        RECT 418.600 227.600 421.200 228.400 ;
        RECT 432.200 228.200 433.800 228.400 ;
        RECT 432.000 227.800 433.800 228.200 ;
        RECT 436.400 228.400 437.000 229.600 ;
        RECT 444.400 228.400 445.000 231.600 ;
        RECT 416.400 227.200 417.200 227.600 ;
        RECT 415.800 226.200 419.400 226.600 ;
        RECT 420.400 226.200 421.000 227.600 ;
        RECT 415.600 226.000 419.600 226.200 ;
        RECT 415.600 222.200 416.400 226.000 ;
        RECT 418.800 222.200 419.600 226.000 ;
        RECT 420.400 222.200 421.200 226.200 ;
        RECT 432.000 222.200 432.800 227.800 ;
        RECT 436.400 227.600 437.200 228.400 ;
        RECT 443.400 228.200 445.000 228.400 ;
        RECT 443.200 227.800 445.000 228.200 ;
        RECT 436.400 224.200 437.000 227.600 ;
        RECT 438.000 224.800 438.800 226.400 ;
        RECT 436.400 222.200 437.200 224.200 ;
        RECT 443.200 222.200 444.000 227.800 ;
        RECT 446.000 226.800 446.800 228.400 ;
        RECT 447.600 226.200 448.400 231.700 ;
        RECT 449.200 231.600 450.000 233.200 ;
        RECT 453.400 232.400 454.200 239.800 ;
        RECT 458.800 235.800 459.600 239.800 ;
        RECT 459.000 235.600 459.600 235.800 ;
        RECT 462.000 235.800 462.800 239.800 ;
        RECT 465.200 235.800 466.000 239.800 ;
        RECT 462.000 235.600 462.600 235.800 ;
        RECT 459.000 235.000 462.600 235.600 ;
        RECT 465.400 235.600 466.000 235.800 ;
        RECT 468.400 235.800 469.200 239.800 ;
        RECT 468.400 235.600 469.000 235.800 ;
        RECT 465.400 235.000 469.000 235.600 ;
        RECT 454.800 233.600 455.600 234.400 ;
        RECT 455.000 232.400 455.600 233.600 ;
        RECT 460.400 232.800 461.200 234.400 ;
        RECT 462.000 232.400 462.600 235.000 ;
        RECT 466.800 232.800 467.600 234.400 ;
        RECT 468.400 232.400 469.000 235.000 ;
        RECT 472.600 232.600 473.400 239.800 ;
        RECT 477.400 232.600 478.200 239.800 ;
        RECT 453.400 231.800 454.400 232.400 ;
        RECT 455.000 231.800 456.400 232.400 ;
        RECT 453.800 230.400 454.400 231.800 ;
        RECT 455.600 231.600 456.400 231.800 ;
        RECT 457.200 230.800 458.000 232.400 ;
        RECT 462.000 231.600 462.800 232.400 ;
        RECT 452.400 228.800 453.200 230.400 ;
        RECT 453.800 229.600 454.800 230.400 ;
        RECT 458.800 229.600 460.400 230.400 ;
        RECT 453.800 228.400 454.400 229.600 ;
        RECT 462.000 228.400 462.600 231.600 ;
        RECT 463.600 230.800 464.400 232.400 ;
        RECT 468.400 231.600 469.200 232.400 ;
        RECT 471.600 231.800 473.400 232.600 ;
        RECT 476.400 231.800 478.200 232.600 ;
        RECT 479.600 232.400 480.400 239.800 ;
        RECT 482.800 232.400 483.600 239.800 ;
        RECT 479.600 231.800 483.600 232.400 ;
        RECT 484.400 231.800 485.200 239.800 ;
        RECT 465.200 229.600 466.800 230.400 ;
        RECT 468.400 228.400 469.000 231.600 ;
        RECT 471.800 228.400 472.400 231.800 ;
        RECT 476.400 231.600 477.200 231.800 ;
        RECT 473.200 229.600 474.000 231.200 ;
        RECT 476.600 228.400 477.200 231.600 ;
        RECT 478.000 229.600 478.800 231.200 ;
        RECT 480.400 230.400 481.200 230.800 ;
        RECT 484.400 230.400 485.000 231.800 ;
        RECT 479.600 229.800 481.200 230.400 ;
        RECT 482.800 229.800 485.200 230.400 ;
        RECT 479.600 229.600 480.400 229.800 ;
        RECT 450.800 228.200 451.600 228.400 ;
        RECT 450.800 227.600 452.400 228.200 ;
        RECT 453.800 227.600 456.400 228.400 ;
        RECT 461.000 228.200 462.600 228.400 ;
        RECT 467.400 228.200 469.000 228.400 ;
        RECT 460.800 227.800 462.600 228.200 ;
        RECT 467.200 227.800 469.000 228.200 ;
        RECT 470.000 228.300 470.800 228.400 ;
        RECT 471.600 228.300 472.400 228.400 ;
        RECT 451.600 227.200 452.400 227.600 ;
        RECT 451.000 226.200 454.600 226.600 ;
        RECT 455.600 226.200 456.200 227.600 ;
        RECT 447.600 225.600 449.400 226.200 ;
        RECT 448.600 222.200 449.400 225.600 ;
        RECT 450.800 226.000 454.800 226.200 ;
        RECT 450.800 222.200 451.600 226.000 ;
        RECT 454.000 222.200 454.800 226.000 ;
        RECT 455.600 222.200 456.400 226.200 ;
        RECT 460.800 222.200 461.600 227.800 ;
        RECT 467.200 222.200 468.000 227.800 ;
        RECT 470.000 227.700 472.400 228.300 ;
        RECT 470.000 227.600 470.800 227.700 ;
        RECT 471.600 227.600 472.400 227.700 ;
        RECT 476.400 227.600 477.200 228.400 ;
        RECT 479.600 228.300 480.400 228.400 ;
        RECT 481.200 228.300 482.000 229.200 ;
        RECT 479.600 227.700 482.000 228.300 ;
        RECT 479.600 227.600 480.400 227.700 ;
        RECT 481.200 227.600 482.000 227.700 ;
        RECT 470.000 224.800 470.800 226.400 ;
        RECT 471.800 224.200 472.400 227.600 ;
        RECT 474.800 224.800 475.600 226.400 ;
        RECT 476.600 224.200 477.200 227.600 ;
        RECT 471.600 222.200 472.400 224.200 ;
        RECT 476.400 222.200 477.200 224.200 ;
        RECT 482.800 226.200 483.400 229.800 ;
        RECT 484.400 229.600 485.200 229.800 ;
        RECT 482.800 222.200 483.600 226.200 ;
        RECT 484.400 225.600 485.200 226.400 ;
        RECT 487.600 226.200 488.400 239.800 ;
        RECT 489.200 232.300 490.000 233.200 ;
        RECT 490.800 232.300 491.600 233.200 ;
        RECT 489.200 231.700 491.600 232.300 ;
        RECT 489.200 231.600 490.000 231.700 ;
        RECT 490.800 231.600 491.600 231.700 ;
        RECT 492.400 226.200 493.200 239.800 ;
        RECT 497.200 232.000 498.000 239.800 ;
        RECT 500.400 235.200 501.200 239.800 ;
        RECT 487.600 225.600 489.400 226.200 ;
        RECT 484.200 224.800 485.000 225.600 ;
        RECT 488.600 222.200 489.400 225.600 ;
        RECT 491.400 225.600 493.200 226.200 ;
        RECT 497.000 231.200 498.000 232.000 ;
        RECT 498.600 234.600 501.200 235.200 ;
        RECT 498.600 233.000 499.200 234.600 ;
        RECT 503.600 234.400 504.400 239.800 ;
        RECT 506.800 237.000 507.600 239.800 ;
        RECT 508.400 237.000 509.200 239.800 ;
        RECT 510.000 237.000 510.800 239.800 ;
        RECT 505.000 234.400 509.200 235.200 ;
        RECT 501.800 233.600 504.400 234.400 ;
        RECT 511.600 233.600 512.400 239.800 ;
        RECT 514.800 235.000 515.600 239.800 ;
        RECT 518.000 235.000 518.800 239.800 ;
        RECT 519.600 237.000 520.400 239.800 ;
        RECT 521.200 237.000 522.000 239.800 ;
        RECT 524.400 235.200 525.200 239.800 ;
        RECT 527.600 236.400 528.400 239.800 ;
        RECT 527.600 235.800 528.600 236.400 ;
        RECT 528.000 235.200 528.600 235.800 ;
        RECT 523.200 234.400 527.400 235.200 ;
        RECT 528.000 234.600 530.000 235.200 ;
        RECT 514.800 233.600 517.400 234.400 ;
        RECT 518.000 233.800 523.800 234.400 ;
        RECT 526.800 234.000 527.400 234.400 ;
        RECT 506.800 233.000 507.600 233.200 ;
        RECT 498.600 232.400 507.600 233.000 ;
        RECT 510.000 233.000 510.800 233.200 ;
        RECT 518.000 233.000 518.600 233.800 ;
        RECT 524.400 233.200 525.800 233.800 ;
        RECT 526.800 233.200 528.400 234.000 ;
        RECT 510.000 232.400 518.600 233.000 ;
        RECT 519.600 233.000 525.800 233.200 ;
        RECT 519.600 232.600 525.000 233.000 ;
        RECT 519.600 232.400 520.400 232.600 ;
        RECT 497.000 226.800 497.800 231.200 ;
        RECT 498.600 230.600 499.200 232.400 ;
        RECT 498.400 230.000 499.200 230.600 ;
        RECT 505.200 230.000 528.600 230.600 ;
        RECT 498.400 228.000 499.000 230.000 ;
        RECT 505.200 229.400 506.000 230.000 ;
        RECT 522.800 229.600 523.600 230.000 ;
        RECT 527.800 229.800 528.600 230.000 ;
        RECT 499.600 228.600 503.400 229.400 ;
        RECT 498.400 227.400 499.600 228.000 ;
        RECT 497.000 226.000 498.000 226.800 ;
        RECT 491.400 224.400 492.200 225.600 ;
        RECT 490.800 223.600 492.200 224.400 ;
        RECT 491.400 222.200 492.200 223.600 ;
        RECT 497.200 222.200 498.000 226.000 ;
        RECT 498.800 222.200 499.600 227.400 ;
        RECT 502.600 227.400 503.400 228.600 ;
        RECT 502.600 226.800 504.400 227.400 ;
        RECT 503.600 226.200 504.400 226.800 ;
        RECT 508.400 226.400 509.200 229.200 ;
        RECT 511.600 228.600 514.800 229.400 ;
        RECT 518.600 228.600 520.600 229.400 ;
        RECT 529.200 229.000 530.000 234.600 ;
        RECT 530.800 231.800 531.600 239.800 ;
        RECT 532.400 232.400 533.200 239.800 ;
        RECT 535.600 232.400 536.400 239.800 ;
        RECT 532.400 231.800 536.400 232.400 ;
        RECT 531.000 230.400 531.600 231.800 ;
        RECT 537.200 231.600 538.000 233.200 ;
        RECT 530.800 229.800 533.200 230.400 ;
        RECT 530.800 229.600 531.600 229.800 ;
        RECT 511.200 227.800 512.000 228.000 ;
        RECT 511.200 227.200 515.600 227.800 ;
        RECT 514.800 227.000 515.600 227.200 ;
        RECT 516.400 226.800 517.200 228.400 ;
        RECT 503.600 225.400 506.000 226.200 ;
        RECT 508.400 225.600 509.400 226.400 ;
        RECT 512.400 225.600 514.000 226.400 ;
        RECT 514.800 226.200 515.600 226.400 ;
        RECT 518.600 226.200 519.400 228.600 ;
        RECT 521.200 228.200 530.000 229.000 ;
        RECT 524.600 226.800 527.600 227.600 ;
        RECT 524.600 226.200 525.400 226.800 ;
        RECT 514.800 225.600 519.400 226.200 ;
        RECT 505.200 222.200 506.000 225.400 ;
        RECT 522.800 225.400 525.400 226.200 ;
        RECT 506.800 222.200 507.600 225.000 ;
        RECT 508.400 222.200 509.200 225.000 ;
        RECT 510.000 222.200 510.800 225.000 ;
        RECT 511.600 222.200 512.400 225.000 ;
        RECT 514.800 222.200 515.600 225.000 ;
        RECT 518.000 222.200 518.800 225.000 ;
        RECT 519.600 222.200 520.400 225.000 ;
        RECT 521.200 222.200 522.000 225.000 ;
        RECT 522.800 222.200 523.600 225.400 ;
        RECT 529.200 222.200 530.000 228.200 ;
        RECT 530.800 225.600 531.600 226.400 ;
        RECT 532.600 226.200 533.200 229.800 ;
        RECT 534.000 228.300 534.800 229.200 ;
        RECT 537.200 228.300 538.000 228.400 ;
        RECT 534.000 227.700 538.000 228.300 ;
        RECT 534.000 227.600 534.800 227.700 ;
        RECT 537.200 227.600 538.000 227.700 ;
        RECT 538.800 226.200 539.600 239.800 ;
        RECT 544.600 232.600 545.400 239.800 ;
        RECT 543.600 231.800 545.400 232.600 ;
        RECT 546.800 232.400 547.600 239.800 ;
        RECT 546.800 231.800 549.000 232.400 ;
        RECT 542.000 230.300 542.800 230.400 ;
        RECT 543.800 230.300 544.400 231.800 ;
        RECT 548.400 231.200 549.000 231.800 ;
        RECT 542.000 229.700 544.400 230.300 ;
        RECT 542.000 229.600 542.800 229.700 ;
        RECT 543.800 228.400 544.400 229.700 ;
        RECT 545.200 229.600 546.000 231.200 ;
        RECT 548.400 230.400 549.600 231.200 ;
        RECT 546.800 228.800 547.600 230.400 ;
        RECT 543.600 227.600 544.400 228.400 ;
        RECT 531.000 224.800 531.800 225.600 ;
        RECT 532.400 222.200 533.200 226.200 ;
        RECT 537.800 225.600 539.600 226.200 ;
        RECT 537.800 224.400 538.600 225.600 ;
        RECT 542.000 224.800 542.800 226.400 ;
        RECT 537.200 223.600 538.600 224.400 ;
        RECT 543.800 224.200 544.400 227.600 ;
        RECT 548.400 227.400 549.000 230.400 ;
        RECT 537.800 222.200 538.600 223.600 ;
        RECT 543.600 222.200 544.400 224.200 ;
        RECT 546.800 226.800 549.000 227.400 ;
        RECT 546.800 222.200 547.600 226.800 ;
        RECT 2.800 212.300 3.600 219.800 ;
        RECT 7.600 217.800 8.400 219.800 ;
        RECT 6.000 215.600 6.800 217.200 ;
        RECT 4.400 213.600 5.200 215.200 ;
        RECT 7.800 214.400 8.400 217.800 ;
        RECT 13.800 218.400 15.400 219.800 ;
        RECT 13.800 217.600 16.400 218.400 ;
        RECT 13.800 215.800 15.400 217.600 ;
        RECT 19.400 216.400 20.200 219.800 ;
        RECT 19.400 215.800 21.200 216.400 ;
        RECT 7.600 214.300 8.400 214.400 ;
        RECT 7.600 213.700 11.500 214.300 ;
        RECT 7.600 213.600 8.400 213.700 ;
        RECT 6.000 212.300 6.800 212.400 ;
        RECT 2.800 211.700 6.800 212.300 ;
        RECT 2.800 202.200 3.600 211.700 ;
        RECT 6.000 211.600 6.800 211.700 ;
        RECT 7.800 210.200 8.400 213.600 ;
        RECT 10.900 212.400 11.500 213.700 ;
        RECT 12.400 212.800 13.200 214.400 ;
        RECT 14.200 212.400 14.800 215.800 ;
        RECT 15.600 214.300 16.400 214.400 ;
        RECT 17.200 214.300 18.000 214.400 ;
        RECT 15.600 213.700 18.000 214.300 ;
        RECT 15.600 213.600 16.400 213.700 ;
        RECT 17.200 213.600 18.000 213.700 ;
        RECT 18.800 214.300 19.600 214.400 ;
        RECT 20.400 214.300 21.200 215.800 ;
        RECT 18.800 213.700 21.200 214.300 ;
        RECT 18.800 213.600 19.600 213.700 ;
        RECT 15.600 213.200 16.200 213.600 ;
        RECT 15.400 212.400 16.200 213.200 ;
        RECT 9.200 210.800 10.000 212.400 ;
        RECT 10.800 212.200 11.600 212.400 ;
        RECT 10.800 211.600 12.400 212.200 ;
        RECT 14.000 211.600 14.800 212.400 ;
        RECT 11.600 211.200 12.400 211.600 ;
        RECT 14.200 211.400 14.800 211.600 ;
        RECT 14.200 210.800 16.200 211.400 ;
        RECT 17.200 210.800 18.000 212.400 ;
        RECT 15.600 210.200 16.200 210.800 ;
        RECT 7.600 209.400 9.400 210.200 ;
        RECT 8.600 202.200 9.400 209.400 ;
        RECT 10.800 209.600 14.800 210.200 ;
        RECT 10.800 202.200 11.600 209.600 ;
        RECT 14.000 202.800 14.800 209.600 ;
        RECT 15.600 203.400 16.400 210.200 ;
        RECT 17.200 202.800 18.000 210.200 ;
        RECT 18.800 208.800 19.600 210.400 ;
        RECT 14.000 202.200 18.000 202.800 ;
        RECT 20.400 202.200 21.200 213.700 ;
        RECT 22.000 213.600 22.800 215.200 ;
        RECT 24.800 214.200 25.600 219.800 ;
        RECT 30.000 215.800 30.800 219.800 ;
        RECT 34.200 216.800 35.000 219.800 ;
        RECT 34.200 215.800 35.600 216.800 ;
        RECT 36.400 215.800 37.200 219.800 ;
        RECT 40.600 216.800 41.400 219.800 ;
        RECT 40.600 215.800 42.000 216.800 ;
        RECT 30.200 215.600 30.800 215.800 ;
        RECT 30.200 215.200 32.000 215.600 ;
        RECT 30.200 215.000 34.400 215.200 ;
        RECT 31.400 214.600 34.400 215.000 ;
        RECT 33.600 214.400 34.400 214.600 ;
        RECT 23.800 213.800 25.600 214.200 ;
        RECT 23.800 213.600 25.400 213.800 ;
        RECT 23.800 210.400 24.400 213.600 ;
        RECT 30.000 212.800 30.800 214.400 ;
        RECT 32.000 213.800 32.800 214.000 ;
        RECT 31.800 213.200 32.800 213.800 ;
        RECT 31.800 212.400 32.400 213.200 ;
        RECT 26.000 211.600 27.600 212.400 ;
        RECT 31.600 211.600 32.400 212.400 ;
        RECT 23.600 209.600 24.400 210.400 ;
        RECT 28.400 209.600 29.200 211.200 ;
        RECT 33.600 211.000 34.200 214.400 ;
        RECT 35.000 212.400 35.600 215.800 ;
        RECT 36.600 215.600 37.200 215.800 ;
        RECT 36.600 215.200 38.400 215.600 ;
        RECT 36.600 215.000 40.800 215.200 ;
        RECT 37.800 214.600 40.800 215.000 ;
        RECT 40.000 214.400 40.800 214.600 ;
        RECT 36.400 212.800 37.200 214.400 ;
        RECT 38.400 213.800 39.200 214.000 ;
        RECT 38.200 213.200 39.200 213.800 ;
        RECT 38.200 212.400 38.800 213.200 ;
        RECT 34.800 211.600 35.600 212.400 ;
        RECT 38.000 211.600 38.800 212.400 ;
        RECT 31.800 210.400 34.200 211.000 ;
        RECT 23.800 207.000 24.400 209.600 ;
        RECT 25.200 208.300 26.000 209.200 ;
        RECT 30.000 208.300 30.800 208.400 ;
        RECT 25.200 207.700 30.800 208.300 ;
        RECT 25.200 207.600 26.000 207.700 ;
        RECT 30.000 207.600 30.800 207.700 ;
        RECT 23.800 206.400 27.400 207.000 ;
        RECT 23.800 206.200 24.400 206.400 ;
        RECT 23.600 202.200 24.400 206.200 ;
        RECT 26.800 202.200 27.600 206.400 ;
        RECT 31.800 206.200 32.400 210.400 ;
        RECT 35.000 210.200 35.600 211.600 ;
        RECT 40.000 211.000 40.600 214.400 ;
        RECT 41.400 212.400 42.000 215.800 ;
        RECT 44.000 214.200 44.800 219.800 ;
        RECT 52.400 218.400 53.200 219.800 ;
        RECT 55.600 218.400 56.400 219.800 ;
        RECT 52.400 217.800 53.400 218.400 ;
        RECT 52.800 217.600 53.400 217.800 ;
        RECT 55.600 217.600 58.000 218.400 ;
        RECT 52.800 217.000 56.800 217.600 ;
        RECT 50.800 215.600 52.600 216.400 ;
        RECT 41.200 211.600 42.000 212.400 ;
        RECT 31.600 202.200 32.400 206.200 ;
        RECT 34.800 202.200 35.600 210.200 ;
        RECT 38.200 210.400 40.600 211.000 ;
        RECT 38.200 206.200 38.800 210.400 ;
        RECT 41.400 210.200 42.000 211.600 ;
        RECT 43.000 213.800 44.800 214.200 ;
        RECT 43.000 213.600 44.600 213.800 ;
        RECT 52.400 213.600 54.000 214.400 ;
        RECT 43.000 210.400 43.600 213.600 ;
        RECT 45.200 211.600 46.800 212.400 ;
        RECT 54.000 211.600 55.600 212.400 ;
        RECT 38.000 202.200 38.800 206.200 ;
        RECT 41.200 202.200 42.000 210.200 ;
        RECT 42.800 209.600 43.600 210.400 ;
        RECT 47.600 209.600 48.400 211.200 ;
        RECT 56.200 210.400 56.800 217.000 ;
        RECT 65.600 214.200 66.400 219.800 ;
        RECT 72.000 214.200 72.800 219.800 ;
        RECT 78.400 216.300 79.200 219.800 ;
        RECT 82.800 217.800 83.600 219.800 ;
        RECT 81.200 216.300 82.000 217.200 ;
        RECT 78.400 215.700 82.000 216.300 ;
        RECT 78.400 214.200 79.200 215.700 ;
        RECT 81.200 215.600 82.000 215.700 ;
        RECT 83.000 215.600 83.600 217.800 ;
        RECT 86.000 215.800 86.800 219.800 ;
        RECT 88.200 216.400 89.000 219.800 ;
        RECT 88.200 215.800 90.000 216.400 ;
        RECT 83.000 215.000 85.400 215.600 ;
        RECT 65.600 213.800 67.400 214.200 ;
        RECT 72.000 213.800 73.800 214.200 ;
        RECT 78.400 213.800 80.200 214.200 ;
        RECT 65.800 213.600 67.400 213.800 ;
        RECT 72.200 213.600 73.800 213.800 ;
        RECT 78.600 213.600 80.200 213.800 ;
        RECT 82.800 213.600 83.800 214.400 ;
        RECT 63.600 211.600 65.200 212.400 ;
        RECT 56.200 209.800 59.600 210.400 ;
        RECT 58.800 209.600 59.600 209.800 ;
        RECT 62.000 209.600 62.800 211.200 ;
        RECT 66.800 210.400 67.400 213.600 ;
        RECT 70.000 211.600 71.600 212.400 ;
        RECT 66.800 209.600 67.600 210.400 ;
        RECT 68.400 209.600 69.200 211.200 ;
        RECT 73.200 210.400 73.800 213.600 ;
        RECT 76.400 211.600 78.000 212.400 ;
        RECT 73.200 209.600 74.000 210.400 ;
        RECT 74.800 209.600 75.600 211.200 ;
        RECT 79.600 210.400 80.200 213.600 ;
        RECT 83.200 212.800 84.000 213.600 ;
        RECT 84.800 212.000 85.400 215.000 ;
        RECT 86.200 212.400 86.800 215.800 ;
        RECT 84.600 211.400 85.400 212.000 ;
        RECT 86.000 211.600 86.800 212.400 ;
        RECT 81.200 211.200 85.400 211.400 ;
        RECT 81.200 210.800 85.200 211.200 ;
        RECT 79.600 209.600 80.400 210.400 ;
        RECT 43.000 207.000 43.600 209.600 ;
        RECT 44.400 207.600 45.200 209.200 ;
        RECT 49.400 208.800 53.000 209.400 ;
        RECT 49.400 208.200 50.000 208.800 ;
        RECT 43.000 206.400 46.600 207.000 ;
        RECT 43.000 206.200 43.600 206.400 ;
        RECT 42.800 202.200 43.600 206.200 ;
        RECT 46.000 206.200 46.600 206.400 ;
        RECT 46.000 202.200 46.800 206.200 ;
        RECT 49.200 202.200 50.000 208.200 ;
        RECT 52.400 208.200 53.000 208.800 ;
        RECT 54.200 209.000 57.800 209.200 ;
        RECT 58.800 209.000 59.400 209.600 ;
        RECT 54.200 208.600 58.000 209.000 ;
        RECT 54.200 208.200 54.800 208.600 ;
        RECT 52.400 202.800 53.200 208.200 ;
        RECT 54.000 203.400 54.800 208.200 ;
        RECT 55.600 202.800 56.400 208.000 ;
        RECT 57.200 203.000 58.000 208.600 ;
        RECT 58.800 203.400 59.600 209.000 ;
        RECT 52.400 202.200 56.400 202.800 ;
        RECT 57.400 202.800 58.000 203.000 ;
        RECT 60.400 203.000 61.200 209.000 ;
        RECT 65.200 207.600 66.000 209.200 ;
        RECT 66.800 207.000 67.400 209.600 ;
        RECT 71.600 207.600 72.400 209.200 ;
        RECT 73.200 207.000 73.800 209.600 ;
        RECT 78.000 207.600 78.800 209.200 ;
        RECT 79.600 207.000 80.200 209.600 ;
        RECT 63.800 206.400 67.400 207.000 ;
        RECT 63.800 206.200 64.400 206.400 ;
        RECT 60.400 202.800 61.000 203.000 ;
        RECT 57.400 202.200 61.000 202.800 ;
        RECT 63.600 202.200 64.400 206.200 ;
        RECT 66.800 206.200 67.400 206.400 ;
        RECT 70.200 206.400 73.800 207.000 ;
        RECT 70.200 206.200 70.800 206.400 ;
        RECT 66.800 202.200 67.600 206.200 ;
        RECT 70.000 202.200 70.800 206.200 ;
        RECT 73.200 206.200 73.800 206.400 ;
        RECT 76.600 206.400 80.200 207.000 ;
        RECT 76.600 206.200 77.200 206.400 ;
        RECT 73.200 202.200 74.000 206.200 ;
        RECT 76.400 202.200 77.200 206.200 ;
        RECT 79.600 206.200 80.200 206.400 ;
        RECT 79.600 202.200 80.400 206.200 ;
        RECT 81.200 202.200 82.000 210.800 ;
        RECT 86.200 210.200 86.800 211.600 ;
        RECT 85.400 209.600 86.800 210.200 ;
        RECT 85.400 202.200 86.200 209.600 ;
        RECT 87.600 208.800 88.400 210.400 ;
        RECT 89.200 202.200 90.000 215.800 ;
        RECT 95.600 215.800 96.400 219.800 ;
        RECT 97.000 216.400 97.800 217.200 ;
        RECT 101.400 216.400 102.200 219.800 ;
        RECT 90.800 214.300 91.600 215.200 ;
        RECT 94.000 214.300 94.800 214.400 ;
        RECT 90.800 213.700 94.800 214.300 ;
        RECT 90.800 213.600 91.600 213.700 ;
        RECT 94.000 212.800 94.800 213.700 ;
        RECT 92.400 212.200 93.200 212.400 ;
        RECT 95.600 212.200 96.200 215.800 ;
        RECT 97.200 215.600 98.000 216.400 ;
        RECT 100.400 215.800 102.200 216.400 ;
        RECT 103.600 216.000 104.400 219.800 ;
        RECT 106.800 216.000 107.600 219.800 ;
        RECT 103.600 215.800 107.600 216.000 ;
        RECT 108.400 218.300 109.200 219.800 ;
        RECT 113.200 218.300 114.000 218.400 ;
        RECT 108.400 217.700 114.000 218.300 ;
        RECT 108.400 215.800 109.200 217.700 ;
        RECT 113.200 217.600 114.000 217.700 ;
        RECT 97.200 214.300 98.000 214.400 ;
        RECT 98.800 214.300 99.600 215.200 ;
        RECT 97.200 213.700 99.600 214.300 ;
        RECT 97.200 213.600 98.000 213.700 ;
        RECT 98.800 213.600 99.600 213.700 ;
        RECT 97.200 212.200 98.000 212.400 ;
        RECT 92.400 211.600 94.000 212.200 ;
        RECT 95.600 211.600 98.000 212.200 ;
        RECT 93.200 211.200 94.000 211.600 ;
        RECT 97.200 210.200 97.800 211.600 ;
        RECT 92.400 209.600 96.400 210.200 ;
        RECT 92.400 202.200 93.200 209.600 ;
        RECT 95.600 202.200 96.400 209.600 ;
        RECT 97.200 202.200 98.000 210.200 ;
        RECT 100.400 202.200 101.200 215.800 ;
        RECT 103.800 215.400 107.400 215.800 ;
        RECT 104.400 214.400 105.200 214.800 ;
        RECT 108.400 214.400 109.000 215.800 ;
        RECT 103.600 213.800 105.200 214.400 ;
        RECT 103.600 213.600 104.400 213.800 ;
        RECT 106.600 213.600 109.200 214.400 ;
        RECT 116.400 213.800 117.200 219.800 ;
        RECT 122.800 216.600 123.600 219.800 ;
        RECT 124.400 217.000 125.200 219.800 ;
        RECT 126.000 217.000 126.800 219.800 ;
        RECT 127.600 217.000 128.400 219.800 ;
        RECT 130.800 217.000 131.600 219.800 ;
        RECT 134.000 217.000 134.800 219.800 ;
        RECT 135.600 217.000 136.400 219.800 ;
        RECT 137.200 217.000 138.000 219.800 ;
        RECT 138.800 217.000 139.600 219.800 ;
        RECT 121.000 215.800 123.600 216.600 ;
        RECT 140.400 216.600 141.200 219.800 ;
        RECT 127.000 215.800 131.600 216.400 ;
        RECT 121.000 215.200 121.800 215.800 ;
        RECT 118.800 214.400 121.800 215.200 ;
        RECT 105.200 211.600 106.000 213.200 ;
        RECT 102.000 208.800 102.800 210.400 ;
        RECT 106.600 210.200 107.200 213.600 ;
        RECT 116.400 213.000 125.200 213.800 ;
        RECT 127.000 213.400 127.800 215.800 ;
        RECT 130.800 215.600 131.600 215.800 ;
        RECT 132.400 215.600 134.000 216.400 ;
        RECT 137.000 215.600 138.000 216.400 ;
        RECT 140.400 215.800 142.800 216.600 ;
        RECT 129.200 213.600 130.000 215.200 ;
        RECT 130.800 214.800 131.600 215.000 ;
        RECT 130.800 214.200 135.200 214.800 ;
        RECT 134.400 214.000 135.200 214.200 ;
        RECT 108.400 210.200 109.200 210.400 ;
        RECT 106.200 209.600 107.200 210.200 ;
        RECT 107.800 209.600 109.200 210.200 ;
        RECT 106.200 202.200 107.000 209.600 ;
        RECT 107.800 208.400 108.400 209.600 ;
        RECT 107.600 207.600 108.400 208.400 ;
        RECT 116.400 207.400 117.200 213.000 ;
        RECT 125.800 212.600 127.800 213.400 ;
        RECT 131.600 212.600 134.800 213.400 ;
        RECT 137.200 212.800 138.000 215.600 ;
        RECT 142.000 215.200 142.800 215.800 ;
        RECT 142.000 214.600 143.800 215.200 ;
        RECT 143.000 213.400 143.800 214.600 ;
        RECT 146.800 214.600 147.600 219.800 ;
        RECT 148.400 216.000 149.200 219.800 ;
        RECT 153.200 217.800 154.000 219.800 ;
        RECT 151.600 216.300 152.400 216.400 ;
        RECT 153.200 216.300 153.800 217.800 ;
        RECT 148.400 215.200 149.400 216.000 ;
        RECT 151.600 215.700 153.900 216.300 ;
        RECT 151.600 215.600 152.400 215.700 ;
        RECT 146.800 214.000 148.000 214.600 ;
        RECT 143.000 212.600 146.800 213.400 ;
        RECT 117.800 212.000 118.600 212.200 ;
        RECT 122.800 212.000 123.600 212.400 ;
        RECT 129.200 212.000 130.000 212.400 ;
        RECT 140.400 212.000 141.200 212.600 ;
        RECT 147.400 212.000 148.000 214.000 ;
        RECT 117.800 211.400 141.200 212.000 ;
        RECT 147.200 211.400 148.000 212.000 ;
        RECT 148.600 212.300 149.400 215.200 ;
        RECT 153.200 214.400 153.800 215.700 ;
        RECT 154.800 215.600 155.600 217.200 ;
        RECT 159.000 216.400 159.800 219.800 ;
        RECT 158.000 215.800 159.800 216.400 ;
        RECT 161.200 216.000 162.000 219.800 ;
        RECT 164.400 216.000 165.200 219.800 ;
        RECT 161.200 215.800 165.200 216.000 ;
        RECT 166.000 215.800 166.800 219.800 ;
        RECT 170.200 216.400 171.800 219.800 ;
        RECT 169.200 215.800 171.800 216.400 ;
        RECT 153.200 213.600 154.000 214.400 ;
        RECT 156.400 213.600 157.200 215.200 ;
        RECT 151.600 212.300 152.400 212.400 ;
        RECT 148.600 211.700 152.400 212.300 ;
        RECT 147.200 209.600 147.800 211.400 ;
        RECT 148.600 210.800 149.400 211.700 ;
        RECT 151.600 210.800 152.400 211.700 ;
        RECT 126.000 209.400 126.800 209.600 ;
        RECT 121.400 209.000 126.800 209.400 ;
        RECT 120.600 208.800 126.800 209.000 ;
        RECT 127.800 209.000 136.400 209.600 ;
        RECT 118.000 208.000 119.600 208.800 ;
        RECT 120.600 208.200 122.000 208.800 ;
        RECT 127.800 208.200 128.400 209.000 ;
        RECT 135.600 208.800 136.400 209.000 ;
        RECT 138.800 209.000 147.800 209.600 ;
        RECT 138.800 208.800 139.600 209.000 ;
        RECT 119.000 207.600 119.600 208.000 ;
        RECT 122.600 207.600 128.400 208.200 ;
        RECT 129.000 207.600 131.600 208.400 ;
        RECT 116.400 206.800 118.400 207.400 ;
        RECT 119.000 206.800 123.200 207.600 ;
        RECT 117.800 206.200 118.400 206.800 ;
        RECT 117.800 205.600 118.800 206.200 ;
        RECT 118.000 202.200 118.800 205.600 ;
        RECT 121.200 202.200 122.000 206.800 ;
        RECT 124.400 202.200 125.200 205.000 ;
        RECT 126.000 202.200 126.800 205.000 ;
        RECT 127.600 202.200 128.400 207.000 ;
        RECT 130.800 202.200 131.600 207.000 ;
        RECT 134.000 202.200 134.800 208.400 ;
        RECT 142.000 207.600 144.600 208.400 ;
        RECT 137.200 206.800 141.400 207.600 ;
        RECT 135.600 202.200 136.400 205.000 ;
        RECT 137.200 202.200 138.000 205.000 ;
        RECT 138.800 202.200 139.600 205.000 ;
        RECT 142.000 202.200 142.800 207.600 ;
        RECT 147.200 207.400 147.800 209.000 ;
        RECT 145.200 206.800 147.800 207.400 ;
        RECT 148.400 210.000 149.400 210.800 ;
        RECT 153.200 210.200 153.800 213.600 ;
        RECT 145.200 202.200 146.000 206.800 ;
        RECT 148.400 202.200 149.200 210.000 ;
        RECT 152.200 209.400 154.000 210.200 ;
        RECT 152.200 202.200 153.000 209.400 ;
        RECT 158.000 202.200 158.800 215.800 ;
        RECT 161.400 215.400 165.000 215.800 ;
        RECT 162.000 214.400 162.800 214.800 ;
        RECT 166.000 214.400 166.600 215.800 ;
        RECT 169.200 215.600 171.400 215.800 ;
        RECT 161.200 213.800 162.800 214.400 ;
        RECT 161.200 213.600 162.000 213.800 ;
        RECT 164.200 213.600 166.800 214.400 ;
        RECT 167.600 214.300 168.400 214.400 ;
        RECT 169.200 214.300 170.000 214.400 ;
        RECT 167.600 213.700 170.000 214.300 ;
        RECT 167.600 213.600 168.400 213.700 ;
        RECT 169.200 213.600 170.000 213.700 ;
        RECT 162.800 211.600 163.600 213.200 ;
        RECT 159.600 208.800 160.400 210.400 ;
        RECT 164.200 210.200 164.800 213.600 ;
        RECT 169.400 213.200 170.000 213.600 ;
        RECT 169.400 212.400 170.200 213.200 ;
        RECT 170.800 212.400 171.400 215.600 ;
        RECT 172.400 214.300 173.200 214.400 ;
        RECT 174.000 214.300 174.800 214.400 ;
        RECT 172.400 213.700 174.800 214.300 ;
        RECT 172.400 212.800 173.200 213.700 ;
        RECT 174.000 213.600 174.800 213.700 ;
        RECT 167.600 212.300 168.400 212.400 ;
        RECT 166.100 211.700 168.400 212.300 ;
        RECT 166.100 210.400 166.700 211.700 ;
        RECT 167.600 210.800 168.400 211.700 ;
        RECT 170.800 211.600 171.600 212.400 ;
        RECT 174.000 212.200 174.800 212.400 ;
        RECT 173.200 211.600 174.800 212.200 ;
        RECT 170.800 211.400 171.400 211.600 ;
        RECT 169.400 210.800 171.400 211.400 ;
        RECT 173.200 211.200 174.000 211.600 ;
        RECT 166.000 210.200 166.800 210.400 ;
        RECT 169.400 210.200 170.000 210.800 ;
        RECT 163.800 209.600 164.800 210.200 ;
        RECT 165.400 209.600 166.800 210.200 ;
        RECT 163.800 202.200 164.600 209.600 ;
        RECT 165.400 208.400 166.000 209.600 ;
        RECT 165.200 207.600 166.000 208.400 ;
        RECT 167.600 202.800 168.400 210.200 ;
        RECT 169.200 203.400 170.000 210.200 ;
        RECT 170.800 209.600 174.800 210.200 ;
        RECT 170.800 202.800 171.600 209.600 ;
        RECT 167.600 202.200 171.600 202.800 ;
        RECT 174.000 202.200 174.800 209.600 ;
        RECT 175.600 202.200 176.400 219.800 ;
        RECT 177.200 215.600 178.000 217.200 ;
        RECT 178.800 215.800 179.600 219.800 ;
        RECT 183.000 216.800 183.800 219.800 ;
        RECT 186.800 217.800 187.600 219.800 ;
        RECT 183.000 215.800 184.400 216.800 ;
        RECT 179.000 215.600 179.600 215.800 ;
        RECT 179.000 215.200 180.800 215.600 ;
        RECT 179.000 215.000 183.200 215.200 ;
        RECT 180.200 214.600 183.200 215.000 ;
        RECT 182.400 214.400 183.200 214.600 ;
        RECT 178.800 212.800 179.600 214.400 ;
        RECT 180.800 213.800 181.600 214.000 ;
        RECT 180.600 213.200 181.600 213.800 ;
        RECT 180.600 212.400 181.200 213.200 ;
        RECT 180.400 211.600 181.200 212.400 ;
        RECT 182.400 211.000 183.000 214.400 ;
        RECT 183.800 212.400 184.400 215.800 ;
        RECT 186.800 214.400 187.400 217.800 ;
        RECT 188.400 215.600 189.200 217.200 ;
        RECT 190.000 216.000 190.800 219.800 ;
        RECT 193.200 216.000 194.000 219.800 ;
        RECT 190.000 215.800 194.000 216.000 ;
        RECT 194.800 215.800 195.600 219.800 ;
        RECT 199.000 216.400 199.800 219.800 ;
        RECT 198.000 215.800 199.800 216.400 ;
        RECT 190.200 215.400 193.800 215.800 ;
        RECT 190.800 214.400 191.600 214.800 ;
        RECT 194.800 214.400 195.400 215.800 ;
        RECT 186.800 214.300 187.600 214.400 ;
        RECT 190.000 214.300 191.600 214.400 ;
        RECT 186.800 213.800 191.600 214.300 ;
        RECT 186.800 213.700 190.800 213.800 ;
        RECT 186.800 213.600 187.600 213.700 ;
        RECT 190.000 213.600 190.800 213.700 ;
        RECT 193.000 213.600 195.600 214.400 ;
        RECT 196.400 213.600 197.200 215.200 ;
        RECT 183.600 211.600 184.400 212.400 ;
        RECT 180.600 210.400 183.000 211.000 ;
        RECT 180.600 206.200 181.200 210.400 ;
        RECT 183.800 210.200 184.400 211.600 ;
        RECT 185.200 210.800 186.000 212.400 ;
        RECT 186.800 210.200 187.400 213.600 ;
        RECT 191.600 211.600 192.400 213.200 ;
        RECT 193.000 210.200 193.600 213.600 ;
        RECT 194.800 210.200 195.600 210.400 ;
        RECT 180.400 202.200 181.200 206.200 ;
        RECT 183.600 202.200 184.400 210.200 ;
        RECT 185.800 209.400 187.600 210.200 ;
        RECT 192.600 209.600 193.600 210.200 ;
        RECT 194.200 209.600 195.600 210.200 ;
        RECT 185.800 202.200 186.600 209.400 ;
        RECT 192.600 208.400 193.400 209.600 ;
        RECT 194.200 208.400 194.800 209.600 ;
        RECT 191.600 207.600 193.400 208.400 ;
        RECT 194.000 207.600 194.800 208.400 ;
        RECT 192.600 202.200 193.400 207.600 ;
        RECT 198.000 202.200 198.800 215.800 ;
        RECT 202.400 214.200 203.200 219.800 ;
        RECT 210.200 218.400 211.800 219.800 ;
        RECT 209.200 217.600 211.800 218.400 ;
        RECT 210.200 215.800 211.800 217.600 ;
        RECT 216.200 216.400 217.000 219.800 ;
        RECT 216.200 215.800 218.000 216.400 ;
        RECT 220.400 216.000 221.200 219.800 ;
        RECT 223.600 216.000 224.400 219.800 ;
        RECT 220.400 215.800 224.400 216.000 ;
        RECT 225.200 215.800 226.000 219.800 ;
        RECT 226.800 216.000 227.600 219.800 ;
        RECT 230.000 216.000 230.800 219.800 ;
        RECT 226.800 215.800 230.800 216.000 ;
        RECT 231.600 215.800 232.400 219.800 ;
        RECT 236.400 215.800 237.200 219.800 ;
        RECT 237.800 216.400 238.600 217.200 ;
        RECT 238.000 216.300 238.800 216.400 ;
        RECT 239.600 216.300 240.400 219.800 ;
        RECT 201.400 213.800 203.200 214.200 ;
        RECT 201.400 213.600 203.000 213.800 ;
        RECT 209.200 213.600 210.000 214.400 ;
        RECT 201.400 210.400 202.000 213.600 ;
        RECT 209.400 213.200 210.000 213.600 ;
        RECT 209.400 212.400 210.200 213.200 ;
        RECT 210.800 212.400 211.400 215.800 ;
        RECT 212.400 214.300 213.200 214.400 ;
        RECT 215.600 214.300 216.400 214.400 ;
        RECT 212.400 213.700 216.400 214.300 ;
        RECT 212.400 212.800 213.200 213.700 ;
        RECT 215.600 213.600 216.400 213.700 ;
        RECT 203.600 211.600 205.200 212.400 ;
        RECT 199.600 208.800 200.400 210.400 ;
        RECT 201.200 209.600 202.000 210.400 ;
        RECT 206.000 209.600 206.800 211.200 ;
        RECT 207.600 210.800 208.400 212.400 ;
        RECT 210.800 211.600 211.600 212.400 ;
        RECT 214.000 212.200 214.800 212.400 ;
        RECT 213.200 211.600 214.800 212.200 ;
        RECT 210.800 211.400 211.400 211.600 ;
        RECT 209.400 210.800 211.400 211.400 ;
        RECT 213.200 211.200 214.000 211.600 ;
        RECT 209.400 210.200 210.000 210.800 ;
        RECT 201.400 207.000 202.000 209.600 ;
        RECT 202.800 207.600 203.600 209.200 ;
        RECT 201.400 206.400 205.000 207.000 ;
        RECT 201.400 206.200 202.000 206.400 ;
        RECT 201.200 202.200 202.000 206.200 ;
        RECT 204.400 206.200 205.000 206.400 ;
        RECT 204.400 202.200 205.200 206.200 ;
        RECT 207.600 202.800 208.400 210.200 ;
        RECT 209.200 203.400 210.000 210.200 ;
        RECT 210.800 209.600 214.800 210.200 ;
        RECT 210.800 202.800 211.600 209.600 ;
        RECT 207.600 202.200 211.600 202.800 ;
        RECT 214.000 202.200 214.800 209.600 ;
        RECT 215.600 208.800 216.400 210.400 ;
        RECT 217.200 202.200 218.000 215.800 ;
        RECT 220.600 215.400 224.200 215.800 ;
        RECT 218.800 213.600 219.600 215.200 ;
        RECT 221.200 214.400 222.000 214.800 ;
        RECT 225.200 214.400 225.800 215.800 ;
        RECT 227.000 215.400 230.600 215.800 ;
        RECT 227.600 214.400 228.400 214.800 ;
        RECT 231.600 214.400 232.200 215.800 ;
        RECT 220.400 213.800 222.000 214.400 ;
        RECT 220.400 213.600 221.200 213.800 ;
        RECT 223.400 213.600 226.000 214.400 ;
        RECT 226.800 213.800 228.400 214.400 ;
        RECT 229.800 214.300 232.400 214.400 ;
        RECT 234.800 214.300 235.600 214.400 ;
        RECT 226.800 213.600 227.600 213.800 ;
        RECT 229.800 213.700 235.600 214.300 ;
        RECT 229.800 213.600 232.400 213.700 ;
        RECT 222.000 211.600 222.800 213.200 ;
        RECT 223.400 212.300 224.000 213.600 ;
        RECT 226.800 212.300 227.600 212.400 ;
        RECT 223.400 211.700 227.600 212.300 ;
        RECT 223.400 210.200 224.000 211.700 ;
        RECT 226.800 211.600 227.600 211.700 ;
        RECT 228.400 211.600 229.200 213.200 ;
        RECT 225.200 210.200 226.000 210.400 ;
        RECT 229.800 210.200 230.400 213.600 ;
        RECT 234.800 212.800 235.600 213.700 ;
        RECT 233.200 212.200 234.000 212.400 ;
        RECT 236.400 212.200 237.000 215.800 ;
        RECT 238.000 215.700 240.400 216.300 ;
        RECT 241.200 216.000 242.000 219.800 ;
        RECT 244.400 216.000 245.200 219.800 ;
        RECT 247.600 216.000 248.400 219.800 ;
        RECT 241.200 215.800 245.200 216.000 ;
        RECT 238.000 215.600 238.800 215.700 ;
        RECT 239.800 214.400 240.400 215.700 ;
        RECT 241.400 215.400 245.000 215.800 ;
        RECT 247.400 215.200 248.400 216.000 ;
        RECT 243.600 214.400 244.400 214.800 ;
        RECT 239.600 213.600 242.200 214.400 ;
        RECT 243.600 213.800 245.200 214.400 ;
        RECT 244.400 213.600 245.200 213.800 ;
        RECT 238.000 212.300 238.800 212.400 ;
        RECT 239.600 212.300 240.400 212.400 ;
        RECT 238.000 212.200 240.400 212.300 ;
        RECT 233.200 211.600 234.800 212.200 ;
        RECT 236.400 211.700 240.400 212.200 ;
        RECT 236.400 211.600 238.800 211.700 ;
        RECT 239.600 211.600 240.400 211.700 ;
        RECT 234.000 211.200 234.800 211.600 ;
        RECT 231.600 210.200 232.400 210.400 ;
        RECT 238.000 210.200 238.600 211.600 ;
        RECT 239.600 210.200 240.400 210.400 ;
        RECT 241.600 210.200 242.200 213.600 ;
        RECT 242.800 212.300 243.600 213.200 ;
        RECT 246.000 212.300 246.800 212.400 ;
        RECT 242.800 211.700 246.800 212.300 ;
        RECT 242.800 211.600 243.600 211.700 ;
        RECT 246.000 211.600 246.800 211.700 ;
        RECT 247.400 210.800 248.200 215.200 ;
        RECT 249.200 214.600 250.000 219.800 ;
        RECT 255.600 216.600 256.400 219.800 ;
        RECT 257.200 217.000 258.000 219.800 ;
        RECT 258.800 217.000 259.600 219.800 ;
        RECT 260.400 217.000 261.200 219.800 ;
        RECT 262.000 217.000 262.800 219.800 ;
        RECT 265.200 217.000 266.000 219.800 ;
        RECT 268.400 217.000 269.200 219.800 ;
        RECT 270.000 217.000 270.800 219.800 ;
        RECT 271.600 217.000 272.400 219.800 ;
        RECT 254.000 215.800 256.400 216.600 ;
        RECT 273.200 216.600 274.000 219.800 ;
        RECT 254.000 215.200 254.800 215.800 ;
        RECT 248.800 214.000 250.000 214.600 ;
        RECT 253.000 214.600 254.800 215.200 ;
        RECT 258.800 215.600 259.800 216.400 ;
        RECT 262.800 215.600 264.400 216.400 ;
        RECT 265.200 215.800 269.800 216.400 ;
        RECT 273.200 215.800 275.800 216.600 ;
        RECT 265.200 215.600 266.000 215.800 ;
        RECT 248.800 212.000 249.400 214.000 ;
        RECT 253.000 213.400 253.800 214.600 ;
        RECT 250.000 212.600 253.800 213.400 ;
        RECT 258.800 212.800 259.600 215.600 ;
        RECT 265.200 214.800 266.000 215.000 ;
        RECT 261.600 214.200 266.000 214.800 ;
        RECT 261.600 214.000 262.400 214.200 ;
        RECT 266.800 213.600 267.600 215.200 ;
        RECT 269.000 213.400 269.800 215.800 ;
        RECT 275.000 215.200 275.800 215.800 ;
        RECT 275.000 214.400 278.000 215.200 ;
        RECT 279.600 213.800 280.400 219.800 ;
        RECT 286.000 216.300 286.800 216.400 ;
        RECT 287.600 216.300 288.400 217.200 ;
        RECT 286.000 215.700 288.400 216.300 ;
        RECT 286.000 215.600 286.800 215.700 ;
        RECT 287.600 215.600 288.400 215.700 ;
        RECT 262.000 212.600 265.200 213.400 ;
        RECT 269.000 212.600 271.000 213.400 ;
        RECT 271.600 213.000 280.400 213.800 ;
        RECT 255.600 212.000 256.400 212.600 ;
        RECT 273.200 212.000 274.000 212.400 ;
        RECT 276.400 212.000 277.200 212.400 ;
        RECT 278.200 212.000 279.000 212.200 ;
        RECT 248.800 211.400 249.600 212.000 ;
        RECT 255.600 211.400 279.000 212.000 ;
        RECT 223.000 209.600 224.000 210.200 ;
        RECT 224.600 209.600 226.000 210.200 ;
        RECT 229.400 209.600 230.400 210.200 ;
        RECT 231.000 209.600 232.400 210.200 ;
        RECT 233.200 209.600 237.200 210.200 ;
        RECT 223.000 202.200 223.800 209.600 ;
        RECT 224.600 208.400 225.200 209.600 ;
        RECT 224.400 207.600 225.200 208.400 ;
        RECT 229.400 202.200 230.200 209.600 ;
        RECT 231.000 208.400 231.600 209.600 ;
        RECT 230.800 207.600 231.600 208.400 ;
        RECT 233.200 202.200 234.000 209.600 ;
        RECT 236.400 202.200 237.200 209.600 ;
        RECT 238.000 202.200 238.800 210.200 ;
        RECT 239.600 209.600 241.000 210.200 ;
        RECT 241.600 209.600 242.600 210.200 ;
        RECT 247.400 210.000 248.400 210.800 ;
        RECT 240.400 208.400 241.000 209.600 ;
        RECT 240.400 207.600 241.200 208.400 ;
        RECT 241.800 202.200 242.600 209.600 ;
        RECT 247.600 202.200 248.400 210.000 ;
        RECT 249.000 209.600 249.600 211.400 ;
        RECT 249.000 209.000 258.000 209.600 ;
        RECT 249.000 207.400 249.600 209.000 ;
        RECT 257.200 208.800 258.000 209.000 ;
        RECT 260.400 209.000 269.000 209.600 ;
        RECT 260.400 208.800 261.200 209.000 ;
        RECT 252.200 207.600 254.800 208.400 ;
        RECT 249.000 206.800 251.600 207.400 ;
        RECT 250.800 202.200 251.600 206.800 ;
        RECT 254.000 202.200 254.800 207.600 ;
        RECT 255.400 206.800 259.600 207.600 ;
        RECT 257.200 202.200 258.000 205.000 ;
        RECT 258.800 202.200 259.600 205.000 ;
        RECT 260.400 202.200 261.200 205.000 ;
        RECT 262.000 202.200 262.800 208.400 ;
        RECT 265.200 207.600 267.800 208.400 ;
        RECT 268.400 208.200 269.000 209.000 ;
        RECT 270.000 209.400 270.800 209.600 ;
        RECT 270.000 209.000 275.400 209.400 ;
        RECT 270.000 208.800 276.200 209.000 ;
        RECT 274.800 208.200 276.200 208.800 ;
        RECT 268.400 207.600 274.200 208.200 ;
        RECT 277.200 208.000 278.800 208.800 ;
        RECT 277.200 207.600 277.800 208.000 ;
        RECT 265.200 202.200 266.000 207.000 ;
        RECT 268.400 202.200 269.200 207.000 ;
        RECT 273.600 206.800 277.800 207.600 ;
        RECT 279.600 207.400 280.400 213.000 ;
        RECT 278.400 206.800 280.400 207.400 ;
        RECT 270.000 202.200 270.800 205.000 ;
        RECT 271.600 202.200 272.400 205.000 ;
        RECT 274.800 202.200 275.600 206.800 ;
        RECT 278.400 206.200 279.000 206.800 ;
        RECT 278.000 205.600 279.000 206.200 ;
        RECT 278.000 202.200 278.800 205.600 ;
        RECT 289.200 202.200 290.000 219.800 ;
        RECT 292.400 216.000 293.200 219.800 ;
        RECT 292.200 215.200 293.200 216.000 ;
        RECT 292.200 210.800 293.000 215.200 ;
        RECT 294.000 214.600 294.800 219.800 ;
        RECT 300.400 216.600 301.200 219.800 ;
        RECT 302.000 217.000 302.800 219.800 ;
        RECT 303.600 217.000 304.400 219.800 ;
        RECT 305.200 217.000 306.000 219.800 ;
        RECT 306.800 217.000 307.600 219.800 ;
        RECT 310.000 217.000 310.800 219.800 ;
        RECT 313.200 217.000 314.000 219.800 ;
        RECT 314.800 217.000 315.600 219.800 ;
        RECT 316.400 217.000 317.200 219.800 ;
        RECT 298.800 215.800 301.200 216.600 ;
        RECT 318.000 216.600 318.800 219.800 ;
        RECT 298.800 215.200 299.600 215.800 ;
        RECT 293.600 214.000 294.800 214.600 ;
        RECT 297.800 214.600 299.600 215.200 ;
        RECT 303.600 215.600 304.600 216.400 ;
        RECT 307.600 215.600 309.200 216.400 ;
        RECT 310.000 215.800 314.600 216.400 ;
        RECT 318.000 215.800 320.600 216.600 ;
        RECT 310.000 215.600 310.800 215.800 ;
        RECT 293.600 212.000 294.200 214.000 ;
        RECT 297.800 213.400 298.600 214.600 ;
        RECT 294.800 212.600 298.600 213.400 ;
        RECT 303.600 212.800 304.400 215.600 ;
        RECT 310.000 214.800 310.800 215.000 ;
        RECT 306.400 214.200 310.800 214.800 ;
        RECT 306.400 214.000 307.200 214.200 ;
        RECT 311.600 213.600 312.400 215.200 ;
        RECT 313.800 213.400 314.600 215.800 ;
        RECT 319.800 215.200 320.600 215.800 ;
        RECT 319.800 214.400 322.800 215.200 ;
        RECT 324.400 213.800 325.200 219.800 ;
        RECT 326.000 215.600 326.800 217.200 ;
        RECT 306.800 212.600 310.000 213.400 ;
        RECT 313.800 212.600 315.800 213.400 ;
        RECT 316.400 213.000 325.200 213.800 ;
        RECT 293.600 211.400 294.400 212.000 ;
        RECT 292.200 210.000 293.200 210.800 ;
        RECT 292.400 202.200 293.200 210.000 ;
        RECT 293.800 209.600 294.400 211.400 ;
        RECT 295.000 210.800 295.800 211.000 ;
        RECT 295.000 210.200 322.000 210.800 ;
        RECT 317.800 210.000 318.800 210.200 ;
        RECT 321.200 209.600 322.000 210.200 ;
        RECT 293.800 209.000 302.800 209.600 ;
        RECT 293.800 207.400 294.400 209.000 ;
        RECT 302.000 208.800 302.800 209.000 ;
        RECT 305.200 209.000 313.800 209.600 ;
        RECT 305.200 208.800 306.000 209.000 ;
        RECT 297.000 207.600 299.600 208.400 ;
        RECT 293.800 206.800 296.400 207.400 ;
        RECT 295.600 202.200 296.400 206.800 ;
        RECT 298.800 202.200 299.600 207.600 ;
        RECT 300.200 206.800 304.400 207.600 ;
        RECT 302.000 202.200 302.800 205.000 ;
        RECT 303.600 202.200 304.400 205.000 ;
        RECT 305.200 202.200 306.000 205.000 ;
        RECT 306.800 202.200 307.600 208.400 ;
        RECT 310.000 207.600 312.600 208.400 ;
        RECT 313.200 208.200 313.800 209.000 ;
        RECT 314.800 209.400 315.600 209.600 ;
        RECT 314.800 209.000 320.200 209.400 ;
        RECT 314.800 208.800 321.000 209.000 ;
        RECT 319.600 208.200 321.000 208.800 ;
        RECT 313.200 207.600 319.000 208.200 ;
        RECT 322.000 208.000 323.600 208.800 ;
        RECT 322.000 207.600 322.600 208.000 ;
        RECT 310.000 202.200 310.800 207.000 ;
        RECT 313.200 202.200 314.000 207.000 ;
        RECT 318.400 206.800 322.600 207.600 ;
        RECT 324.400 207.400 325.200 213.000 ;
        RECT 323.200 206.800 325.200 207.400 ;
        RECT 327.600 214.300 328.400 219.800 ;
        RECT 329.200 216.000 330.000 219.800 ;
        RECT 332.400 216.000 333.200 219.800 ;
        RECT 329.200 215.800 333.200 216.000 ;
        RECT 334.000 215.800 334.800 219.800 ;
        RECT 335.600 215.800 336.400 219.800 ;
        RECT 337.200 216.000 338.000 219.800 ;
        RECT 340.400 216.000 341.200 219.800 ;
        RECT 337.200 215.800 341.200 216.000 ;
        RECT 329.400 215.400 333.000 215.800 ;
        RECT 330.000 214.400 330.800 214.800 ;
        RECT 334.000 214.400 334.600 215.800 ;
        RECT 335.800 214.400 336.400 215.800 ;
        RECT 337.400 215.400 341.000 215.800 ;
        RECT 342.000 215.600 342.800 217.200 ;
        RECT 339.600 214.400 340.400 214.800 ;
        RECT 329.200 214.300 330.800 214.400 ;
        RECT 327.600 213.800 330.800 214.300 ;
        RECT 327.600 213.700 330.000 213.800 ;
        RECT 314.800 202.200 315.600 205.000 ;
        RECT 316.400 202.200 317.200 205.000 ;
        RECT 319.600 202.200 320.400 206.800 ;
        RECT 323.200 206.200 323.800 206.800 ;
        RECT 322.800 205.600 323.800 206.200 ;
        RECT 322.800 202.200 323.600 205.600 ;
        RECT 327.600 202.200 328.400 213.700 ;
        RECT 329.200 213.600 330.000 213.700 ;
        RECT 332.200 213.600 334.800 214.400 ;
        RECT 335.600 213.600 338.200 214.400 ;
        RECT 339.600 214.300 341.200 214.400 ;
        RECT 342.000 214.300 342.800 214.400 ;
        RECT 339.600 213.800 342.800 214.300 ;
        RECT 340.400 213.700 342.800 213.800 ;
        RECT 340.400 213.600 341.200 213.700 ;
        RECT 342.000 213.600 342.800 213.700 ;
        RECT 330.800 211.600 331.600 213.200 ;
        RECT 332.200 210.200 332.800 213.600 ;
        RECT 337.600 212.300 338.200 213.600 ;
        RECT 334.100 211.700 338.200 212.300 ;
        RECT 334.100 210.400 334.700 211.700 ;
        RECT 334.000 210.200 334.800 210.400 ;
        RECT 331.800 209.600 332.800 210.200 ;
        RECT 333.400 209.600 334.800 210.200 ;
        RECT 335.600 210.200 336.400 210.400 ;
        RECT 337.600 210.200 338.200 211.700 ;
        RECT 335.600 209.600 337.000 210.200 ;
        RECT 337.600 209.600 338.600 210.200 ;
        RECT 331.800 202.200 332.600 209.600 ;
        RECT 333.400 208.400 334.000 209.600 ;
        RECT 333.200 207.600 334.000 208.400 ;
        RECT 336.400 208.400 337.000 209.600 ;
        RECT 336.400 207.600 337.200 208.400 ;
        RECT 337.800 202.200 338.600 209.600 ;
        RECT 343.600 202.200 344.400 219.800 ;
        RECT 345.200 215.400 346.000 219.800 ;
        RECT 349.400 218.400 350.600 219.800 ;
        RECT 349.400 217.800 350.800 218.400 ;
        RECT 354.000 217.800 354.800 219.800 ;
        RECT 358.400 218.400 359.200 219.800 ;
        RECT 358.400 217.800 360.400 218.400 ;
        RECT 350.000 217.000 350.800 217.800 ;
        RECT 354.200 217.200 354.800 217.800 ;
        RECT 354.200 216.600 357.000 217.200 ;
        RECT 356.200 216.400 357.000 216.600 ;
        RECT 358.000 216.400 358.800 217.200 ;
        RECT 359.600 217.000 360.400 217.800 ;
        RECT 348.200 215.400 349.000 215.600 ;
        RECT 345.200 214.800 349.000 215.400 ;
        RECT 345.200 211.400 346.000 214.800 ;
        RECT 352.200 214.200 353.000 214.400 ;
        RECT 358.000 214.200 358.600 216.400 ;
        RECT 362.800 215.000 363.600 219.800 ;
        RECT 364.400 215.800 365.200 219.800 ;
        RECT 366.000 216.000 366.800 219.800 ;
        RECT 369.200 216.000 370.000 219.800 ;
        RECT 366.000 215.800 370.000 216.000 ;
        RECT 370.800 219.200 374.800 219.800 ;
        RECT 370.800 215.800 371.600 219.200 ;
        RECT 372.400 215.800 373.200 218.600 ;
        RECT 374.000 216.000 374.800 219.200 ;
        RECT 377.200 216.000 378.000 219.800 ;
        RECT 379.000 216.400 379.800 217.200 ;
        RECT 374.000 215.800 378.000 216.000 ;
        RECT 364.600 214.400 365.200 215.800 ;
        RECT 366.200 215.400 369.800 215.800 ;
        RECT 368.400 214.400 369.200 214.800 ;
        RECT 372.400 214.400 373.000 215.800 ;
        RECT 374.200 215.400 377.800 215.800 ;
        RECT 378.800 215.600 379.600 216.400 ;
        RECT 380.400 215.800 381.200 219.800 ;
        RECT 387.800 218.400 388.600 219.800 ;
        RECT 387.800 217.600 389.200 218.400 ;
        RECT 387.800 216.400 388.600 217.600 ;
        RECT 376.400 214.400 377.200 214.800 ;
        RECT 380.600 214.400 381.200 215.800 ;
        RECT 386.800 215.800 388.600 216.400 ;
        RECT 390.000 216.000 390.800 219.800 ;
        RECT 393.200 216.000 394.000 219.800 ;
        RECT 390.000 215.800 394.000 216.000 ;
        RECT 394.800 215.800 395.600 219.800 ;
        RECT 396.400 219.200 400.400 219.800 ;
        RECT 396.400 215.800 397.200 219.200 ;
        RECT 398.000 215.800 398.800 218.600 ;
        RECT 399.600 216.000 400.400 219.200 ;
        RECT 402.800 216.000 403.600 219.800 ;
        RECT 399.600 215.800 403.600 216.000 ;
        RECT 404.400 219.200 408.400 219.800 ;
        RECT 404.400 215.800 405.200 219.200 ;
        RECT 406.000 215.800 406.800 218.600 ;
        RECT 407.600 216.000 408.400 219.200 ;
        RECT 410.800 216.000 411.600 219.800 ;
        RECT 407.600 215.800 411.600 216.000 ;
        RECT 414.000 217.800 414.800 219.800 ;
        RECT 361.200 214.200 362.800 214.400 ;
        RECT 351.800 213.600 362.800 214.200 ;
        RECT 364.400 213.600 367.000 214.400 ;
        RECT 368.400 213.800 370.000 214.400 ;
        RECT 369.200 213.600 370.000 213.800 ;
        RECT 350.000 212.800 350.800 213.000 ;
        RECT 347.000 212.200 350.800 212.800 ;
        RECT 347.000 212.000 347.800 212.200 ;
        RECT 348.600 211.400 349.400 211.600 ;
        RECT 345.200 210.800 349.400 211.400 ;
        RECT 345.200 202.200 346.000 210.800 ;
        RECT 351.800 210.400 352.400 213.600 ;
        RECT 359.000 213.400 359.800 213.600 ;
        RECT 358.000 212.400 358.800 212.600 ;
        RECT 360.600 212.400 361.400 212.600 ;
        RECT 356.400 211.800 361.400 212.400 ;
        RECT 356.400 211.600 357.200 211.800 ;
        RECT 358.000 211.000 363.600 211.200 ;
        RECT 357.800 210.800 363.600 211.000 ;
        RECT 350.000 209.800 352.400 210.400 ;
        RECT 353.800 210.600 363.600 210.800 ;
        RECT 353.800 210.200 358.600 210.600 ;
        RECT 350.000 208.800 350.600 209.800 ;
        RECT 349.200 208.000 350.600 208.800 ;
        RECT 352.200 209.000 353.000 209.200 ;
        RECT 353.800 209.000 354.400 210.200 ;
        RECT 352.200 208.400 354.400 209.000 ;
        RECT 355.000 209.000 360.400 209.600 ;
        RECT 355.000 208.800 355.800 209.000 ;
        RECT 359.600 208.800 360.400 209.000 ;
        RECT 353.400 207.400 354.200 207.600 ;
        RECT 356.200 207.400 357.000 207.600 ;
        RECT 350.000 206.200 350.800 207.000 ;
        RECT 353.400 206.800 357.000 207.400 ;
        RECT 354.200 206.200 354.800 206.800 ;
        RECT 359.600 206.200 360.400 207.000 ;
        RECT 349.400 202.200 350.600 206.200 ;
        RECT 354.000 202.200 354.800 206.200 ;
        RECT 358.400 205.600 360.400 206.200 ;
        RECT 358.400 202.200 359.200 205.600 ;
        RECT 362.800 202.200 363.600 210.600 ;
        RECT 364.400 210.200 365.200 210.400 ;
        RECT 366.400 210.200 367.000 213.600 ;
        RECT 367.600 211.600 368.400 213.200 ;
        RECT 370.800 212.800 371.600 214.400 ;
        RECT 372.400 213.800 374.800 214.400 ;
        RECT 376.400 214.300 378.000 214.400 ;
        RECT 378.800 214.300 379.600 214.400 ;
        RECT 376.400 213.800 379.600 214.300 ;
        RECT 374.000 213.600 374.800 213.800 ;
        RECT 377.200 213.700 379.600 213.800 ;
        RECT 377.200 213.600 378.000 213.700 ;
        RECT 378.800 213.600 379.600 213.700 ;
        RECT 380.400 213.600 381.200 214.400 ;
        RECT 372.400 211.600 373.200 213.200 ;
        RECT 374.200 210.200 374.800 213.600 ;
        RECT 375.600 212.300 376.400 213.200 ;
        RECT 377.200 212.300 378.000 212.400 ;
        RECT 375.600 211.700 378.000 212.300 ;
        RECT 375.600 211.600 376.400 211.700 ;
        RECT 377.200 211.600 378.000 211.700 ;
        RECT 378.800 212.200 379.600 212.400 ;
        RECT 380.600 212.200 381.200 213.600 ;
        RECT 382.000 212.800 382.800 214.400 ;
        RECT 385.200 213.600 386.000 215.200 ;
        RECT 383.600 212.200 384.400 212.400 ;
        RECT 378.800 211.600 381.200 212.200 ;
        RECT 382.800 211.600 384.400 212.200 ;
        RECT 379.000 210.200 379.600 211.600 ;
        RECT 382.800 211.200 383.600 211.600 ;
        RECT 364.400 209.600 365.800 210.200 ;
        RECT 366.400 209.600 367.400 210.200 ;
        RECT 365.200 208.400 365.800 209.600 ;
        RECT 365.200 207.600 366.000 208.400 ;
        RECT 366.600 202.200 367.400 209.600 ;
        RECT 373.400 202.200 375.400 210.200 ;
        RECT 378.800 202.200 379.600 210.200 ;
        RECT 380.400 209.600 384.400 210.200 ;
        RECT 380.400 202.200 381.200 209.600 ;
        RECT 383.600 202.200 384.400 209.600 ;
        RECT 386.800 202.200 387.600 215.800 ;
        RECT 390.200 215.400 393.800 215.800 ;
        RECT 390.800 214.400 391.600 214.800 ;
        RECT 394.800 214.400 395.400 215.800 ;
        RECT 398.000 214.400 398.600 215.800 ;
        RECT 399.800 215.400 403.400 215.800 ;
        RECT 402.000 214.400 402.800 214.800 ;
        RECT 406.000 214.400 406.600 215.800 ;
        RECT 407.800 215.400 411.400 215.800 ;
        RECT 410.000 214.400 410.800 214.800 ;
        RECT 414.000 214.400 414.600 217.800 ;
        RECT 415.600 215.600 416.400 217.200 ;
        RECT 417.200 215.800 418.000 219.800 ;
        RECT 418.800 216.000 419.600 219.800 ;
        RECT 422.000 216.000 422.800 219.800 ;
        RECT 418.800 215.800 422.800 216.000 ;
        RECT 432.600 215.800 434.200 219.800 ;
        RECT 439.600 217.800 440.400 219.800 ;
        RECT 417.400 214.400 418.000 215.800 ;
        RECT 419.000 215.400 422.600 215.800 ;
        RECT 421.200 214.400 422.000 214.800 ;
        RECT 390.000 213.800 391.600 214.400 ;
        RECT 390.000 213.600 390.800 213.800 ;
        RECT 393.000 213.600 395.600 214.400 ;
        RECT 391.600 211.600 392.400 213.200 ;
        RECT 388.400 208.800 389.200 210.400 ;
        RECT 393.000 210.200 393.600 213.600 ;
        RECT 396.400 212.800 397.200 214.400 ;
        RECT 398.000 213.800 400.400 214.400 ;
        RECT 402.000 213.800 403.600 214.400 ;
        RECT 399.600 213.600 400.400 213.800 ;
        RECT 402.800 213.600 403.600 213.800 ;
        RECT 398.000 211.600 398.800 213.200 ;
        RECT 394.800 210.200 395.600 210.400 ;
        RECT 399.800 210.200 400.400 213.600 ;
        RECT 401.200 211.600 402.000 213.200 ;
        RECT 404.400 212.800 405.200 214.400 ;
        RECT 406.000 213.800 408.400 214.400 ;
        RECT 410.000 213.800 411.600 214.400 ;
        RECT 407.600 213.600 408.400 213.800 ;
        RECT 410.800 213.600 411.600 213.800 ;
        RECT 414.000 213.600 414.800 214.400 ;
        RECT 415.600 214.300 416.400 214.400 ;
        RECT 417.200 214.300 419.800 214.400 ;
        RECT 415.600 213.700 419.800 214.300 ;
        RECT 421.200 214.300 422.800 214.400 ;
        RECT 423.600 214.300 424.400 214.400 ;
        RECT 421.200 213.800 424.400 214.300 ;
        RECT 415.600 213.600 416.400 213.700 ;
        RECT 417.200 213.600 419.800 213.700 ;
        RECT 422.000 213.700 424.400 213.800 ;
        RECT 422.000 213.600 422.800 213.700 ;
        RECT 423.600 213.600 424.400 213.700 ;
        RECT 428.400 214.300 429.200 214.400 ;
        RECT 431.600 214.300 432.400 214.400 ;
        RECT 428.400 213.700 432.400 214.300 ;
        RECT 428.400 213.600 429.200 213.700 ;
        RECT 431.600 213.600 432.400 213.700 ;
        RECT 406.000 211.600 406.800 213.200 ;
        RECT 407.800 210.200 408.400 213.600 ;
        RECT 409.200 211.600 410.000 213.200 ;
        RECT 412.400 210.800 413.200 212.400 ;
        RECT 414.000 210.200 414.600 213.600 ;
        RECT 417.200 210.200 418.000 210.400 ;
        RECT 419.200 210.200 419.800 213.600 ;
        RECT 431.800 213.200 432.400 213.600 ;
        RECT 420.400 212.300 421.200 213.200 ;
        RECT 431.800 212.400 432.600 213.200 ;
        RECT 433.200 212.400 433.800 215.800 ;
        RECT 438.000 215.600 438.800 217.200 ;
        RECT 439.800 216.300 440.400 217.800 ;
        RECT 444.400 217.800 445.200 219.800 ;
        RECT 447.600 219.200 451.600 219.800 ;
        RECT 441.200 216.300 442.000 216.400 ;
        RECT 439.700 215.700 442.000 216.300 ;
        RECT 439.800 214.400 440.400 215.700 ;
        RECT 441.200 215.600 442.000 215.700 ;
        RECT 434.800 212.800 435.600 214.400 ;
        RECT 439.600 213.600 440.400 214.400 ;
        RECT 428.400 212.300 429.200 212.400 ;
        RECT 420.400 211.700 429.200 212.300 ;
        RECT 420.400 211.600 421.200 211.700 ;
        RECT 428.400 211.600 429.200 211.700 ;
        RECT 430.000 210.800 430.800 212.400 ;
        RECT 433.200 211.600 434.000 212.400 ;
        RECT 436.400 212.200 437.200 212.400 ;
        RECT 435.600 211.600 437.200 212.200 ;
        RECT 433.200 211.400 433.800 211.600 ;
        RECT 431.800 210.800 433.800 211.400 ;
        RECT 435.600 211.200 436.400 211.600 ;
        RECT 431.800 210.200 432.400 210.800 ;
        RECT 439.800 210.200 440.400 213.600 ;
        RECT 444.400 214.400 445.000 217.800 ;
        RECT 446.000 215.600 446.800 217.200 ;
        RECT 447.600 215.800 448.400 219.200 ;
        RECT 449.200 215.800 450.000 218.600 ;
        RECT 450.800 216.000 451.600 219.200 ;
        RECT 454.000 216.000 454.800 219.800 ;
        RECT 450.800 215.800 454.800 216.000 ;
        RECT 455.600 216.000 456.400 219.800 ;
        RECT 458.800 219.200 462.800 219.800 ;
        RECT 458.800 216.000 459.600 219.200 ;
        RECT 455.600 215.800 459.600 216.000 ;
        RECT 460.400 215.800 461.200 218.600 ;
        RECT 462.000 215.800 462.800 219.200 ;
        RECT 463.600 217.000 464.400 219.000 ;
        RECT 449.200 214.400 449.800 215.800 ;
        RECT 451.000 215.400 454.600 215.800 ;
        RECT 455.800 215.400 459.400 215.800 ;
        RECT 453.200 214.400 454.000 214.800 ;
        RECT 456.400 214.400 457.200 214.800 ;
        RECT 460.600 214.400 461.200 215.800 ;
        RECT 463.600 214.800 464.200 217.000 ;
        RECT 467.800 216.000 468.600 219.000 ;
        RECT 473.200 216.000 474.000 219.800 ;
        RECT 476.400 216.000 477.200 219.800 ;
        RECT 467.800 215.400 469.400 216.000 ;
        RECT 473.200 215.800 477.200 216.000 ;
        RECT 478.000 215.800 478.800 219.800 ;
        RECT 481.200 216.000 482.000 219.800 ;
        RECT 473.400 215.400 477.000 215.800 ;
        RECT 468.600 215.000 469.400 215.400 ;
        RECT 444.400 213.600 445.200 214.400 ;
        RECT 441.200 210.800 442.000 212.400 ;
        RECT 442.800 210.800 443.600 212.400 ;
        RECT 444.400 210.200 445.000 213.600 ;
        RECT 447.600 212.800 448.400 214.400 ;
        RECT 449.200 213.800 451.600 214.400 ;
        RECT 453.200 213.800 454.800 214.400 ;
        RECT 450.800 213.600 451.600 213.800 ;
        RECT 454.000 213.600 454.800 213.800 ;
        RECT 455.600 213.800 457.200 214.400 ;
        RECT 458.800 213.800 461.200 214.400 ;
        RECT 455.600 213.600 456.400 213.800 ;
        RECT 458.800 213.600 459.600 213.800 ;
        RECT 449.200 211.600 450.000 213.200 ;
        RECT 451.000 210.200 451.600 213.600 ;
        RECT 452.400 212.300 453.200 213.200 ;
        RECT 457.200 212.300 458.000 213.200 ;
        RECT 452.400 211.700 458.000 212.300 ;
        RECT 452.400 211.600 453.200 211.700 ;
        RECT 457.200 211.600 458.000 211.700 ;
        RECT 458.800 210.200 459.400 213.600 ;
        RECT 460.400 211.600 461.200 213.200 ;
        RECT 462.000 212.800 462.800 214.400 ;
        RECT 463.600 214.200 467.800 214.800 ;
        RECT 466.800 213.800 467.800 214.200 ;
        RECT 468.800 214.400 469.400 215.000 ;
        RECT 474.000 214.400 474.800 214.800 ;
        RECT 478.000 214.400 478.600 215.800 ;
        RECT 481.000 215.200 482.000 216.000 ;
        RECT 463.600 211.600 464.400 213.200 ;
        RECT 465.200 211.600 466.000 213.200 ;
        RECT 466.800 213.000 468.200 213.800 ;
        RECT 468.800 213.600 470.800 214.400 ;
        RECT 473.200 213.800 474.800 214.400 ;
        RECT 473.200 213.600 474.000 213.800 ;
        RECT 476.200 213.600 478.800 214.400 ;
        RECT 466.800 211.000 467.400 213.000 ;
        RECT 463.600 210.400 467.400 211.000 ;
        RECT 392.600 209.600 393.600 210.200 ;
        RECT 394.200 209.600 395.600 210.200 ;
        RECT 392.600 202.200 393.400 209.600 ;
        RECT 394.200 208.400 394.800 209.600 ;
        RECT 394.000 207.600 394.800 208.400 ;
        RECT 399.000 204.400 401.000 210.200 ;
        RECT 399.000 203.600 402.000 204.400 ;
        RECT 399.000 202.200 401.000 203.600 ;
        RECT 407.000 202.200 409.000 210.200 ;
        RECT 413.000 209.400 414.800 210.200 ;
        RECT 417.200 209.600 418.600 210.200 ;
        RECT 419.200 209.600 420.200 210.200 ;
        RECT 413.000 204.400 413.800 209.400 ;
        RECT 418.000 208.400 418.600 209.600 ;
        RECT 418.000 207.600 418.800 208.400 ;
        RECT 413.000 203.600 414.800 204.400 ;
        RECT 413.000 202.200 413.800 203.600 ;
        RECT 419.400 202.200 420.200 209.600 ;
        RECT 430.000 202.800 430.800 210.200 ;
        RECT 431.600 203.400 432.400 210.200 ;
        RECT 433.200 209.600 437.200 210.200 ;
        RECT 433.200 202.800 434.000 209.600 ;
        RECT 430.000 202.200 434.000 202.800 ;
        RECT 436.400 202.200 437.200 209.600 ;
        RECT 439.600 209.400 441.400 210.200 ;
        RECT 440.600 202.200 441.400 209.400 ;
        RECT 443.400 209.400 445.200 210.200 ;
        RECT 443.400 208.400 444.200 209.400 ;
        RECT 450.200 208.400 452.200 210.200 ;
        RECT 443.400 207.600 445.200 208.400 ;
        RECT 449.200 207.600 452.200 208.400 ;
        RECT 443.400 202.200 444.200 207.600 ;
        RECT 450.200 202.200 452.200 207.600 ;
        RECT 458.200 202.200 460.200 210.200 ;
        RECT 463.600 207.000 464.200 210.400 ;
        RECT 468.800 209.800 469.400 213.600 ;
        RECT 470.000 212.300 470.800 212.400 ;
        RECT 471.600 212.300 472.400 212.400 ;
        RECT 470.000 211.700 472.400 212.300 ;
        RECT 470.000 210.800 470.800 211.700 ;
        RECT 471.600 211.600 472.400 211.700 ;
        RECT 474.800 211.600 475.600 213.200 ;
        RECT 476.200 212.400 476.800 213.600 ;
        RECT 476.200 211.600 477.200 212.400 ;
        RECT 476.200 210.200 476.800 211.600 ;
        RECT 481.000 210.800 481.800 215.200 ;
        RECT 482.800 214.600 483.600 219.800 ;
        RECT 489.200 216.600 490.000 219.800 ;
        RECT 490.800 217.000 491.600 219.800 ;
        RECT 492.400 217.000 493.200 219.800 ;
        RECT 494.000 217.000 494.800 219.800 ;
        RECT 495.600 217.000 496.400 219.800 ;
        RECT 498.800 217.000 499.600 219.800 ;
        RECT 502.000 217.000 502.800 219.800 ;
        RECT 503.600 217.000 504.400 219.800 ;
        RECT 505.200 217.000 506.000 219.800 ;
        RECT 487.600 215.800 490.000 216.600 ;
        RECT 506.800 216.600 507.600 219.800 ;
        RECT 487.600 215.200 488.400 215.800 ;
        RECT 482.400 214.000 483.600 214.600 ;
        RECT 486.600 214.600 488.400 215.200 ;
        RECT 492.400 215.600 493.400 216.400 ;
        RECT 496.400 215.600 498.000 216.400 ;
        RECT 498.800 215.800 503.400 216.400 ;
        RECT 506.800 215.800 509.400 216.600 ;
        RECT 498.800 215.600 499.600 215.800 ;
        RECT 482.400 212.000 483.000 214.000 ;
        RECT 486.600 213.400 487.400 214.600 ;
        RECT 483.600 212.600 487.400 213.400 ;
        RECT 492.400 212.800 493.200 215.600 ;
        RECT 498.800 214.800 499.600 215.000 ;
        RECT 495.200 214.200 499.600 214.800 ;
        RECT 495.200 214.000 496.000 214.200 ;
        RECT 500.400 213.600 501.200 215.200 ;
        RECT 502.600 213.400 503.400 215.800 ;
        RECT 508.600 215.200 509.400 215.800 ;
        RECT 508.600 214.400 511.600 215.200 ;
        RECT 513.200 213.800 514.000 219.800 ;
        RECT 495.600 212.600 498.800 213.400 ;
        RECT 502.600 212.600 504.600 213.400 ;
        RECT 505.200 213.000 514.000 213.800 ;
        RECT 489.200 212.000 490.000 212.600 ;
        RECT 506.800 212.000 507.600 212.400 ;
        RECT 511.800 212.000 512.600 212.200 ;
        RECT 482.400 211.400 483.200 212.000 ;
        RECT 489.200 211.400 512.600 212.000 ;
        RECT 478.000 210.200 478.800 210.400 ;
        RECT 467.800 209.200 469.400 209.800 ;
        RECT 475.800 209.600 476.800 210.200 ;
        RECT 477.400 209.600 478.800 210.200 ;
        RECT 481.000 210.000 482.000 210.800 ;
        RECT 463.600 203.000 464.400 207.000 ;
        RECT 467.800 204.400 468.600 209.200 ;
        RECT 467.800 203.600 469.200 204.400 ;
        RECT 467.800 202.200 468.600 203.600 ;
        RECT 475.800 202.200 476.600 209.600 ;
        RECT 477.400 208.400 478.000 209.600 ;
        RECT 477.200 207.600 478.000 208.400 ;
        RECT 481.200 202.200 482.000 210.000 ;
        RECT 482.600 209.600 483.200 211.400 ;
        RECT 482.600 209.000 491.600 209.600 ;
        RECT 482.600 207.400 483.200 209.000 ;
        RECT 490.800 208.800 491.600 209.000 ;
        RECT 494.000 209.000 502.600 209.600 ;
        RECT 494.000 208.800 494.800 209.000 ;
        RECT 485.800 207.600 488.400 208.400 ;
        RECT 482.600 206.800 485.200 207.400 ;
        RECT 484.400 202.200 485.200 206.800 ;
        RECT 487.600 202.200 488.400 207.600 ;
        RECT 489.000 206.800 493.200 207.600 ;
        RECT 490.800 202.200 491.600 205.000 ;
        RECT 492.400 202.200 493.200 205.000 ;
        RECT 494.000 202.200 494.800 205.000 ;
        RECT 495.600 202.200 496.400 208.400 ;
        RECT 498.800 207.600 501.400 208.400 ;
        RECT 502.000 208.200 502.600 209.000 ;
        RECT 503.600 209.400 504.400 209.600 ;
        RECT 503.600 209.000 509.000 209.400 ;
        RECT 503.600 208.800 509.800 209.000 ;
        RECT 508.400 208.200 509.800 208.800 ;
        RECT 502.000 207.600 507.800 208.200 ;
        RECT 510.800 208.000 512.400 208.800 ;
        RECT 510.800 207.600 511.400 208.000 ;
        RECT 498.800 202.200 499.600 207.000 ;
        RECT 502.000 202.200 502.800 207.000 ;
        RECT 507.200 206.800 511.400 207.600 ;
        RECT 513.200 207.400 514.000 213.000 ;
        RECT 512.000 206.800 514.000 207.400 ;
        RECT 514.800 213.800 515.600 219.800 ;
        RECT 521.200 216.600 522.000 219.800 ;
        RECT 522.800 217.000 523.600 219.800 ;
        RECT 524.400 217.000 525.200 219.800 ;
        RECT 526.000 217.000 526.800 219.800 ;
        RECT 529.200 217.000 530.000 219.800 ;
        RECT 532.400 217.000 533.200 219.800 ;
        RECT 534.000 217.000 534.800 219.800 ;
        RECT 535.600 217.000 536.400 219.800 ;
        RECT 537.200 217.000 538.000 219.800 ;
        RECT 519.400 215.800 522.000 216.600 ;
        RECT 538.800 216.600 539.600 219.800 ;
        RECT 525.400 215.800 530.000 216.400 ;
        RECT 519.400 215.200 520.200 215.800 ;
        RECT 517.200 214.400 520.200 215.200 ;
        RECT 514.800 213.000 523.600 213.800 ;
        RECT 525.400 213.400 526.200 215.800 ;
        RECT 529.200 215.600 530.000 215.800 ;
        RECT 530.800 215.600 532.400 216.400 ;
        RECT 535.400 215.600 536.400 216.400 ;
        RECT 538.800 215.800 541.200 216.600 ;
        RECT 527.600 213.600 528.400 215.200 ;
        RECT 529.200 214.800 530.000 215.000 ;
        RECT 529.200 214.200 533.600 214.800 ;
        RECT 532.800 214.000 533.600 214.200 ;
        RECT 514.800 207.400 515.600 213.000 ;
        RECT 524.200 212.600 526.200 213.400 ;
        RECT 530.000 212.600 533.200 213.400 ;
        RECT 535.600 212.800 536.400 215.600 ;
        RECT 540.400 215.200 541.200 215.800 ;
        RECT 540.400 214.600 542.200 215.200 ;
        RECT 541.400 213.400 542.200 214.600 ;
        RECT 545.200 214.600 546.000 219.800 ;
        RECT 546.800 216.000 547.600 219.800 ;
        RECT 546.800 215.200 547.800 216.000 ;
        RECT 545.200 214.000 546.400 214.600 ;
        RECT 541.400 212.600 545.200 213.400 ;
        RECT 516.200 212.000 517.000 212.200 ;
        RECT 518.000 212.000 518.800 212.400 ;
        RECT 521.200 212.000 522.000 212.400 ;
        RECT 538.800 212.000 539.600 212.600 ;
        RECT 545.800 212.000 546.400 214.000 ;
        RECT 516.200 211.400 539.600 212.000 ;
        RECT 545.600 211.400 546.400 212.000 ;
        RECT 545.600 209.600 546.200 211.400 ;
        RECT 547.000 210.800 547.800 215.200 ;
        RECT 524.400 209.400 525.200 209.600 ;
        RECT 519.800 209.000 525.200 209.400 ;
        RECT 519.000 208.800 525.200 209.000 ;
        RECT 526.200 209.000 534.800 209.600 ;
        RECT 516.400 208.000 518.000 208.800 ;
        RECT 519.000 208.200 520.400 208.800 ;
        RECT 526.200 208.200 526.800 209.000 ;
        RECT 534.000 208.800 534.800 209.000 ;
        RECT 537.200 209.000 546.200 209.600 ;
        RECT 537.200 208.800 538.000 209.000 ;
        RECT 517.400 207.600 518.000 208.000 ;
        RECT 521.000 207.600 526.800 208.200 ;
        RECT 527.400 207.600 530.000 208.400 ;
        RECT 514.800 206.800 516.800 207.400 ;
        RECT 517.400 206.800 521.600 207.600 ;
        RECT 503.600 202.200 504.400 205.000 ;
        RECT 505.200 202.200 506.000 205.000 ;
        RECT 508.400 202.200 509.200 206.800 ;
        RECT 512.000 206.200 512.600 206.800 ;
        RECT 511.600 205.600 512.600 206.200 ;
        RECT 516.200 206.200 516.800 206.800 ;
        RECT 516.200 205.600 517.200 206.200 ;
        RECT 511.600 202.200 512.400 205.600 ;
        RECT 516.400 202.200 517.200 205.600 ;
        RECT 519.600 202.200 520.400 206.800 ;
        RECT 522.800 202.200 523.600 205.000 ;
        RECT 524.400 202.200 525.200 205.000 ;
        RECT 526.000 202.200 526.800 207.000 ;
        RECT 529.200 202.200 530.000 207.000 ;
        RECT 532.400 202.200 533.200 208.400 ;
        RECT 540.400 207.600 543.000 208.400 ;
        RECT 535.600 206.800 539.800 207.600 ;
        RECT 534.000 202.200 534.800 205.000 ;
        RECT 535.600 202.200 536.400 205.000 ;
        RECT 537.200 202.200 538.000 205.000 ;
        RECT 540.400 202.200 541.200 207.600 ;
        RECT 545.600 207.400 546.200 209.000 ;
        RECT 543.600 206.800 546.200 207.400 ;
        RECT 546.800 210.000 547.800 210.800 ;
        RECT 546.800 208.300 547.600 210.000 ;
        RECT 550.000 208.300 550.800 208.400 ;
        RECT 546.800 207.700 550.800 208.300 ;
        RECT 543.600 202.200 544.400 206.800 ;
        RECT 546.800 202.200 547.600 207.700 ;
        RECT 550.000 207.600 550.800 207.700 ;
        RECT 1.200 186.800 2.000 188.400 ;
        RECT 2.800 186.200 3.600 199.800 ;
        RECT 4.400 191.600 5.200 193.200 ;
        RECT 6.000 191.600 6.800 193.200 ;
        RECT 7.600 186.200 8.400 199.800 ;
        RECT 11.400 192.600 12.200 199.800 ;
        RECT 17.200 195.800 18.000 199.800 ;
        RECT 11.400 191.800 13.200 192.600 ;
        RECT 10.800 189.600 11.600 191.200 ;
        RECT 12.400 188.400 13.000 191.800 ;
        RECT 17.400 191.600 18.000 195.800 ;
        RECT 20.400 191.800 21.200 199.800 ;
        RECT 24.600 192.600 25.400 199.800 ;
        RECT 23.600 191.800 25.400 192.600 ;
        RECT 17.400 191.000 19.800 191.600 ;
        RECT 17.200 189.600 18.000 190.400 ;
        RECT 9.200 186.800 10.000 188.400 ;
        RECT 12.400 188.300 13.200 188.400 ;
        RECT 15.600 188.300 16.400 189.200 ;
        RECT 17.400 188.800 18.000 189.600 ;
        RECT 12.400 187.700 16.400 188.300 ;
        RECT 17.200 188.000 18.400 188.800 ;
        RECT 12.400 187.600 13.200 187.700 ;
        RECT 15.600 187.600 16.400 187.700 ;
        RECT 19.200 187.600 19.800 191.000 ;
        RECT 20.600 190.400 21.200 191.800 ;
        RECT 20.400 189.600 21.200 190.400 ;
        RECT 22.000 190.300 22.800 190.400 ;
        RECT 23.800 190.300 24.400 191.800 ;
        RECT 26.800 191.200 27.600 199.800 ;
        RECT 31.000 196.400 31.800 199.800 ;
        RECT 31.000 195.600 32.400 196.400 ;
        RECT 34.800 195.800 35.600 199.800 ;
        RECT 35.000 195.600 35.600 195.800 ;
        RECT 38.000 195.800 38.800 199.800 ;
        RECT 39.600 195.800 40.400 199.800 ;
        RECT 38.000 195.600 38.600 195.800 ;
        RECT 31.000 192.400 31.800 195.600 ;
        RECT 35.000 195.000 38.600 195.600 ;
        RECT 36.400 192.800 37.200 194.400 ;
        RECT 38.000 192.400 38.600 195.000 ;
        RECT 39.800 195.600 40.400 195.800 ;
        RECT 42.800 195.800 43.600 199.800 ;
        RECT 42.800 195.600 43.400 195.800 ;
        RECT 39.800 195.000 43.400 195.600 ;
        RECT 39.800 192.400 40.400 195.000 ;
        RECT 41.200 192.800 42.000 194.400 ;
        RECT 31.000 191.800 32.400 192.400 ;
        RECT 22.000 189.700 24.400 190.300 ;
        RECT 22.000 189.600 22.800 189.700 ;
        RECT 2.800 185.600 4.600 186.200 ;
        RECT 3.800 184.400 4.600 185.600 ;
        RECT 6.600 185.600 8.400 186.200 ;
        RECT 6.600 184.400 7.400 185.600 ;
        RECT 3.800 183.600 5.200 184.400 ;
        RECT 6.600 183.600 8.400 184.400 ;
        RECT 12.400 184.200 13.000 187.600 ;
        RECT 19.200 187.400 20.000 187.600 ;
        RECT 17.000 187.000 20.000 187.400 ;
        RECT 15.800 186.800 20.000 187.000 ;
        RECT 15.800 186.400 17.600 186.800 ;
        RECT 14.000 184.800 14.800 186.400 ;
        RECT 15.800 186.200 16.400 186.400 ;
        RECT 20.600 186.200 21.200 189.600 ;
        RECT 23.800 188.400 24.400 189.700 ;
        RECT 25.200 189.600 26.000 191.200 ;
        RECT 26.800 190.800 30.800 191.200 ;
        RECT 26.800 190.600 31.000 190.800 ;
        RECT 30.200 190.000 31.000 190.600 ;
        RECT 31.800 190.400 32.400 191.800 ;
        RECT 33.200 190.800 34.000 192.400 ;
        RECT 38.000 191.600 38.800 192.400 ;
        RECT 39.600 191.600 40.400 192.400 ;
        RECT 28.800 188.400 29.600 189.200 ;
        RECT 23.600 187.600 24.400 188.400 ;
        RECT 28.400 187.600 29.400 188.400 ;
        RECT 3.800 182.200 4.600 183.600 ;
        RECT 6.600 182.200 7.400 183.600 ;
        RECT 12.400 182.200 13.200 184.200 ;
        RECT 15.600 182.200 16.400 186.200 ;
        RECT 19.800 185.200 21.200 186.200 ;
        RECT 19.800 184.400 20.600 185.200 ;
        RECT 22.000 184.800 22.800 186.400 ;
        RECT 19.800 183.600 21.200 184.400 ;
        RECT 23.800 184.200 24.400 187.600 ;
        RECT 30.400 187.000 31.000 190.000 ;
        RECT 31.600 189.600 32.400 190.400 ;
        RECT 34.800 189.600 36.400 190.400 ;
        RECT 28.600 186.400 31.000 187.000 ;
        RECT 26.800 184.800 27.600 186.400 ;
        RECT 28.600 184.200 29.200 186.400 ;
        RECT 31.800 186.200 32.400 189.600 ;
        RECT 38.000 188.400 38.600 191.600 ;
        RECT 34.800 188.300 35.600 188.400 ;
        RECT 37.000 188.300 38.600 188.400 ;
        RECT 34.800 187.800 38.600 188.300 ;
        RECT 39.800 188.400 40.400 191.600 ;
        RECT 44.400 190.800 45.200 192.400 ;
        RECT 42.000 189.600 43.600 190.400 ;
        RECT 39.800 188.200 41.400 188.400 ;
        RECT 39.800 187.800 41.600 188.200 ;
        RECT 34.800 187.700 37.600 187.800 ;
        RECT 34.800 187.600 35.600 187.700 ;
        RECT 36.400 187.600 37.600 187.700 ;
        RECT 19.800 182.200 20.600 183.600 ;
        RECT 23.600 182.200 24.400 184.200 ;
        RECT 28.400 182.200 29.200 184.200 ;
        RECT 31.600 182.200 32.400 186.200 ;
        RECT 36.800 182.200 37.600 187.600 ;
        RECT 40.800 182.200 41.600 187.800 ;
        RECT 46.000 184.800 46.800 186.400 ;
        RECT 47.600 182.200 48.400 199.800 ;
        RECT 49.200 186.800 50.000 188.400 ;
        RECT 50.800 186.200 51.600 199.800 ;
        RECT 54.000 195.800 54.800 199.800 ;
        RECT 54.200 195.600 54.800 195.800 ;
        RECT 57.200 195.800 58.000 199.800 ;
        RECT 62.000 195.800 62.800 199.800 ;
        RECT 57.200 195.600 57.800 195.800 ;
        RECT 54.200 195.000 57.800 195.600 ;
        RECT 52.400 191.600 53.200 193.200 ;
        RECT 54.200 192.400 54.800 195.000 ;
        RECT 55.600 192.800 56.400 194.400 ;
        RECT 54.000 191.600 54.800 192.400 ;
        RECT 54.200 188.400 54.800 191.600 ;
        RECT 58.800 190.800 59.600 192.400 ;
        RECT 62.200 191.600 62.800 195.800 ;
        RECT 65.200 191.800 66.000 199.800 ;
        RECT 68.400 196.400 69.200 199.800 ;
        RECT 68.200 195.800 69.200 196.400 ;
        RECT 68.200 195.200 68.800 195.800 ;
        RECT 71.600 195.200 72.400 199.800 ;
        RECT 74.800 197.000 75.600 199.800 ;
        RECT 76.400 197.000 77.200 199.800 ;
        RECT 62.200 191.000 64.600 191.600 ;
        RECT 56.400 189.600 58.000 190.400 ;
        RECT 62.000 189.600 62.800 190.400 ;
        RECT 54.200 188.200 55.800 188.400 ;
        RECT 54.200 187.800 56.000 188.200 ;
        RECT 50.800 185.600 52.600 186.200 ;
        RECT 51.800 184.400 52.600 185.600 ;
        RECT 51.800 183.600 53.200 184.400 ;
        RECT 51.800 182.200 52.600 183.600 ;
        RECT 55.200 182.200 56.000 187.800 ;
        RECT 60.400 187.600 61.200 189.200 ;
        RECT 62.200 188.800 62.800 189.600 ;
        RECT 62.200 188.200 63.200 188.800 ;
        RECT 62.400 188.000 63.200 188.200 ;
        RECT 64.000 187.600 64.600 191.000 ;
        RECT 65.400 190.400 66.000 191.800 ;
        RECT 65.200 189.600 66.000 190.400 ;
        RECT 64.000 187.400 64.800 187.600 ;
        RECT 61.800 187.000 64.800 187.400 ;
        RECT 60.600 186.800 64.800 187.000 ;
        RECT 60.600 186.400 62.400 186.800 ;
        RECT 60.600 186.200 61.200 186.400 ;
        RECT 65.400 186.200 66.000 189.600 ;
        RECT 60.400 182.200 61.200 186.200 ;
        RECT 64.600 185.200 66.000 186.200 ;
        RECT 66.800 194.600 68.800 195.200 ;
        RECT 66.800 189.000 67.600 194.600 ;
        RECT 69.400 194.400 73.600 195.200 ;
        RECT 78.000 195.000 78.800 199.800 ;
        RECT 81.200 195.000 82.000 199.800 ;
        RECT 69.400 194.000 70.000 194.400 ;
        RECT 68.400 193.200 70.000 194.000 ;
        RECT 73.000 193.800 78.800 194.400 ;
        RECT 71.000 193.200 72.400 193.800 ;
        RECT 71.000 193.000 77.200 193.200 ;
        RECT 71.800 192.600 77.200 193.000 ;
        RECT 76.400 192.400 77.200 192.600 ;
        RECT 78.200 193.000 78.800 193.800 ;
        RECT 79.400 193.600 82.000 194.400 ;
        RECT 84.400 193.600 85.200 199.800 ;
        RECT 86.000 197.000 86.800 199.800 ;
        RECT 87.600 197.000 88.400 199.800 ;
        RECT 89.200 197.000 90.000 199.800 ;
        RECT 87.600 194.400 91.800 195.200 ;
        RECT 92.400 194.400 93.200 199.800 ;
        RECT 95.600 195.200 96.400 199.800 ;
        RECT 95.600 194.600 98.200 195.200 ;
        RECT 92.400 193.600 95.000 194.400 ;
        RECT 86.000 193.000 86.800 193.200 ;
        RECT 78.200 192.400 86.800 193.000 ;
        RECT 89.200 193.000 90.000 193.200 ;
        RECT 97.600 193.000 98.200 194.600 ;
        RECT 89.200 192.400 98.200 193.000 ;
        RECT 97.600 190.600 98.200 192.400 ;
        RECT 98.800 192.000 99.600 199.800 ;
        RECT 103.600 192.000 104.400 199.800 ;
        RECT 106.800 195.200 107.600 199.800 ;
        RECT 98.800 191.200 99.800 192.000 ;
        RECT 68.200 190.000 91.600 190.600 ;
        RECT 97.600 190.000 98.400 190.600 ;
        RECT 68.200 189.800 69.000 190.000 ;
        RECT 73.200 189.600 74.000 190.000 ;
        RECT 90.800 189.400 91.600 190.000 ;
        RECT 66.800 188.200 75.600 189.000 ;
        RECT 76.200 188.600 78.200 189.400 ;
        RECT 82.000 188.600 85.200 189.400 ;
        RECT 64.600 182.200 65.400 185.200 ;
        RECT 66.800 182.200 67.600 188.200 ;
        RECT 69.200 186.800 72.200 187.600 ;
        RECT 71.400 186.200 72.200 186.800 ;
        RECT 77.400 186.200 78.200 188.600 ;
        RECT 79.600 186.800 80.400 188.400 ;
        RECT 84.800 187.800 85.600 188.000 ;
        RECT 81.200 187.200 85.600 187.800 ;
        RECT 81.200 187.000 82.000 187.200 ;
        RECT 87.600 186.400 88.400 189.200 ;
        RECT 93.400 188.600 97.200 189.400 ;
        RECT 93.400 187.400 94.200 188.600 ;
        RECT 97.800 188.000 98.400 190.000 ;
        RECT 81.200 186.200 82.000 186.400 ;
        RECT 71.400 185.400 74.000 186.200 ;
        RECT 77.400 185.600 82.000 186.200 ;
        RECT 82.800 185.600 84.400 186.400 ;
        RECT 87.400 185.600 88.400 186.400 ;
        RECT 92.400 186.800 94.200 187.400 ;
        RECT 97.200 187.400 98.400 188.000 ;
        RECT 92.400 186.200 93.200 186.800 ;
        RECT 73.200 182.200 74.000 185.400 ;
        RECT 90.800 185.400 93.200 186.200 ;
        RECT 74.800 182.200 75.600 185.000 ;
        RECT 76.400 182.200 77.200 185.000 ;
        RECT 78.000 182.200 78.800 185.000 ;
        RECT 81.200 182.200 82.000 185.000 ;
        RECT 84.400 182.200 85.200 185.000 ;
        RECT 86.000 182.200 86.800 185.000 ;
        RECT 87.600 182.200 88.400 185.000 ;
        RECT 89.200 182.200 90.000 185.000 ;
        RECT 90.800 182.200 91.600 185.400 ;
        RECT 97.200 182.200 98.000 187.400 ;
        RECT 99.000 186.800 99.800 191.200 ;
        RECT 98.800 186.000 99.800 186.800 ;
        RECT 103.400 191.200 104.400 192.000 ;
        RECT 105.000 194.600 107.600 195.200 ;
        RECT 105.000 193.000 105.600 194.600 ;
        RECT 110.000 194.400 110.800 199.800 ;
        RECT 113.200 197.000 114.000 199.800 ;
        RECT 114.800 197.000 115.600 199.800 ;
        RECT 116.400 197.000 117.200 199.800 ;
        RECT 111.400 194.400 115.600 195.200 ;
        RECT 108.200 193.600 110.800 194.400 ;
        RECT 118.000 193.600 118.800 199.800 ;
        RECT 121.200 195.000 122.000 199.800 ;
        RECT 124.400 195.000 125.200 199.800 ;
        RECT 126.000 197.000 126.800 199.800 ;
        RECT 127.600 197.000 128.400 199.800 ;
        RECT 130.800 195.200 131.600 199.800 ;
        RECT 134.000 196.400 134.800 199.800 ;
        RECT 145.200 196.400 146.000 199.800 ;
        RECT 134.000 195.800 135.000 196.400 ;
        RECT 134.400 195.200 135.000 195.800 ;
        RECT 145.000 195.800 146.000 196.400 ;
        RECT 145.000 195.200 145.600 195.800 ;
        RECT 148.400 195.200 149.200 199.800 ;
        RECT 151.600 197.000 152.400 199.800 ;
        RECT 153.200 197.000 154.000 199.800 ;
        RECT 129.600 194.400 133.800 195.200 ;
        RECT 134.400 194.600 136.400 195.200 ;
        RECT 121.200 193.600 123.800 194.400 ;
        RECT 124.400 193.800 130.200 194.400 ;
        RECT 133.200 194.000 133.800 194.400 ;
        RECT 113.200 193.000 114.000 193.200 ;
        RECT 105.000 192.400 114.000 193.000 ;
        RECT 116.400 193.000 117.200 193.200 ;
        RECT 124.400 193.000 125.000 193.800 ;
        RECT 130.800 193.200 132.200 193.800 ;
        RECT 133.200 193.200 134.800 194.000 ;
        RECT 116.400 192.400 125.000 193.000 ;
        RECT 126.000 193.000 132.200 193.200 ;
        RECT 126.000 192.600 131.400 193.000 ;
        RECT 126.000 192.400 126.800 192.600 ;
        RECT 103.400 186.800 104.200 191.200 ;
        RECT 105.000 190.600 105.600 192.400 ;
        RECT 129.000 191.800 130.000 192.000 ;
        RECT 132.400 191.800 133.200 192.400 ;
        RECT 106.200 191.200 133.200 191.800 ;
        RECT 106.200 191.000 107.000 191.200 ;
        RECT 104.800 190.000 105.600 190.600 ;
        RECT 104.800 188.000 105.400 190.000 ;
        RECT 106.000 188.600 109.800 189.400 ;
        RECT 104.800 187.400 106.000 188.000 ;
        RECT 103.400 186.000 104.400 186.800 ;
        RECT 98.800 182.200 99.600 186.000 ;
        RECT 103.600 182.200 104.400 186.000 ;
        RECT 105.200 182.200 106.000 187.400 ;
        RECT 109.000 187.400 109.800 188.600 ;
        RECT 109.000 186.800 110.800 187.400 ;
        RECT 110.000 186.200 110.800 186.800 ;
        RECT 114.800 186.400 115.600 189.200 ;
        RECT 118.000 188.600 121.200 189.400 ;
        RECT 125.000 188.600 127.000 189.400 ;
        RECT 135.600 189.000 136.400 194.600 ;
        RECT 117.600 187.800 118.400 188.000 ;
        RECT 117.600 187.200 122.000 187.800 ;
        RECT 121.200 187.000 122.000 187.200 ;
        RECT 122.800 186.800 123.600 188.400 ;
        RECT 110.000 185.400 112.400 186.200 ;
        RECT 114.800 185.600 115.800 186.400 ;
        RECT 118.800 185.600 120.400 186.400 ;
        RECT 121.200 186.200 122.000 186.400 ;
        RECT 125.000 186.200 125.800 188.600 ;
        RECT 127.600 188.200 136.400 189.000 ;
        RECT 131.000 186.800 134.000 187.600 ;
        RECT 131.000 186.200 131.800 186.800 ;
        RECT 121.200 185.600 125.800 186.200 ;
        RECT 111.600 182.200 112.400 185.400 ;
        RECT 129.200 185.400 131.800 186.200 ;
        RECT 113.200 182.200 114.000 185.000 ;
        RECT 114.800 182.200 115.600 185.000 ;
        RECT 116.400 182.200 117.200 185.000 ;
        RECT 118.000 182.200 118.800 185.000 ;
        RECT 121.200 182.200 122.000 185.000 ;
        RECT 124.400 182.200 125.200 185.000 ;
        RECT 126.000 182.200 126.800 185.000 ;
        RECT 127.600 182.200 128.400 185.000 ;
        RECT 129.200 182.200 130.000 185.400 ;
        RECT 135.600 182.200 136.400 188.200 ;
        RECT 143.600 194.600 145.600 195.200 ;
        RECT 143.600 189.000 144.400 194.600 ;
        RECT 146.200 194.400 150.400 195.200 ;
        RECT 154.800 195.000 155.600 199.800 ;
        RECT 158.000 195.000 158.800 199.800 ;
        RECT 146.200 194.000 146.800 194.400 ;
        RECT 145.200 193.200 146.800 194.000 ;
        RECT 149.800 193.800 155.600 194.400 ;
        RECT 147.800 193.200 149.200 193.800 ;
        RECT 147.800 193.000 154.000 193.200 ;
        RECT 148.600 192.600 154.000 193.000 ;
        RECT 153.200 192.400 154.000 192.600 ;
        RECT 155.000 193.000 155.600 193.800 ;
        RECT 156.200 193.600 158.800 194.400 ;
        RECT 161.200 193.600 162.000 199.800 ;
        RECT 162.800 197.000 163.600 199.800 ;
        RECT 164.400 197.000 165.200 199.800 ;
        RECT 166.000 197.000 166.800 199.800 ;
        RECT 164.400 194.400 168.600 195.200 ;
        RECT 169.200 194.400 170.000 199.800 ;
        RECT 172.400 195.200 173.200 199.800 ;
        RECT 172.400 194.600 175.000 195.200 ;
        RECT 169.200 193.600 171.800 194.400 ;
        RECT 162.800 193.000 163.600 193.200 ;
        RECT 155.000 192.400 163.600 193.000 ;
        RECT 166.000 193.000 166.800 193.200 ;
        RECT 174.400 193.000 175.000 194.600 ;
        RECT 166.000 192.400 175.000 193.000 ;
        RECT 174.400 190.600 175.000 192.400 ;
        RECT 175.600 192.000 176.400 199.800 ;
        RECT 175.600 191.200 176.600 192.000 ;
        RECT 145.000 190.000 168.400 190.600 ;
        RECT 174.400 190.000 175.200 190.600 ;
        RECT 145.000 189.800 145.800 190.000 ;
        RECT 148.400 189.600 149.200 190.000 ;
        RECT 150.000 189.600 150.800 190.000 ;
        RECT 167.600 189.400 168.400 190.000 ;
        RECT 143.600 188.200 152.400 189.000 ;
        RECT 153.000 188.600 155.000 189.400 ;
        RECT 158.800 188.600 162.000 189.400 ;
        RECT 143.600 182.200 144.400 188.200 ;
        RECT 146.000 186.800 149.000 187.600 ;
        RECT 148.200 186.200 149.000 186.800 ;
        RECT 154.200 186.200 155.000 188.600 ;
        RECT 156.400 186.800 157.200 188.400 ;
        RECT 161.600 187.800 162.400 188.000 ;
        RECT 158.000 187.200 162.400 187.800 ;
        RECT 158.000 187.000 158.800 187.200 ;
        RECT 164.400 186.400 165.200 189.200 ;
        RECT 170.200 188.600 174.000 189.400 ;
        RECT 170.200 187.400 171.000 188.600 ;
        RECT 174.600 188.000 175.200 190.000 ;
        RECT 158.000 186.200 158.800 186.400 ;
        RECT 148.200 185.400 150.800 186.200 ;
        RECT 154.200 185.600 158.800 186.200 ;
        RECT 159.600 185.600 161.200 186.400 ;
        RECT 164.200 185.600 165.200 186.400 ;
        RECT 169.200 186.800 171.000 187.400 ;
        RECT 174.000 187.400 175.200 188.000 ;
        RECT 169.200 186.200 170.000 186.800 ;
        RECT 150.000 182.200 150.800 185.400 ;
        RECT 167.600 185.400 170.000 186.200 ;
        RECT 151.600 182.200 152.400 185.000 ;
        RECT 153.200 182.200 154.000 185.000 ;
        RECT 154.800 182.200 155.600 185.000 ;
        RECT 158.000 182.200 158.800 185.000 ;
        RECT 161.200 182.200 162.000 185.000 ;
        RECT 162.800 182.200 163.600 185.000 ;
        RECT 164.400 182.200 165.200 185.000 ;
        RECT 166.000 182.200 166.800 185.000 ;
        RECT 167.600 182.200 168.400 185.400 ;
        RECT 174.000 182.200 174.800 187.400 ;
        RECT 175.800 186.800 176.600 191.200 ;
        RECT 175.600 186.000 176.600 186.800 ;
        RECT 175.600 182.200 176.400 186.000 ;
        RECT 178.800 182.200 179.600 199.800 ;
        RECT 183.600 192.000 184.400 199.800 ;
        RECT 186.800 195.200 187.600 199.800 ;
        RECT 183.400 191.200 184.400 192.000 ;
        RECT 185.000 194.600 187.600 195.200 ;
        RECT 185.000 193.000 185.600 194.600 ;
        RECT 190.000 194.400 190.800 199.800 ;
        RECT 193.200 197.000 194.000 199.800 ;
        RECT 194.800 197.000 195.600 199.800 ;
        RECT 196.400 197.000 197.200 199.800 ;
        RECT 191.400 194.400 195.600 195.200 ;
        RECT 188.200 193.600 190.800 194.400 ;
        RECT 198.000 193.600 198.800 199.800 ;
        RECT 201.200 195.000 202.000 199.800 ;
        RECT 204.400 195.000 205.200 199.800 ;
        RECT 206.000 197.000 206.800 199.800 ;
        RECT 207.600 197.000 208.400 199.800 ;
        RECT 210.800 195.200 211.600 199.800 ;
        RECT 214.000 196.400 214.800 199.800 ;
        RECT 214.000 195.800 215.000 196.400 ;
        RECT 214.400 195.200 215.000 195.800 ;
        RECT 209.600 194.400 213.800 195.200 ;
        RECT 214.400 194.600 216.400 195.200 ;
        RECT 201.200 193.600 203.800 194.400 ;
        RECT 204.400 193.800 210.200 194.400 ;
        RECT 213.200 194.000 213.800 194.400 ;
        RECT 193.200 193.000 194.000 193.200 ;
        RECT 185.000 192.400 194.000 193.000 ;
        RECT 196.400 193.000 197.200 193.200 ;
        RECT 204.400 193.000 205.000 193.800 ;
        RECT 210.800 193.200 212.200 193.800 ;
        RECT 213.200 193.200 214.800 194.000 ;
        RECT 196.400 192.400 205.000 193.000 ;
        RECT 206.000 193.000 212.200 193.200 ;
        RECT 206.000 192.600 211.400 193.000 ;
        RECT 206.000 192.400 206.800 192.600 ;
        RECT 180.400 188.300 181.200 188.400 ;
        RECT 182.000 188.300 182.800 188.400 ;
        RECT 180.400 187.700 182.800 188.300 ;
        RECT 180.400 186.800 181.200 187.700 ;
        RECT 182.000 187.600 182.800 187.700 ;
        RECT 183.400 186.800 184.200 191.200 ;
        RECT 185.000 190.600 185.600 192.400 ;
        RECT 184.800 190.000 185.600 190.600 ;
        RECT 191.600 190.000 215.000 190.600 ;
        RECT 184.800 188.000 185.400 190.000 ;
        RECT 191.600 189.400 192.400 190.000 ;
        RECT 209.200 189.600 210.000 190.000 ;
        RECT 210.800 189.600 211.600 190.000 ;
        RECT 214.200 189.800 215.000 190.000 ;
        RECT 186.000 188.600 189.800 189.400 ;
        RECT 184.800 187.400 186.000 188.000 ;
        RECT 183.400 186.000 184.400 186.800 ;
        RECT 183.600 182.200 184.400 186.000 ;
        RECT 185.200 182.200 186.000 187.400 ;
        RECT 189.000 187.400 189.800 188.600 ;
        RECT 189.000 186.800 190.800 187.400 ;
        RECT 190.000 186.200 190.800 186.800 ;
        RECT 194.800 186.400 195.600 189.200 ;
        RECT 198.000 188.600 201.200 189.400 ;
        RECT 205.000 188.600 207.000 189.400 ;
        RECT 215.600 189.000 216.400 194.600 ;
        RECT 197.600 187.800 198.400 188.000 ;
        RECT 197.600 187.200 202.000 187.800 ;
        RECT 201.200 187.000 202.000 187.200 ;
        RECT 202.800 186.800 203.600 188.400 ;
        RECT 190.000 185.400 192.400 186.200 ;
        RECT 194.800 185.600 195.800 186.400 ;
        RECT 198.800 185.600 200.400 186.400 ;
        RECT 201.200 186.200 202.000 186.400 ;
        RECT 205.000 186.200 205.800 188.600 ;
        RECT 207.600 188.200 216.400 189.000 ;
        RECT 211.000 186.800 214.000 187.600 ;
        RECT 211.000 186.200 211.800 186.800 ;
        RECT 201.200 185.600 205.800 186.200 ;
        RECT 191.600 182.200 192.400 185.400 ;
        RECT 209.200 185.400 211.800 186.200 ;
        RECT 193.200 182.200 194.000 185.000 ;
        RECT 194.800 182.200 195.600 185.000 ;
        RECT 196.400 182.200 197.200 185.000 ;
        RECT 198.000 182.200 198.800 185.000 ;
        RECT 201.200 182.200 202.000 185.000 ;
        RECT 204.400 182.200 205.200 185.000 ;
        RECT 206.000 182.200 206.800 185.000 ;
        RECT 207.600 182.200 208.400 185.000 ;
        RECT 209.200 182.200 210.000 185.400 ;
        RECT 215.600 182.200 216.400 188.200 ;
        RECT 217.200 190.300 218.000 199.800 ;
        RECT 220.400 195.800 221.200 199.800 ;
        RECT 220.600 195.600 221.200 195.800 ;
        RECT 223.600 195.800 224.400 199.800 ;
        RECT 223.600 195.600 224.200 195.800 ;
        RECT 220.600 195.000 224.200 195.600 ;
        RECT 220.600 192.400 221.200 195.000 ;
        RECT 222.000 192.800 222.800 194.400 ;
        RECT 220.400 191.600 221.200 192.400 ;
        RECT 218.800 190.300 219.600 190.400 ;
        RECT 217.200 189.700 219.600 190.300 ;
        RECT 217.200 182.200 218.000 189.700 ;
        RECT 218.800 189.600 219.600 189.700 ;
        RECT 220.600 188.400 221.200 191.600 ;
        RECT 225.200 192.300 226.000 192.400 ;
        RECT 226.800 192.300 227.600 199.800 ;
        RECT 225.200 191.700 227.600 192.300 ;
        RECT 225.200 190.800 226.000 191.700 ;
        RECT 222.800 189.600 224.400 190.400 ;
        RECT 220.600 188.200 222.200 188.400 ;
        RECT 220.600 187.800 222.400 188.200 ;
        RECT 218.800 184.800 219.600 186.400 ;
        RECT 221.600 182.200 222.400 187.800 ;
        RECT 226.800 182.200 227.600 191.700 ;
        RECT 230.000 186.800 230.800 188.400 ;
        RECT 228.400 184.800 229.200 186.400 ;
        RECT 231.600 186.200 232.400 199.800 ;
        RECT 233.200 191.600 234.000 193.200 ;
        RECT 235.400 192.600 236.200 199.800 ;
        RECT 235.400 191.800 237.200 192.600 ;
        RECT 234.800 189.600 235.600 191.200 ;
        RECT 236.400 190.300 237.000 191.800 ;
        RECT 239.600 191.600 240.400 193.200 ;
        RECT 239.700 190.300 240.300 191.600 ;
        RECT 236.400 189.700 240.300 190.300 ;
        RECT 236.400 188.400 237.000 189.700 ;
        RECT 236.400 187.600 237.200 188.400 ;
        RECT 231.600 185.600 233.400 186.200 ;
        RECT 232.600 184.400 233.400 185.600 ;
        RECT 232.600 183.600 234.000 184.400 ;
        RECT 236.400 184.200 237.000 187.600 ;
        RECT 238.000 184.800 238.800 186.400 ;
        RECT 241.200 186.200 242.000 199.800 ;
        RECT 242.800 188.300 243.600 188.400 ;
        RECT 246.000 188.300 246.800 199.800 ;
        RECT 250.200 192.400 251.000 199.800 ;
        RECT 251.600 193.600 252.400 194.400 ;
        RECT 251.800 192.400 252.400 193.600 ;
        RECT 254.000 192.400 254.800 199.800 ;
        RECT 257.200 192.400 258.000 199.800 ;
        RECT 250.200 191.800 251.200 192.400 ;
        RECT 251.800 191.800 253.200 192.400 ;
        RECT 254.000 191.800 258.000 192.400 ;
        RECT 258.800 191.800 259.600 199.800 ;
        RECT 268.400 192.000 269.200 199.800 ;
        RECT 271.600 195.200 272.400 199.800 ;
        RECT 249.200 188.800 250.000 190.400 ;
        RECT 250.600 188.400 251.200 191.800 ;
        RECT 252.400 191.600 253.200 191.800 ;
        RECT 254.800 190.400 255.600 190.800 ;
        RECT 258.800 190.400 259.400 191.800 ;
        RECT 268.200 191.200 269.200 192.000 ;
        RECT 269.800 194.600 272.400 195.200 ;
        RECT 269.800 193.000 270.400 194.600 ;
        RECT 274.800 194.400 275.600 199.800 ;
        RECT 278.000 197.000 278.800 199.800 ;
        RECT 279.600 197.000 280.400 199.800 ;
        RECT 281.200 197.000 282.000 199.800 ;
        RECT 276.200 194.400 280.400 195.200 ;
        RECT 273.000 193.600 275.600 194.400 ;
        RECT 282.800 193.600 283.600 199.800 ;
        RECT 286.000 195.000 286.800 199.800 ;
        RECT 289.200 195.000 290.000 199.800 ;
        RECT 290.800 197.000 291.600 199.800 ;
        RECT 292.400 197.000 293.200 199.800 ;
        RECT 295.600 195.200 296.400 199.800 ;
        RECT 298.800 196.400 299.600 199.800 ;
        RECT 298.800 195.800 299.800 196.400 ;
        RECT 299.200 195.200 299.800 195.800 ;
        RECT 294.400 194.400 298.600 195.200 ;
        RECT 299.200 194.600 301.200 195.200 ;
        RECT 286.000 193.600 288.600 194.400 ;
        RECT 289.200 193.800 295.000 194.400 ;
        RECT 298.000 194.000 298.600 194.400 ;
        RECT 278.000 193.000 278.800 193.200 ;
        RECT 269.800 192.400 278.800 193.000 ;
        RECT 281.200 193.000 282.000 193.200 ;
        RECT 289.200 193.000 289.800 193.800 ;
        RECT 295.600 193.200 297.000 193.800 ;
        RECT 298.000 193.200 299.600 194.000 ;
        RECT 281.200 192.400 289.800 193.000 ;
        RECT 290.800 193.000 297.000 193.200 ;
        RECT 290.800 192.600 296.200 193.000 ;
        RECT 290.800 192.400 291.600 192.600 ;
        RECT 254.000 189.800 255.600 190.400 ;
        RECT 257.200 189.800 259.600 190.400 ;
        RECT 254.000 189.600 254.800 189.800 ;
        RECT 247.600 188.300 248.400 188.400 ;
        RECT 242.800 187.700 245.100 188.300 ;
        RECT 242.800 186.800 243.600 187.700 ;
        RECT 244.500 186.400 245.100 187.700 ;
        RECT 246.000 188.200 248.400 188.300 ;
        RECT 250.600 188.300 253.200 188.400 ;
        RECT 255.600 188.300 256.400 189.200 ;
        RECT 246.000 187.700 249.200 188.200 ;
        RECT 240.200 185.600 242.000 186.200 ;
        RECT 240.200 184.400 241.000 185.600 ;
        RECT 244.400 184.800 245.200 186.400 ;
        RECT 232.600 182.200 233.400 183.600 ;
        RECT 236.400 182.200 237.200 184.200 ;
        RECT 239.600 183.600 241.000 184.400 ;
        RECT 240.200 182.200 241.000 183.600 ;
        RECT 246.000 182.200 246.800 187.700 ;
        RECT 247.600 187.600 249.200 187.700 ;
        RECT 250.600 187.700 256.400 188.300 ;
        RECT 250.600 187.600 253.200 187.700 ;
        RECT 255.600 187.600 256.400 187.700 ;
        RECT 257.200 188.300 257.800 189.800 ;
        RECT 258.800 189.600 259.600 189.800 ;
        RECT 266.800 188.300 267.600 188.400 ;
        RECT 257.200 187.700 267.600 188.300 ;
        RECT 248.400 187.200 249.200 187.600 ;
        RECT 247.800 186.200 251.400 186.600 ;
        RECT 252.400 186.200 253.000 187.600 ;
        RECT 257.200 186.200 257.800 187.700 ;
        RECT 266.800 187.600 267.600 187.700 ;
        RECT 268.200 186.800 269.000 191.200 ;
        RECT 269.800 190.600 270.400 192.400 ;
        RECT 269.600 190.000 270.400 190.600 ;
        RECT 276.400 190.000 299.800 190.600 ;
        RECT 269.600 188.000 270.200 190.000 ;
        RECT 276.400 189.400 277.200 190.000 ;
        RECT 294.000 189.600 294.800 190.000 ;
        RECT 297.200 189.600 298.000 190.000 ;
        RECT 299.000 189.800 299.800 190.000 ;
        RECT 270.800 188.600 274.600 189.400 ;
        RECT 269.600 187.400 270.800 188.000 ;
        RECT 258.800 186.300 259.600 186.400 ;
        RECT 263.600 186.300 264.400 186.400 ;
        RECT 247.600 186.000 251.600 186.200 ;
        RECT 247.600 182.200 248.400 186.000 ;
        RECT 250.800 182.200 251.600 186.000 ;
        RECT 252.400 182.200 253.200 186.200 ;
        RECT 257.200 182.200 258.000 186.200 ;
        RECT 258.800 185.700 264.400 186.300 ;
        RECT 268.200 186.000 269.200 186.800 ;
        RECT 258.800 185.600 259.600 185.700 ;
        RECT 263.600 185.600 264.400 185.700 ;
        RECT 258.600 184.800 259.400 185.600 ;
        RECT 268.400 182.200 269.200 186.000 ;
        RECT 270.000 182.200 270.800 187.400 ;
        RECT 273.800 187.400 274.600 188.600 ;
        RECT 273.800 186.800 275.600 187.400 ;
        RECT 274.800 186.200 275.600 186.800 ;
        RECT 279.600 186.400 280.400 189.200 ;
        RECT 282.800 188.600 286.000 189.400 ;
        RECT 289.800 188.600 291.800 189.400 ;
        RECT 300.400 189.000 301.200 194.600 ;
        RECT 303.600 192.000 304.400 199.800 ;
        RECT 306.800 195.200 307.600 199.800 ;
        RECT 282.400 187.800 283.200 188.000 ;
        RECT 282.400 187.200 286.800 187.800 ;
        RECT 286.000 187.000 286.800 187.200 ;
        RECT 287.600 186.800 288.400 188.400 ;
        RECT 274.800 185.400 277.200 186.200 ;
        RECT 279.600 185.600 280.600 186.400 ;
        RECT 283.600 185.600 285.200 186.400 ;
        RECT 286.000 186.200 286.800 186.400 ;
        RECT 289.800 186.200 290.600 188.600 ;
        RECT 292.400 188.200 301.200 189.000 ;
        RECT 295.800 186.800 298.800 187.600 ;
        RECT 295.800 186.200 296.600 186.800 ;
        RECT 286.000 185.600 290.600 186.200 ;
        RECT 276.400 182.200 277.200 185.400 ;
        RECT 294.000 185.400 296.600 186.200 ;
        RECT 278.000 182.200 278.800 185.000 ;
        RECT 279.600 182.200 280.400 185.000 ;
        RECT 281.200 182.200 282.000 185.000 ;
        RECT 282.800 182.200 283.600 185.000 ;
        RECT 286.000 182.200 286.800 185.000 ;
        RECT 289.200 182.200 290.000 185.000 ;
        RECT 290.800 182.200 291.600 185.000 ;
        RECT 292.400 182.200 293.200 185.000 ;
        RECT 294.000 182.200 294.800 185.400 ;
        RECT 300.400 182.200 301.200 188.200 ;
        RECT 303.400 191.200 304.400 192.000 ;
        RECT 305.000 194.600 307.600 195.200 ;
        RECT 305.000 193.000 305.600 194.600 ;
        RECT 310.000 194.400 310.800 199.800 ;
        RECT 313.200 197.000 314.000 199.800 ;
        RECT 314.800 197.000 315.600 199.800 ;
        RECT 316.400 197.000 317.200 199.800 ;
        RECT 311.400 194.400 315.600 195.200 ;
        RECT 308.200 193.600 310.800 194.400 ;
        RECT 318.000 193.600 318.800 199.800 ;
        RECT 321.200 195.000 322.000 199.800 ;
        RECT 324.400 195.000 325.200 199.800 ;
        RECT 326.000 197.000 326.800 199.800 ;
        RECT 327.600 197.000 328.400 199.800 ;
        RECT 330.800 195.200 331.600 199.800 ;
        RECT 334.000 196.400 334.800 199.800 ;
        RECT 334.000 195.800 335.000 196.400 ;
        RECT 334.400 195.200 335.000 195.800 ;
        RECT 329.600 194.400 333.800 195.200 ;
        RECT 334.400 194.600 336.400 195.200 ;
        RECT 321.200 193.600 323.800 194.400 ;
        RECT 324.400 193.800 330.200 194.400 ;
        RECT 333.200 194.000 333.800 194.400 ;
        RECT 313.200 193.000 314.000 193.200 ;
        RECT 305.000 192.400 314.000 193.000 ;
        RECT 316.400 193.000 317.200 193.200 ;
        RECT 324.400 193.000 325.000 193.800 ;
        RECT 330.800 193.200 332.200 193.800 ;
        RECT 333.200 193.200 334.800 194.000 ;
        RECT 316.400 192.400 325.000 193.000 ;
        RECT 326.000 193.000 332.200 193.200 ;
        RECT 326.000 192.600 331.400 193.000 ;
        RECT 326.000 192.400 326.800 192.600 ;
        RECT 303.400 186.800 304.200 191.200 ;
        RECT 305.000 190.600 305.600 192.400 ;
        RECT 329.000 191.800 329.800 192.000 ;
        RECT 332.400 191.800 333.200 192.400 ;
        RECT 306.200 191.200 333.200 191.800 ;
        RECT 306.200 191.000 307.000 191.200 ;
        RECT 304.800 190.000 305.600 190.600 ;
        RECT 304.800 188.000 305.400 190.000 ;
        RECT 306.000 188.600 309.800 189.400 ;
        RECT 304.800 187.400 306.000 188.000 ;
        RECT 303.400 186.000 304.400 186.800 ;
        RECT 303.600 182.200 304.400 186.000 ;
        RECT 305.200 182.200 306.000 187.400 ;
        RECT 309.000 187.400 309.800 188.600 ;
        RECT 309.000 186.800 310.800 187.400 ;
        RECT 310.000 186.200 310.800 186.800 ;
        RECT 314.800 186.400 315.600 189.200 ;
        RECT 318.000 188.600 321.200 189.400 ;
        RECT 325.000 188.600 327.000 189.400 ;
        RECT 335.600 189.000 336.400 194.600 ;
        RECT 317.600 187.800 318.400 188.000 ;
        RECT 317.600 187.200 322.000 187.800 ;
        RECT 321.200 187.000 322.000 187.200 ;
        RECT 322.800 186.800 323.600 188.400 ;
        RECT 310.000 185.400 312.400 186.200 ;
        RECT 314.800 185.600 315.800 186.400 ;
        RECT 318.800 185.600 320.400 186.400 ;
        RECT 321.200 186.200 322.000 186.400 ;
        RECT 325.000 186.200 325.800 188.600 ;
        RECT 327.600 188.200 336.400 189.000 ;
        RECT 331.000 186.800 334.000 187.600 ;
        RECT 331.000 186.200 331.800 186.800 ;
        RECT 321.200 185.600 325.800 186.200 ;
        RECT 311.600 182.200 312.400 185.400 ;
        RECT 329.200 185.400 331.800 186.200 ;
        RECT 313.200 182.200 314.000 185.000 ;
        RECT 314.800 182.200 315.600 185.000 ;
        RECT 316.400 182.200 317.200 185.000 ;
        RECT 318.000 182.200 318.800 185.000 ;
        RECT 321.200 182.200 322.000 185.000 ;
        RECT 324.400 182.200 325.200 185.000 ;
        RECT 326.000 182.200 326.800 185.000 ;
        RECT 327.600 182.200 328.400 185.000 ;
        RECT 329.200 182.200 330.000 185.400 ;
        RECT 335.600 182.200 336.400 188.200 ;
        RECT 338.800 188.300 339.600 199.800 ;
        RECT 343.000 192.400 343.800 199.800 ;
        RECT 348.400 196.400 349.200 199.800 ;
        RECT 348.200 195.800 349.200 196.400 ;
        RECT 348.200 195.200 348.800 195.800 ;
        RECT 351.600 195.200 352.400 199.800 ;
        RECT 354.800 197.000 355.600 199.800 ;
        RECT 356.400 197.000 357.200 199.800 ;
        RECT 346.800 194.600 348.800 195.200 ;
        RECT 344.400 193.600 345.200 194.400 ;
        RECT 344.600 192.400 345.200 193.600 ;
        RECT 343.000 191.800 344.000 192.400 ;
        RECT 344.600 191.800 346.000 192.400 ;
        RECT 342.000 188.800 342.800 190.400 ;
        RECT 343.400 188.400 344.000 191.800 ;
        RECT 345.200 191.600 346.000 191.800 ;
        RECT 346.800 189.000 347.600 194.600 ;
        RECT 349.400 194.400 353.600 195.200 ;
        RECT 358.000 195.000 358.800 199.800 ;
        RECT 361.200 195.000 362.000 199.800 ;
        RECT 349.400 194.000 350.000 194.400 ;
        RECT 348.400 193.200 350.000 194.000 ;
        RECT 353.000 193.800 358.800 194.400 ;
        RECT 351.000 193.200 352.400 193.800 ;
        RECT 351.000 193.000 357.200 193.200 ;
        RECT 351.800 192.600 357.200 193.000 ;
        RECT 356.400 192.400 357.200 192.600 ;
        RECT 358.200 193.000 358.800 193.800 ;
        RECT 359.400 193.600 362.000 194.400 ;
        RECT 364.400 193.600 365.200 199.800 ;
        RECT 366.000 197.000 366.800 199.800 ;
        RECT 367.600 197.000 368.400 199.800 ;
        RECT 369.200 197.000 370.000 199.800 ;
        RECT 367.600 194.400 371.800 195.200 ;
        RECT 372.400 194.400 373.200 199.800 ;
        RECT 375.600 195.200 376.400 199.800 ;
        RECT 375.600 194.600 378.200 195.200 ;
        RECT 372.400 193.600 375.000 194.400 ;
        RECT 366.000 193.000 366.800 193.200 ;
        RECT 358.200 192.400 366.800 193.000 ;
        RECT 369.200 193.000 370.000 193.200 ;
        RECT 377.600 193.000 378.200 194.600 ;
        RECT 369.200 192.400 378.200 193.000 ;
        RECT 350.000 191.800 350.800 192.400 ;
        RECT 353.200 191.800 354.200 192.000 ;
        RECT 350.000 191.200 377.000 191.800 ;
        RECT 376.200 191.000 377.000 191.200 ;
        RECT 377.600 190.600 378.200 192.400 ;
        RECT 378.800 192.000 379.600 199.800 ;
        RECT 382.800 193.600 383.600 194.400 ;
        RECT 382.800 192.400 383.400 193.600 ;
        RECT 384.200 192.400 385.000 199.800 ;
        RECT 390.000 195.800 390.800 199.800 ;
        RECT 390.200 195.600 390.800 195.800 ;
        RECT 393.200 195.800 394.000 199.800 ;
        RECT 393.200 195.600 393.800 195.800 ;
        RECT 390.200 195.000 393.800 195.600 ;
        RECT 391.600 192.800 392.400 194.400 ;
        RECT 393.200 192.400 393.800 195.000 ;
        RECT 380.400 192.300 381.200 192.400 ;
        RECT 382.000 192.300 383.400 192.400 ;
        RECT 378.800 191.200 379.800 192.000 ;
        RECT 380.400 191.800 383.400 192.300 ;
        RECT 384.000 191.800 385.000 192.400 ;
        RECT 380.400 191.700 382.800 191.800 ;
        RECT 380.400 191.600 381.200 191.700 ;
        RECT 382.000 191.600 382.800 191.700 ;
        RECT 377.600 190.000 378.400 190.600 ;
        RECT 340.400 188.300 341.200 188.400 ;
        RECT 338.800 188.200 341.200 188.300 ;
        RECT 338.800 187.700 342.000 188.200 ;
        RECT 337.200 184.800 338.000 186.400 ;
        RECT 338.800 182.200 339.600 187.700 ;
        RECT 340.400 187.600 342.000 187.700 ;
        RECT 343.400 187.600 346.000 188.400 ;
        RECT 346.800 188.200 355.600 189.000 ;
        RECT 356.200 188.600 358.200 189.400 ;
        RECT 362.000 188.600 365.200 189.400 ;
        RECT 341.200 187.200 342.000 187.600 ;
        RECT 340.600 186.200 344.200 186.600 ;
        RECT 345.200 186.200 345.800 187.600 ;
        RECT 340.400 186.000 344.400 186.200 ;
        RECT 340.400 182.200 341.200 186.000 ;
        RECT 343.600 182.200 344.400 186.000 ;
        RECT 345.200 182.200 346.000 186.200 ;
        RECT 346.800 182.200 347.600 188.200 ;
        RECT 349.200 186.800 352.200 187.600 ;
        RECT 351.400 186.200 352.200 186.800 ;
        RECT 357.400 186.200 358.200 188.600 ;
        RECT 359.600 186.800 360.400 188.400 ;
        RECT 364.800 187.800 365.600 188.000 ;
        RECT 361.200 187.200 365.600 187.800 ;
        RECT 361.200 187.000 362.000 187.200 ;
        RECT 367.600 186.400 368.400 189.200 ;
        RECT 373.400 188.600 377.200 189.400 ;
        RECT 373.400 187.400 374.200 188.600 ;
        RECT 377.800 188.000 378.400 190.000 ;
        RECT 361.200 186.200 362.000 186.400 ;
        RECT 351.400 185.400 354.000 186.200 ;
        RECT 357.400 185.600 362.000 186.200 ;
        RECT 362.800 185.600 364.400 186.400 ;
        RECT 367.400 185.600 368.400 186.400 ;
        RECT 372.400 186.800 374.200 187.400 ;
        RECT 377.200 187.400 378.400 188.000 ;
        RECT 372.400 186.200 373.200 186.800 ;
        RECT 353.200 182.200 354.000 185.400 ;
        RECT 370.800 185.400 373.200 186.200 ;
        RECT 354.800 182.200 355.600 185.000 ;
        RECT 356.400 182.200 357.200 185.000 ;
        RECT 358.000 182.200 358.800 185.000 ;
        RECT 361.200 182.200 362.000 185.000 ;
        RECT 364.400 182.200 365.200 185.000 ;
        RECT 366.000 182.200 366.800 185.000 ;
        RECT 367.600 182.200 368.400 185.000 ;
        RECT 369.200 182.200 370.000 185.000 ;
        RECT 370.800 182.200 371.600 185.400 ;
        RECT 377.200 182.200 378.000 187.400 ;
        RECT 379.000 186.800 379.800 191.200 ;
        RECT 384.000 188.400 384.600 191.800 ;
        RECT 388.400 190.800 389.200 192.400 ;
        RECT 393.200 191.600 394.000 192.400 ;
        RECT 394.800 191.600 395.600 193.200 ;
        RECT 385.200 188.800 386.000 190.400 ;
        RECT 390.000 189.600 391.600 190.400 ;
        RECT 393.200 188.400 393.800 191.600 ;
        RECT 382.000 187.600 384.600 188.400 ;
        RECT 386.800 188.200 387.600 188.400 ;
        RECT 392.200 188.200 393.800 188.400 ;
        RECT 386.000 187.600 387.600 188.200 ;
        RECT 392.000 187.800 393.800 188.200 ;
        RECT 378.800 186.000 379.800 186.800 ;
        RECT 380.400 186.300 381.200 186.400 ;
        RECT 382.200 186.300 382.800 187.600 ;
        RECT 386.000 187.200 386.800 187.600 ;
        RECT 378.800 182.200 379.600 186.000 ;
        RECT 380.400 185.700 382.800 186.300 ;
        RECT 383.800 186.200 387.400 186.600 ;
        RECT 380.400 185.600 381.200 185.700 ;
        RECT 382.000 182.200 382.800 185.700 ;
        RECT 383.600 186.000 387.600 186.200 ;
        RECT 383.600 182.200 384.400 186.000 ;
        RECT 386.800 182.200 387.600 186.000 ;
        RECT 392.000 182.200 392.800 187.800 ;
        RECT 396.400 186.400 397.200 199.800 ;
        RECT 402.200 192.400 403.000 199.800 ;
        RECT 403.600 193.600 404.400 194.400 ;
        RECT 403.800 192.400 404.400 193.600 ;
        RECT 402.200 191.800 403.200 192.400 ;
        RECT 403.800 191.800 405.200 192.400 ;
        RECT 401.200 188.800 402.000 190.400 ;
        RECT 402.600 188.400 403.200 191.800 ;
        RECT 404.400 191.600 405.200 191.800 ;
        RECT 398.000 186.800 398.800 188.400 ;
        RECT 399.600 188.200 400.400 188.400 ;
        RECT 399.600 187.600 401.200 188.200 ;
        RECT 402.600 187.600 405.200 188.400 ;
        RECT 400.400 187.200 401.200 187.600 ;
        RECT 394.800 185.600 397.200 186.400 ;
        RECT 399.800 186.200 403.400 186.600 ;
        RECT 404.400 186.200 405.000 187.600 ;
        RECT 399.600 186.000 403.600 186.200 ;
        RECT 395.400 182.200 396.200 185.600 ;
        RECT 399.600 182.200 400.400 186.000 ;
        RECT 402.800 182.200 403.600 186.000 ;
        RECT 404.400 182.200 405.200 186.200 ;
        RECT 407.600 182.200 408.400 199.800 ;
        RECT 410.800 195.800 411.600 199.800 ;
        RECT 411.000 195.600 411.600 195.800 ;
        RECT 414.000 195.800 414.800 199.800 ;
        RECT 414.000 195.600 414.600 195.800 ;
        RECT 411.000 195.000 414.600 195.600 ;
        RECT 412.400 192.800 413.200 194.400 ;
        RECT 414.000 192.400 414.600 195.000 ;
        RECT 409.200 190.800 410.000 192.400 ;
        RECT 414.000 191.600 414.800 192.400 ;
        RECT 410.800 189.600 412.400 190.400 ;
        RECT 414.000 188.400 414.600 191.600 ;
        RECT 413.000 188.200 414.600 188.400 ;
        RECT 412.800 187.800 414.600 188.200 ;
        RECT 412.800 182.200 413.600 187.800 ;
        RECT 415.600 182.200 416.400 199.800 ;
        RECT 421.400 198.400 422.200 199.800 ;
        RECT 420.400 197.600 422.200 198.400 ;
        RECT 421.400 192.400 422.200 197.600 ;
        RECT 422.800 194.300 423.600 194.400 ;
        RECT 430.000 194.300 430.800 194.400 ;
        RECT 422.800 193.700 430.800 194.300 ;
        RECT 422.800 193.600 423.600 193.700 ;
        RECT 430.000 193.600 430.800 193.700 ;
        RECT 423.000 192.400 423.600 193.600 ;
        RECT 421.400 191.800 422.400 192.400 ;
        RECT 423.000 191.800 424.400 192.400 ;
        RECT 417.200 190.300 418.000 190.400 ;
        RECT 420.400 190.300 421.200 190.400 ;
        RECT 417.200 189.700 421.200 190.300 ;
        RECT 417.200 189.600 418.000 189.700 ;
        RECT 420.400 188.800 421.200 189.700 ;
        RECT 421.800 188.400 422.400 191.800 ;
        RECT 423.600 191.600 424.400 191.800 ;
        RECT 431.600 192.300 432.400 199.800 ;
        RECT 434.800 195.000 435.600 199.000 ;
        RECT 433.200 192.300 434.000 192.400 ;
        RECT 431.600 191.700 434.000 192.300 ;
        RECT 418.800 188.200 419.600 188.400 ;
        RECT 418.800 187.600 420.400 188.200 ;
        RECT 421.800 187.600 424.400 188.400 ;
        RECT 419.600 187.200 420.400 187.600 ;
        RECT 417.200 184.800 418.000 186.400 ;
        RECT 419.000 186.200 422.600 186.600 ;
        RECT 423.600 186.200 424.200 187.600 ;
        RECT 418.800 186.000 422.800 186.200 ;
        RECT 418.800 182.200 419.600 186.000 ;
        RECT 422.000 182.200 422.800 186.000 ;
        RECT 423.600 182.200 424.400 186.200 ;
        RECT 431.600 182.200 432.400 191.700 ;
        RECT 433.200 191.600 434.000 191.700 ;
        RECT 434.800 191.600 435.400 195.000 ;
        RECT 439.000 192.800 439.800 199.800 ;
        RECT 444.400 195.800 445.200 199.800 ;
        RECT 444.600 195.600 445.200 195.800 ;
        RECT 447.600 195.800 448.400 199.800 ;
        RECT 447.600 195.600 448.200 195.800 ;
        RECT 444.600 195.000 448.200 195.600 ;
        RECT 439.000 192.200 440.600 192.800 ;
        RECT 444.600 192.400 445.200 195.000 ;
        RECT 446.000 192.800 446.800 194.400 ;
        RECT 434.800 191.000 438.600 191.600 ;
        RECT 434.800 188.800 435.600 190.400 ;
        RECT 436.400 188.800 437.200 190.400 ;
        RECT 438.000 189.000 438.600 191.000 ;
        RECT 438.000 188.200 439.400 189.000 ;
        RECT 440.000 188.400 440.600 192.200 ;
        RECT 444.400 191.600 445.200 192.400 ;
        RECT 450.800 192.400 451.600 199.800 ;
        RECT 450.800 191.800 453.000 192.400 ;
        RECT 454.000 191.800 454.800 199.800 ;
        RECT 455.600 195.800 456.400 199.800 ;
        RECT 455.800 195.600 456.400 195.800 ;
        RECT 458.800 195.800 459.600 199.800 ;
        RECT 464.200 198.400 465.000 199.800 ;
        RECT 464.200 197.600 466.000 198.400 ;
        RECT 458.800 195.600 459.400 195.800 ;
        RECT 455.800 195.000 459.400 195.600 ;
        RECT 455.800 192.400 456.400 195.000 ;
        RECT 457.200 194.300 458.000 194.400 ;
        RECT 460.400 194.300 461.200 194.400 ;
        RECT 457.200 193.700 461.200 194.300 ;
        RECT 457.200 192.800 458.000 193.700 ;
        RECT 460.400 193.600 461.200 193.700 ;
        RECT 462.800 193.600 463.600 194.400 ;
        RECT 462.800 192.400 463.400 193.600 ;
        RECT 464.200 192.400 465.000 197.600 ;
        RECT 441.200 189.600 442.000 191.200 ;
        RECT 444.600 188.400 445.200 191.600 ;
        RECT 452.400 191.200 453.000 191.800 ;
        RECT 452.400 190.400 453.600 191.200 ;
        RECT 446.800 189.600 448.400 190.400 ;
        RECT 438.000 187.800 439.000 188.200 ;
        RECT 434.800 187.200 439.000 187.800 ;
        RECT 440.000 187.600 442.000 188.400 ;
        RECT 444.600 188.200 446.200 188.400 ;
        RECT 444.600 187.800 446.400 188.200 ;
        RECT 433.200 184.800 434.000 186.400 ;
        RECT 434.800 185.000 435.400 187.200 ;
        RECT 440.000 187.000 440.600 187.600 ;
        RECT 439.800 186.600 440.600 187.000 ;
        RECT 439.000 186.000 440.600 186.600 ;
        RECT 434.800 183.000 435.600 185.000 ;
        RECT 439.000 184.400 439.800 186.000 ;
        RECT 439.000 183.600 440.400 184.400 ;
        RECT 439.000 183.000 439.800 183.600 ;
        RECT 445.600 182.200 446.400 187.800 ;
        RECT 452.400 187.400 453.000 190.400 ;
        RECT 454.200 189.600 454.800 191.800 ;
        RECT 455.600 191.600 456.400 192.400 ;
        RECT 450.800 186.800 453.000 187.400 ;
        RECT 450.800 182.200 451.600 186.800 ;
        RECT 454.000 182.200 454.800 189.600 ;
        RECT 455.800 188.400 456.400 191.600 ;
        RECT 460.400 190.800 461.200 192.400 ;
        RECT 462.000 191.800 463.400 192.400 ;
        RECT 464.000 191.800 465.000 192.400 ;
        RECT 470.000 192.000 470.800 199.800 ;
        RECT 473.200 195.200 474.000 199.800 ;
        RECT 462.000 191.600 462.800 191.800 ;
        RECT 458.000 189.600 459.600 190.400 ;
        RECT 464.000 188.400 464.600 191.800 ;
        RECT 469.800 191.200 470.800 192.000 ;
        RECT 471.400 194.600 474.000 195.200 ;
        RECT 471.400 193.000 472.000 194.600 ;
        RECT 476.400 194.400 477.200 199.800 ;
        RECT 479.600 197.000 480.400 199.800 ;
        RECT 481.200 197.000 482.000 199.800 ;
        RECT 482.800 197.000 483.600 199.800 ;
        RECT 477.800 194.400 482.000 195.200 ;
        RECT 474.600 193.600 477.200 194.400 ;
        RECT 484.400 193.600 485.200 199.800 ;
        RECT 487.600 195.000 488.400 199.800 ;
        RECT 490.800 195.000 491.600 199.800 ;
        RECT 492.400 197.000 493.200 199.800 ;
        RECT 494.000 197.000 494.800 199.800 ;
        RECT 497.200 195.200 498.000 199.800 ;
        RECT 500.400 196.400 501.200 199.800 ;
        RECT 506.200 198.400 508.200 199.800 ;
        RECT 506.200 197.600 509.200 198.400 ;
        RECT 500.400 195.800 501.400 196.400 ;
        RECT 500.800 195.200 501.400 195.800 ;
        RECT 496.000 194.400 500.200 195.200 ;
        RECT 500.800 194.600 502.800 195.200 ;
        RECT 487.600 193.600 490.200 194.400 ;
        RECT 490.800 193.800 496.600 194.400 ;
        RECT 499.600 194.000 500.200 194.400 ;
        RECT 479.600 193.000 480.400 193.200 ;
        RECT 471.400 192.400 480.400 193.000 ;
        RECT 482.800 193.000 483.600 193.200 ;
        RECT 490.800 193.000 491.400 193.800 ;
        RECT 497.200 193.200 498.600 193.800 ;
        RECT 499.600 193.200 501.200 194.000 ;
        RECT 482.800 192.400 491.400 193.000 ;
        RECT 492.400 193.000 498.600 193.200 ;
        RECT 492.400 192.600 497.800 193.000 ;
        RECT 492.400 192.400 493.200 192.600 ;
        RECT 465.200 188.800 466.000 190.400 ;
        RECT 455.800 188.300 457.400 188.400 ;
        RECT 458.800 188.300 459.600 188.400 ;
        RECT 455.800 187.800 459.600 188.300 ;
        RECT 456.800 187.700 459.600 187.800 ;
        RECT 456.800 187.600 458.000 187.700 ;
        RECT 458.800 187.600 459.600 187.700 ;
        RECT 462.000 187.600 464.600 188.400 ;
        RECT 466.800 188.200 467.600 188.400 ;
        RECT 466.000 187.600 467.600 188.200 ;
        RECT 456.800 182.200 457.600 187.600 ;
        RECT 462.200 186.200 462.800 187.600 ;
        RECT 466.000 187.200 466.800 187.600 ;
        RECT 469.800 186.800 470.600 191.200 ;
        RECT 471.400 190.600 472.000 192.400 ;
        RECT 471.200 190.000 472.000 190.600 ;
        RECT 478.000 190.000 501.400 190.600 ;
        RECT 471.200 188.000 471.800 190.000 ;
        RECT 478.000 189.400 478.800 190.000 ;
        RECT 495.600 189.600 496.400 190.000 ;
        RECT 497.200 189.600 498.000 190.000 ;
        RECT 500.600 189.800 501.400 190.000 ;
        RECT 472.400 188.600 476.200 189.400 ;
        RECT 471.200 187.400 472.400 188.000 ;
        RECT 463.800 186.200 467.400 186.600 ;
        RECT 462.000 182.200 462.800 186.200 ;
        RECT 463.600 186.000 467.600 186.200 ;
        RECT 469.800 186.000 470.800 186.800 ;
        RECT 463.600 182.200 464.400 186.000 ;
        RECT 466.800 182.200 467.600 186.000 ;
        RECT 470.000 182.200 470.800 186.000 ;
        RECT 471.600 182.200 472.400 187.400 ;
        RECT 475.400 187.400 476.200 188.600 ;
        RECT 475.400 186.800 477.200 187.400 ;
        RECT 476.400 186.200 477.200 186.800 ;
        RECT 481.200 186.400 482.000 189.200 ;
        RECT 484.400 188.600 487.600 189.400 ;
        RECT 491.400 188.600 493.400 189.400 ;
        RECT 502.000 189.000 502.800 194.600 ;
        RECT 506.200 191.800 508.200 197.600 ;
        RECT 511.600 195.000 512.400 199.000 ;
        RECT 515.800 198.400 516.600 199.800 ;
        RECT 514.800 197.600 516.600 198.400 ;
        RECT 484.000 187.800 484.800 188.000 ;
        RECT 484.000 187.200 488.400 187.800 ;
        RECT 487.600 187.000 488.400 187.200 ;
        RECT 489.200 186.800 490.000 188.400 ;
        RECT 476.400 185.400 478.800 186.200 ;
        RECT 481.200 185.600 482.200 186.400 ;
        RECT 485.200 185.600 486.800 186.400 ;
        RECT 487.600 186.200 488.400 186.400 ;
        RECT 491.400 186.200 492.200 188.600 ;
        RECT 494.000 188.200 502.800 189.000 ;
        RECT 505.200 188.800 506.000 190.400 ;
        RECT 506.800 188.400 507.400 191.800 ;
        RECT 511.600 191.600 512.200 195.000 ;
        RECT 515.800 192.800 516.600 197.600 ;
        RECT 515.800 192.200 517.400 192.800 ;
        RECT 511.600 191.000 515.400 191.600 ;
        RECT 508.400 188.800 509.200 190.400 ;
        RECT 497.400 186.800 500.400 187.600 ;
        RECT 497.400 186.200 498.200 186.800 ;
        RECT 487.600 185.600 492.200 186.200 ;
        RECT 478.000 182.200 478.800 185.400 ;
        RECT 495.600 185.400 498.200 186.200 ;
        RECT 479.600 182.200 480.400 185.000 ;
        RECT 481.200 182.200 482.000 185.000 ;
        RECT 482.800 182.200 483.600 185.000 ;
        RECT 484.400 182.200 485.200 185.000 ;
        RECT 487.600 182.200 488.400 185.000 ;
        RECT 490.800 182.200 491.600 185.000 ;
        RECT 492.400 182.200 493.200 185.000 ;
        RECT 494.000 182.200 494.800 185.000 ;
        RECT 495.600 182.200 496.400 185.400 ;
        RECT 502.000 182.200 502.800 188.200 ;
        RECT 503.600 188.200 504.400 188.400 ;
        RECT 506.800 188.200 507.600 188.400 ;
        RECT 503.600 187.600 505.200 188.200 ;
        RECT 506.800 187.600 509.200 188.200 ;
        RECT 510.000 187.600 510.800 189.200 ;
        RECT 511.600 188.800 512.400 190.400 ;
        RECT 513.200 188.800 514.000 190.400 ;
        RECT 514.800 189.000 515.400 191.000 ;
        RECT 514.800 188.200 516.200 189.000 ;
        RECT 516.800 188.400 517.400 192.200 ;
        RECT 521.200 191.400 522.000 199.800 ;
        RECT 525.600 196.400 526.400 199.800 ;
        RECT 524.400 195.800 526.400 196.400 ;
        RECT 530.000 195.800 530.800 199.800 ;
        RECT 534.200 195.800 535.400 199.800 ;
        RECT 524.400 195.000 525.200 195.800 ;
        RECT 530.000 195.200 530.600 195.800 ;
        RECT 527.800 194.600 531.400 195.200 ;
        RECT 534.000 195.000 534.800 195.800 ;
        RECT 527.800 194.400 528.600 194.600 ;
        RECT 530.600 194.400 531.400 194.600 ;
        RECT 524.400 193.000 525.200 193.200 ;
        RECT 529.000 193.000 529.800 193.200 ;
        RECT 524.400 192.400 529.800 193.000 ;
        RECT 530.400 193.000 532.600 193.600 ;
        RECT 530.400 191.800 531.000 193.000 ;
        RECT 531.800 192.800 532.600 193.000 ;
        RECT 534.200 193.200 535.600 194.000 ;
        RECT 534.200 192.200 534.800 193.200 ;
        RECT 526.200 191.400 531.000 191.800 ;
        RECT 521.200 191.200 531.000 191.400 ;
        RECT 532.400 191.600 534.800 192.200 ;
        RECT 518.000 189.600 518.800 191.200 ;
        RECT 521.200 191.000 527.000 191.200 ;
        RECT 521.200 190.800 526.800 191.000 ;
        RECT 527.600 190.200 528.400 190.400 ;
        RECT 523.400 189.600 528.400 190.200 ;
        RECT 530.800 190.300 531.600 190.400 ;
        RECT 532.400 190.300 533.000 191.600 ;
        RECT 538.800 191.200 539.600 199.800 ;
        RECT 543.000 198.400 543.800 199.800 ;
        RECT 542.000 197.600 543.800 198.400 ;
        RECT 543.000 192.400 543.800 197.600 ;
        RECT 544.400 193.600 545.200 194.400 ;
        RECT 544.600 192.400 545.200 193.600 ;
        RECT 543.000 191.800 544.000 192.400 ;
        RECT 544.600 191.800 546.000 192.400 ;
        RECT 535.400 190.600 539.600 191.200 ;
        RECT 535.400 190.400 536.200 190.600 ;
        RECT 530.800 189.700 533.100 190.300 ;
        RECT 537.000 189.800 537.800 190.000 ;
        RECT 530.800 189.600 531.600 189.700 ;
        RECT 523.400 189.400 524.200 189.600 ;
        RECT 525.000 188.400 525.800 188.600 ;
        RECT 532.400 188.400 533.000 189.700 ;
        RECT 534.000 189.200 537.800 189.800 ;
        RECT 534.000 189.000 534.800 189.200 ;
        RECT 514.800 187.800 515.800 188.200 ;
        RECT 504.400 187.200 505.200 187.600 ;
        RECT 503.800 186.200 507.400 186.600 ;
        RECT 508.600 186.200 509.200 187.600 ;
        RECT 511.600 187.200 515.800 187.800 ;
        RECT 516.800 187.600 518.800 188.400 ;
        RECT 522.000 187.800 533.000 188.400 ;
        RECT 522.000 187.600 523.600 187.800 ;
        RECT 503.600 186.000 507.600 186.200 ;
        RECT 503.600 182.200 504.400 186.000 ;
        RECT 506.800 182.800 507.600 186.000 ;
        RECT 508.400 183.400 509.200 186.200 ;
        RECT 510.000 182.800 510.800 186.200 ;
        RECT 511.600 185.000 512.200 187.200 ;
        RECT 516.800 187.000 517.400 187.600 ;
        RECT 516.600 186.600 517.400 187.000 ;
        RECT 515.800 186.000 517.400 186.600 ;
        RECT 511.600 183.000 512.400 185.000 ;
        RECT 515.800 183.000 516.600 186.000 ;
        RECT 506.800 182.200 510.800 182.800 ;
        RECT 521.200 182.200 522.000 187.000 ;
        RECT 526.200 185.600 526.800 187.800 ;
        RECT 531.800 187.600 532.600 187.800 ;
        RECT 538.800 187.200 539.600 190.600 ;
        RECT 542.000 188.800 542.800 190.400 ;
        RECT 543.400 188.400 544.000 191.800 ;
        RECT 545.200 191.600 546.000 191.800 ;
        RECT 546.800 191.600 547.600 193.200 ;
        RECT 545.300 190.300 545.900 191.600 ;
        RECT 548.400 190.300 549.200 199.800 ;
        RECT 545.300 189.700 549.200 190.300 ;
        RECT 540.400 188.200 541.200 188.400 ;
        RECT 540.400 187.600 542.000 188.200 ;
        RECT 543.400 187.600 546.000 188.400 ;
        RECT 541.200 187.200 542.000 187.600 ;
        RECT 535.800 186.600 539.600 187.200 ;
        RECT 535.800 186.400 536.600 186.600 ;
        RECT 524.400 184.200 525.200 185.000 ;
        RECT 526.000 184.800 526.800 185.600 ;
        RECT 527.800 185.400 528.600 185.600 ;
        RECT 527.800 184.800 530.600 185.400 ;
        RECT 530.000 184.200 530.600 184.800 ;
        RECT 534.000 184.200 534.800 185.000 ;
        RECT 524.400 183.600 526.400 184.200 ;
        RECT 525.600 182.200 526.400 183.600 ;
        RECT 530.000 182.200 530.800 184.200 ;
        RECT 534.000 183.600 535.400 184.200 ;
        RECT 534.200 182.200 535.400 183.600 ;
        RECT 538.800 182.200 539.600 186.600 ;
        RECT 540.600 186.200 544.200 186.600 ;
        RECT 545.200 186.200 545.800 187.600 ;
        RECT 548.400 186.200 549.200 189.700 ;
        RECT 550.000 186.800 550.800 188.400 ;
        RECT 540.400 186.000 544.400 186.200 ;
        RECT 540.400 182.200 541.200 186.000 ;
        RECT 543.600 182.200 544.400 186.000 ;
        RECT 545.200 182.200 546.000 186.200 ;
        RECT 547.400 185.600 549.200 186.200 ;
        RECT 547.400 182.200 548.200 185.600 ;
        RECT 1.200 175.600 2.000 177.200 ;
        RECT 2.800 172.300 3.600 179.800 ;
        RECT 6.000 177.800 6.800 179.800 ;
        RECT 10.800 177.800 11.600 179.800 ;
        RECT 6.000 174.400 6.600 177.800 ;
        RECT 7.600 175.600 8.400 177.200 ;
        RECT 9.200 175.600 10.000 177.200 ;
        RECT 11.000 176.300 11.600 177.800 ;
        RECT 15.600 177.800 16.400 179.800 ;
        RECT 12.400 176.300 13.200 176.400 ;
        RECT 10.900 175.700 13.200 176.300 ;
        RECT 11.000 174.400 11.600 175.700 ;
        RECT 12.400 175.600 13.200 175.700 ;
        RECT 6.000 173.600 6.800 174.400 ;
        RECT 10.800 173.600 11.600 174.400 ;
        RECT 4.400 172.300 5.200 172.400 ;
        RECT 2.800 171.700 5.200 172.300 ;
        RECT 2.800 162.200 3.600 171.700 ;
        RECT 4.400 170.800 5.200 171.700 ;
        RECT 6.000 172.300 6.600 173.600 ;
        RECT 9.200 172.300 10.000 172.400 ;
        RECT 6.000 171.700 10.000 172.300 ;
        RECT 6.000 170.200 6.600 171.700 ;
        RECT 9.200 171.600 10.000 171.700 ;
        RECT 11.000 170.200 11.600 173.600 ;
        RECT 15.600 174.400 16.200 177.800 ;
        RECT 17.200 176.300 18.000 177.200 ;
        RECT 18.800 176.300 19.600 177.200 ;
        RECT 17.200 175.700 19.600 176.300 ;
        RECT 17.200 175.600 18.000 175.700 ;
        RECT 18.800 175.600 19.600 175.700 ;
        RECT 15.600 173.600 16.400 174.400 ;
        RECT 12.400 170.800 13.200 172.400 ;
        RECT 14.000 170.800 14.800 172.400 ;
        RECT 15.600 170.400 16.200 173.600 ;
        RECT 15.600 170.200 16.400 170.400 ;
        RECT 5.000 169.400 6.800 170.200 ;
        RECT 10.800 169.400 12.600 170.200 ;
        RECT 5.000 162.200 5.800 169.400 ;
        RECT 11.800 162.200 12.600 169.400 ;
        RECT 14.600 169.400 16.400 170.200 ;
        RECT 14.600 162.200 15.400 169.400 ;
        RECT 20.400 162.200 21.200 179.800 ;
        RECT 22.000 162.200 22.800 179.800 ;
        RECT 23.600 175.600 24.400 177.200 ;
        RECT 26.400 174.200 27.200 179.800 ;
        RECT 25.400 173.800 27.200 174.200 ;
        RECT 35.200 178.400 36.000 179.800 ;
        RECT 35.200 177.600 37.200 178.400 ;
        RECT 35.200 174.200 36.000 177.600 ;
        RECT 38.000 176.000 38.800 179.800 ;
        RECT 41.200 179.200 45.200 179.800 ;
        RECT 41.200 176.000 42.000 179.200 ;
        RECT 38.000 175.800 42.000 176.000 ;
        RECT 38.200 175.400 41.800 175.800 ;
        RECT 42.800 175.600 43.600 178.600 ;
        RECT 44.400 175.800 45.200 179.200 ;
        RECT 48.600 178.400 49.400 179.800 ;
        RECT 51.400 178.400 52.200 179.800 ;
        RECT 48.600 177.600 50.000 178.400 ;
        RECT 51.400 177.600 53.200 178.400 ;
        RECT 48.600 176.400 49.400 177.600 ;
        RECT 47.600 175.800 49.400 176.400 ;
        RECT 51.400 176.400 52.200 177.600 ;
        RECT 51.400 175.800 53.200 176.400 ;
        RECT 57.200 176.000 58.000 179.800 ;
        RECT 38.800 174.400 39.600 174.800 ;
        RECT 43.000 174.400 43.600 175.600 ;
        RECT 35.200 173.800 37.000 174.200 ;
        RECT 25.400 173.600 27.000 173.800 ;
        RECT 35.400 173.600 37.000 173.800 ;
        RECT 38.000 173.800 39.600 174.400 ;
        RECT 41.200 173.800 43.600 174.400 ;
        RECT 38.000 173.600 38.800 173.800 ;
        RECT 41.200 173.600 42.000 173.800 ;
        RECT 25.400 170.400 26.000 173.600 ;
        RECT 27.600 171.600 29.200 172.400 ;
        RECT 33.200 171.600 34.800 172.400 ;
        RECT 25.200 169.600 26.000 170.400 ;
        RECT 30.000 170.300 30.800 171.200 ;
        RECT 31.600 170.300 32.400 171.200 ;
        RECT 30.000 169.700 32.400 170.300 ;
        RECT 30.000 169.600 30.800 169.700 ;
        RECT 31.600 169.600 32.400 169.700 ;
        RECT 36.400 170.400 37.000 173.600 ;
        RECT 39.600 171.600 40.400 173.200 ;
        RECT 36.400 169.600 37.200 170.400 ;
        RECT 41.200 170.200 41.800 173.600 ;
        RECT 42.800 171.600 43.600 173.200 ;
        RECT 44.400 172.800 45.200 174.400 ;
        RECT 46.000 173.600 46.800 175.200 ;
        RECT 25.400 167.000 26.000 169.600 ;
        RECT 26.800 168.300 27.600 169.200 ;
        RECT 30.000 168.300 30.800 168.400 ;
        RECT 31.600 168.300 32.400 168.400 ;
        RECT 34.800 168.300 35.600 169.200 ;
        RECT 26.800 167.700 35.600 168.300 ;
        RECT 26.800 167.600 27.600 167.700 ;
        RECT 30.000 167.600 30.800 167.700 ;
        RECT 31.600 167.600 32.400 167.700 ;
        RECT 34.800 167.600 35.600 167.700 ;
        RECT 36.400 167.000 37.000 169.600 ;
        RECT 25.400 166.400 29.000 167.000 ;
        RECT 25.400 166.200 26.000 166.400 ;
        RECT 25.200 162.200 26.000 166.200 ;
        RECT 28.400 166.200 29.000 166.400 ;
        RECT 33.400 166.400 37.000 167.000 ;
        RECT 33.400 166.200 34.000 166.400 ;
        RECT 28.400 162.200 29.200 166.200 ;
        RECT 33.200 162.200 34.000 166.200 ;
        RECT 36.400 166.200 37.000 166.400 ;
        RECT 36.400 162.200 37.200 166.200 ;
        RECT 40.600 162.200 42.600 170.200 ;
        RECT 47.600 162.200 48.400 175.800 ;
        RECT 49.200 170.300 50.000 170.400 ;
        RECT 50.800 170.300 51.600 170.400 ;
        RECT 49.200 169.700 51.600 170.300 ;
        RECT 49.200 168.800 50.000 169.700 ;
        RECT 50.800 168.800 51.600 169.700 ;
        RECT 52.400 162.200 53.200 175.800 ;
        RECT 57.000 175.200 58.000 176.000 ;
        RECT 54.000 173.600 54.800 175.200 ;
        RECT 57.000 170.800 57.800 175.200 ;
        RECT 58.800 174.600 59.600 179.800 ;
        RECT 65.200 176.600 66.000 179.800 ;
        RECT 66.800 177.000 67.600 179.800 ;
        RECT 68.400 177.000 69.200 179.800 ;
        RECT 70.000 177.000 70.800 179.800 ;
        RECT 71.600 177.000 72.400 179.800 ;
        RECT 74.800 177.000 75.600 179.800 ;
        RECT 78.000 177.000 78.800 179.800 ;
        RECT 79.600 177.000 80.400 179.800 ;
        RECT 81.200 177.000 82.000 179.800 ;
        RECT 63.600 175.800 66.000 176.600 ;
        RECT 82.800 176.600 83.600 179.800 ;
        RECT 63.600 175.200 64.400 175.800 ;
        RECT 58.400 174.000 59.600 174.600 ;
        RECT 62.600 174.600 64.400 175.200 ;
        RECT 68.400 175.600 69.400 176.400 ;
        RECT 72.400 175.600 74.000 176.400 ;
        RECT 74.800 175.800 79.400 176.400 ;
        RECT 82.800 175.800 85.400 176.600 ;
        RECT 74.800 175.600 75.600 175.800 ;
        RECT 58.400 172.000 59.000 174.000 ;
        RECT 62.600 173.400 63.400 174.600 ;
        RECT 59.600 172.600 63.400 173.400 ;
        RECT 68.400 172.800 69.200 175.600 ;
        RECT 74.800 174.800 75.600 175.000 ;
        RECT 71.200 174.200 75.600 174.800 ;
        RECT 71.200 174.000 72.000 174.200 ;
        RECT 76.400 173.600 77.200 175.200 ;
        RECT 78.600 173.400 79.400 175.800 ;
        RECT 84.600 175.200 85.400 175.800 ;
        RECT 84.600 174.400 87.600 175.200 ;
        RECT 89.200 173.800 90.000 179.800 ;
        RECT 90.800 176.000 91.600 179.800 ;
        RECT 94.000 176.000 94.800 179.800 ;
        RECT 90.800 175.800 94.800 176.000 ;
        RECT 95.600 175.800 96.400 179.800 ;
        RECT 98.800 177.800 99.600 179.800 ;
        RECT 91.000 175.400 94.600 175.800 ;
        RECT 91.600 174.400 92.400 174.800 ;
        RECT 95.600 174.400 96.200 175.800 ;
        RECT 98.800 174.400 99.400 177.800 ;
        RECT 100.400 175.600 101.200 177.200 ;
        RECT 104.600 175.800 106.200 179.800 ;
        RECT 118.000 176.000 118.800 179.800 ;
        RECT 105.200 174.400 105.800 175.800 ;
        RECT 117.800 175.200 118.800 176.000 ;
        RECT 71.600 172.600 74.800 173.400 ;
        RECT 78.600 172.600 80.600 173.400 ;
        RECT 81.200 173.000 90.000 173.800 ;
        RECT 90.800 173.800 92.400 174.400 ;
        RECT 90.800 173.600 91.600 173.800 ;
        RECT 93.800 173.600 96.400 174.400 ;
        RECT 98.800 174.300 99.600 174.400 ;
        RECT 103.600 174.300 104.400 174.400 ;
        RECT 98.800 173.700 104.400 174.300 ;
        RECT 98.800 173.600 99.600 173.700 ;
        RECT 103.600 173.600 104.400 173.700 ;
        RECT 65.200 172.000 66.000 172.600 ;
        RECT 82.800 172.000 83.600 172.400 ;
        RECT 86.000 172.000 86.800 172.400 ;
        RECT 87.800 172.000 88.600 172.200 ;
        RECT 58.400 171.400 59.200 172.000 ;
        RECT 65.200 171.400 88.600 172.000 ;
        RECT 57.000 170.000 58.000 170.800 ;
        RECT 57.200 162.200 58.000 170.000 ;
        RECT 58.600 169.600 59.200 171.400 ;
        RECT 58.600 169.000 67.600 169.600 ;
        RECT 58.600 167.400 59.200 169.000 ;
        RECT 66.800 168.800 67.600 169.000 ;
        RECT 70.000 169.000 78.600 169.600 ;
        RECT 70.000 168.800 70.800 169.000 ;
        RECT 61.800 167.600 64.400 168.400 ;
        RECT 58.600 166.800 61.200 167.400 ;
        RECT 60.400 162.200 61.200 166.800 ;
        RECT 63.600 162.200 64.400 167.600 ;
        RECT 65.000 166.800 69.200 167.600 ;
        RECT 66.800 162.200 67.600 165.000 ;
        RECT 68.400 162.200 69.200 165.000 ;
        RECT 70.000 162.200 70.800 165.000 ;
        RECT 71.600 162.200 72.400 168.400 ;
        RECT 74.800 167.600 77.400 168.400 ;
        RECT 78.000 168.200 78.600 169.000 ;
        RECT 79.600 169.400 80.400 169.600 ;
        RECT 79.600 169.000 85.000 169.400 ;
        RECT 79.600 168.800 85.800 169.000 ;
        RECT 84.400 168.200 85.800 168.800 ;
        RECT 78.000 167.600 83.800 168.200 ;
        RECT 86.800 168.000 88.400 168.800 ;
        RECT 86.800 167.600 87.400 168.000 ;
        RECT 74.800 162.200 75.600 167.000 ;
        RECT 78.000 162.200 78.800 167.000 ;
        RECT 83.200 166.800 87.400 167.600 ;
        RECT 89.200 167.400 90.000 173.000 ;
        RECT 92.400 171.600 93.200 173.200 ;
        RECT 93.800 172.300 94.400 173.600 ;
        RECT 97.200 172.300 98.000 172.400 ;
        RECT 93.800 171.700 98.000 172.300 ;
        RECT 93.800 170.200 94.400 171.700 ;
        RECT 97.200 170.800 98.000 171.700 ;
        RECT 95.600 170.200 96.400 170.400 ;
        RECT 98.800 170.200 99.400 173.600 ;
        RECT 103.800 173.200 104.400 173.600 ;
        RECT 105.200 173.600 106.000 174.400 ;
        RECT 103.800 172.400 104.600 173.200 ;
        RECT 105.200 172.400 105.800 173.600 ;
        RECT 106.800 172.800 107.600 174.400 ;
        RECT 100.400 172.300 101.200 172.400 ;
        RECT 102.000 172.300 102.800 172.400 ;
        RECT 100.400 171.700 102.800 172.300 ;
        RECT 100.400 171.600 101.200 171.700 ;
        RECT 102.000 170.800 102.800 171.700 ;
        RECT 105.200 171.600 106.000 172.400 ;
        RECT 108.400 172.300 109.200 172.400 ;
        RECT 110.000 172.300 110.800 172.400 ;
        RECT 108.400 172.200 110.800 172.300 ;
        RECT 107.600 171.700 110.800 172.200 ;
        RECT 107.600 171.600 109.200 171.700 ;
        RECT 110.000 171.600 110.800 171.700 ;
        RECT 105.200 171.400 105.800 171.600 ;
        RECT 103.800 170.800 105.800 171.400 ;
        RECT 107.600 171.200 108.400 171.600 ;
        RECT 117.800 170.800 118.600 175.200 ;
        RECT 119.600 174.600 120.400 179.800 ;
        RECT 126.000 176.600 126.800 179.800 ;
        RECT 127.600 177.000 128.400 179.800 ;
        RECT 129.200 177.000 130.000 179.800 ;
        RECT 130.800 177.000 131.600 179.800 ;
        RECT 132.400 177.000 133.200 179.800 ;
        RECT 135.600 177.000 136.400 179.800 ;
        RECT 138.800 177.000 139.600 179.800 ;
        RECT 140.400 177.000 141.200 179.800 ;
        RECT 142.000 177.000 142.800 179.800 ;
        RECT 124.400 175.800 126.800 176.600 ;
        RECT 143.600 176.600 144.400 179.800 ;
        RECT 124.400 175.200 125.200 175.800 ;
        RECT 119.200 174.000 120.400 174.600 ;
        RECT 123.400 174.600 125.200 175.200 ;
        RECT 129.200 175.600 130.200 176.400 ;
        RECT 133.200 175.600 134.800 176.400 ;
        RECT 135.600 175.800 140.200 176.400 ;
        RECT 143.600 175.800 146.200 176.600 ;
        RECT 135.600 175.600 136.400 175.800 ;
        RECT 119.200 172.000 119.800 174.000 ;
        RECT 123.400 173.400 124.200 174.600 ;
        RECT 120.400 172.600 124.200 173.400 ;
        RECT 129.200 172.800 130.000 175.600 ;
        RECT 135.600 174.800 136.400 175.000 ;
        RECT 132.000 174.200 136.400 174.800 ;
        RECT 132.000 174.000 132.800 174.200 ;
        RECT 137.200 173.600 138.000 175.200 ;
        RECT 139.400 173.400 140.200 175.800 ;
        RECT 145.400 175.200 146.200 175.800 ;
        RECT 145.400 174.400 148.400 175.200 ;
        RECT 150.000 173.800 150.800 179.800 ;
        RECT 132.400 172.600 135.600 173.400 ;
        RECT 139.400 172.600 141.400 173.400 ;
        RECT 142.000 173.000 150.800 173.800 ;
        RECT 119.200 171.400 120.000 172.000 ;
        RECT 103.800 170.200 104.400 170.800 ;
        RECT 88.000 166.800 90.000 167.400 ;
        RECT 93.400 169.600 94.400 170.200 ;
        RECT 95.000 169.600 96.400 170.200 ;
        RECT 79.600 162.200 80.400 165.000 ;
        RECT 81.200 162.200 82.000 165.000 ;
        RECT 84.400 162.200 85.200 166.800 ;
        RECT 88.000 166.200 88.600 166.800 ;
        RECT 87.600 165.600 88.600 166.200 ;
        RECT 87.600 162.200 88.400 165.600 ;
        RECT 93.400 162.200 94.200 169.600 ;
        RECT 95.000 168.400 95.600 169.600 ;
        RECT 94.800 167.600 95.600 168.400 ;
        RECT 97.800 169.400 99.600 170.200 ;
        RECT 97.800 162.200 98.600 169.400 ;
        RECT 102.000 162.800 102.800 170.200 ;
        RECT 103.600 163.400 104.400 170.200 ;
        RECT 105.200 169.600 109.200 170.200 ;
        RECT 117.800 170.000 118.800 170.800 ;
        RECT 105.200 162.800 106.000 169.600 ;
        RECT 102.000 162.200 106.000 162.800 ;
        RECT 108.400 162.200 109.200 169.600 ;
        RECT 118.000 162.200 118.800 170.000 ;
        RECT 119.400 169.600 120.000 171.400 ;
        RECT 120.600 170.800 121.400 171.000 ;
        RECT 120.600 170.200 147.600 170.800 ;
        RECT 143.400 170.000 144.200 170.200 ;
        RECT 146.800 169.600 147.600 170.200 ;
        RECT 119.400 169.000 128.400 169.600 ;
        RECT 119.400 167.400 120.000 169.000 ;
        RECT 127.600 168.800 128.400 169.000 ;
        RECT 130.800 169.000 139.400 169.600 ;
        RECT 130.800 168.800 131.600 169.000 ;
        RECT 122.600 167.600 125.200 168.400 ;
        RECT 119.400 166.800 122.000 167.400 ;
        RECT 121.200 162.200 122.000 166.800 ;
        RECT 124.400 162.200 125.200 167.600 ;
        RECT 125.800 166.800 130.000 167.600 ;
        RECT 127.600 162.200 128.400 165.000 ;
        RECT 129.200 162.200 130.000 165.000 ;
        RECT 130.800 162.200 131.600 165.000 ;
        RECT 132.400 162.200 133.200 168.400 ;
        RECT 135.600 167.600 138.200 168.400 ;
        RECT 138.800 168.200 139.400 169.000 ;
        RECT 140.400 169.400 141.200 169.600 ;
        RECT 140.400 169.000 145.800 169.400 ;
        RECT 140.400 168.800 146.600 169.000 ;
        RECT 145.200 168.200 146.600 168.800 ;
        RECT 138.800 167.600 144.600 168.200 ;
        RECT 147.600 168.000 149.200 168.800 ;
        RECT 147.600 167.600 148.200 168.000 ;
        RECT 135.600 162.200 136.400 167.000 ;
        RECT 138.800 162.200 139.600 167.000 ;
        RECT 144.000 166.800 148.200 167.600 ;
        RECT 150.000 167.400 150.800 173.000 ;
        RECT 148.800 166.800 150.800 167.400 ;
        RECT 151.600 173.800 152.400 179.800 ;
        RECT 158.000 176.600 158.800 179.800 ;
        RECT 159.600 177.000 160.400 179.800 ;
        RECT 161.200 177.000 162.000 179.800 ;
        RECT 162.800 177.000 163.600 179.800 ;
        RECT 166.000 177.000 166.800 179.800 ;
        RECT 169.200 177.000 170.000 179.800 ;
        RECT 170.800 177.000 171.600 179.800 ;
        RECT 172.400 177.000 173.200 179.800 ;
        RECT 174.000 177.000 174.800 179.800 ;
        RECT 156.200 175.800 158.800 176.600 ;
        RECT 175.600 176.600 176.400 179.800 ;
        RECT 162.200 175.800 166.800 176.400 ;
        RECT 156.200 175.200 157.000 175.800 ;
        RECT 154.000 174.400 157.000 175.200 ;
        RECT 151.600 173.000 160.400 173.800 ;
        RECT 162.200 173.400 163.000 175.800 ;
        RECT 166.000 175.600 166.800 175.800 ;
        RECT 167.600 175.600 169.200 176.400 ;
        RECT 172.200 175.600 173.200 176.400 ;
        RECT 175.600 175.800 178.000 176.600 ;
        RECT 164.400 173.600 165.200 175.200 ;
        RECT 166.000 174.800 166.800 175.000 ;
        RECT 166.000 174.200 170.400 174.800 ;
        RECT 169.600 174.000 170.400 174.200 ;
        RECT 151.600 167.400 152.400 173.000 ;
        RECT 161.000 172.600 163.000 173.400 ;
        RECT 166.800 172.600 170.000 173.400 ;
        RECT 172.400 172.800 173.200 175.600 ;
        RECT 177.200 175.200 178.000 175.800 ;
        RECT 177.200 174.600 179.000 175.200 ;
        RECT 178.200 173.400 179.000 174.600 ;
        RECT 182.000 174.600 182.800 179.800 ;
        RECT 183.600 176.000 184.400 179.800 ;
        RECT 189.400 176.400 190.200 179.800 ;
        RECT 191.800 176.400 192.600 177.200 ;
        RECT 188.400 176.300 190.200 176.400 ;
        RECT 191.600 176.300 192.400 176.400 ;
        RECT 183.600 175.200 184.600 176.000 ;
        RECT 188.400 175.700 192.400 176.300 ;
        RECT 182.000 174.000 183.200 174.600 ;
        RECT 178.200 172.600 182.000 173.400 ;
        RECT 153.200 172.200 154.000 172.400 ;
        RECT 153.000 172.000 154.000 172.200 ;
        RECT 158.000 172.000 158.800 172.400 ;
        RECT 175.600 172.000 176.400 172.600 ;
        RECT 182.600 172.000 183.200 174.000 ;
        RECT 153.000 171.400 176.400 172.000 ;
        RECT 182.400 171.400 183.200 172.000 ;
        RECT 182.400 169.600 183.000 171.400 ;
        RECT 183.800 170.800 184.600 175.200 ;
        RECT 186.800 173.600 187.600 175.200 ;
        RECT 161.200 169.400 162.000 169.600 ;
        RECT 156.600 169.000 162.000 169.400 ;
        RECT 155.800 168.800 162.000 169.000 ;
        RECT 163.000 169.000 171.600 169.600 ;
        RECT 153.200 168.000 154.800 168.800 ;
        RECT 155.800 168.200 157.200 168.800 ;
        RECT 163.000 168.200 163.600 169.000 ;
        RECT 170.800 168.800 171.600 169.000 ;
        RECT 174.000 169.000 183.000 169.600 ;
        RECT 174.000 168.800 174.800 169.000 ;
        RECT 154.200 167.600 154.800 168.000 ;
        RECT 157.800 167.600 163.600 168.200 ;
        RECT 164.200 167.600 166.800 168.400 ;
        RECT 151.600 166.800 153.600 167.400 ;
        RECT 154.200 166.800 158.400 167.600 ;
        RECT 140.400 162.200 141.200 165.000 ;
        RECT 142.000 162.200 142.800 165.000 ;
        RECT 145.200 162.200 146.000 166.800 ;
        RECT 148.800 166.200 149.400 166.800 ;
        RECT 148.400 165.600 149.400 166.200 ;
        RECT 153.000 166.200 153.600 166.800 ;
        RECT 153.000 165.600 154.000 166.200 ;
        RECT 148.400 162.200 149.200 165.600 ;
        RECT 153.200 162.200 154.000 165.600 ;
        RECT 156.400 162.200 157.200 166.800 ;
        RECT 159.600 162.200 160.400 165.000 ;
        RECT 161.200 162.200 162.000 165.000 ;
        RECT 162.800 162.200 163.600 167.000 ;
        RECT 166.000 162.200 166.800 167.000 ;
        RECT 169.200 162.200 170.000 168.400 ;
        RECT 177.200 167.600 179.800 168.400 ;
        RECT 172.400 166.800 176.600 167.600 ;
        RECT 170.800 162.200 171.600 165.000 ;
        RECT 172.400 162.200 173.200 165.000 ;
        RECT 174.000 162.200 174.800 165.000 ;
        RECT 177.200 162.200 178.000 167.600 ;
        RECT 182.400 167.400 183.000 169.000 ;
        RECT 180.400 166.800 183.000 167.400 ;
        RECT 183.600 170.000 184.600 170.800 ;
        RECT 180.400 162.200 181.200 166.800 ;
        RECT 183.600 162.200 184.400 170.000 ;
        RECT 188.400 162.200 189.200 175.700 ;
        RECT 191.600 175.600 192.400 175.700 ;
        RECT 193.200 175.600 194.000 179.800 ;
        RECT 191.600 172.200 192.400 172.400 ;
        RECT 193.400 172.200 194.000 175.600 ;
        RECT 194.800 174.300 195.600 174.400 ;
        RECT 198.000 174.300 198.800 179.800 ;
        RECT 199.600 175.600 200.400 177.200 ;
        RECT 202.800 176.000 203.600 179.800 ;
        RECT 194.800 173.700 198.800 174.300 ;
        RECT 194.800 172.800 195.600 173.700 ;
        RECT 196.400 172.200 197.200 172.400 ;
        RECT 191.600 171.600 194.000 172.200 ;
        RECT 195.600 171.600 197.200 172.200 ;
        RECT 190.000 168.800 190.800 170.400 ;
        RECT 191.800 170.200 192.400 171.600 ;
        RECT 195.600 171.200 196.400 171.600 ;
        RECT 191.600 162.200 192.400 170.200 ;
        RECT 193.200 169.600 197.200 170.200 ;
        RECT 193.200 162.200 194.000 169.600 ;
        RECT 196.400 162.200 197.200 169.600 ;
        RECT 198.000 162.200 198.800 173.700 ;
        RECT 202.600 175.200 203.600 176.000 ;
        RECT 202.600 170.800 203.400 175.200 ;
        RECT 204.400 174.600 205.200 179.800 ;
        RECT 210.800 176.600 211.600 179.800 ;
        RECT 212.400 177.000 213.200 179.800 ;
        RECT 214.000 177.000 214.800 179.800 ;
        RECT 215.600 177.000 216.400 179.800 ;
        RECT 217.200 177.000 218.000 179.800 ;
        RECT 220.400 177.000 221.200 179.800 ;
        RECT 223.600 177.000 224.400 179.800 ;
        RECT 225.200 177.000 226.000 179.800 ;
        RECT 226.800 177.000 227.600 179.800 ;
        RECT 209.200 175.800 211.600 176.600 ;
        RECT 228.400 176.600 229.200 179.800 ;
        RECT 209.200 175.200 210.000 175.800 ;
        RECT 204.000 174.000 205.200 174.600 ;
        RECT 208.200 174.600 210.000 175.200 ;
        RECT 214.000 175.600 215.000 176.400 ;
        RECT 218.000 175.600 219.600 176.400 ;
        RECT 220.400 175.800 225.000 176.400 ;
        RECT 228.400 175.800 231.000 176.600 ;
        RECT 220.400 175.600 221.200 175.800 ;
        RECT 204.000 172.000 204.600 174.000 ;
        RECT 208.200 173.400 209.000 174.600 ;
        RECT 205.200 172.600 209.000 173.400 ;
        RECT 214.000 172.800 214.800 175.600 ;
        RECT 220.400 174.800 221.200 175.000 ;
        RECT 216.800 174.200 221.200 174.800 ;
        RECT 216.800 174.000 217.600 174.200 ;
        RECT 222.000 173.600 222.800 175.200 ;
        RECT 224.200 173.400 225.000 175.800 ;
        RECT 230.200 175.200 231.000 175.800 ;
        RECT 230.200 174.400 233.200 175.200 ;
        RECT 234.800 173.800 235.600 179.800 ;
        RECT 236.600 176.400 237.400 177.200 ;
        RECT 236.400 175.600 237.200 176.400 ;
        RECT 238.000 175.800 238.800 179.800 ;
        RECT 238.200 174.400 238.800 175.800 ;
        RECT 217.200 172.600 220.400 173.400 ;
        RECT 224.200 172.600 226.200 173.400 ;
        RECT 226.800 173.000 235.600 173.800 ;
        RECT 238.000 173.600 238.800 174.400 ;
        RECT 210.800 172.000 211.600 172.600 ;
        RECT 222.000 172.000 222.800 172.400 ;
        RECT 228.400 172.000 229.200 172.400 ;
        RECT 233.400 172.000 234.200 172.200 ;
        RECT 204.000 171.400 204.800 172.000 ;
        RECT 210.800 171.400 234.200 172.000 ;
        RECT 202.600 170.000 203.600 170.800 ;
        RECT 202.800 162.200 203.600 170.000 ;
        RECT 204.200 169.600 204.800 171.400 ;
        RECT 204.200 169.000 213.200 169.600 ;
        RECT 204.200 167.400 204.800 169.000 ;
        RECT 212.400 168.800 213.200 169.000 ;
        RECT 215.600 169.000 224.200 169.600 ;
        RECT 215.600 168.800 216.400 169.000 ;
        RECT 207.400 167.600 210.000 168.400 ;
        RECT 204.200 166.800 206.800 167.400 ;
        RECT 206.000 162.200 206.800 166.800 ;
        RECT 209.200 162.200 210.000 167.600 ;
        RECT 210.600 166.800 214.800 167.600 ;
        RECT 212.400 162.200 213.200 165.000 ;
        RECT 214.000 162.200 214.800 165.000 ;
        RECT 215.600 162.200 216.400 165.000 ;
        RECT 217.200 162.200 218.000 168.400 ;
        RECT 220.400 167.600 223.000 168.400 ;
        RECT 223.600 168.200 224.200 169.000 ;
        RECT 225.200 169.400 226.000 169.600 ;
        RECT 225.200 169.000 230.600 169.400 ;
        RECT 225.200 168.800 231.400 169.000 ;
        RECT 230.000 168.200 231.400 168.800 ;
        RECT 223.600 167.600 229.400 168.200 ;
        RECT 232.400 168.000 234.000 168.800 ;
        RECT 232.400 167.600 233.000 168.000 ;
        RECT 220.400 162.200 221.200 167.000 ;
        RECT 223.600 162.200 224.400 167.000 ;
        RECT 228.800 166.800 233.000 167.600 ;
        RECT 234.800 167.400 235.600 173.000 ;
        RECT 236.400 172.200 237.200 172.400 ;
        RECT 238.200 172.200 238.800 173.600 ;
        RECT 239.600 174.300 240.400 174.400 ;
        RECT 242.800 174.300 243.600 179.800 ;
        RECT 244.400 175.600 245.200 177.200 ;
        RECT 246.000 175.800 246.800 179.800 ;
        RECT 247.600 176.000 248.400 179.800 ;
        RECT 250.800 176.000 251.600 179.800 ;
        RECT 247.600 175.800 251.600 176.000 ;
        RECT 253.000 178.400 253.800 179.800 ;
        RECT 253.000 177.600 254.800 178.400 ;
        RECT 253.000 176.400 253.800 177.600 ;
        RECT 257.400 176.400 258.200 177.200 ;
        RECT 253.000 175.800 254.800 176.400 ;
        RECT 246.200 174.400 246.800 175.800 ;
        RECT 247.800 175.400 251.400 175.800 ;
        RECT 250.000 174.400 250.800 174.800 ;
        RECT 239.600 173.700 243.600 174.300 ;
        RECT 239.600 172.800 240.400 173.700 ;
        RECT 241.200 172.200 242.000 172.400 ;
        RECT 236.400 171.600 238.800 172.200 ;
        RECT 240.400 171.600 242.000 172.200 ;
        RECT 236.600 170.200 237.200 171.600 ;
        RECT 240.400 171.200 241.200 171.600 ;
        RECT 233.600 166.800 235.600 167.400 ;
        RECT 225.200 162.200 226.000 165.000 ;
        RECT 226.800 162.200 227.600 165.000 ;
        RECT 230.000 162.200 230.800 166.800 ;
        RECT 233.600 166.200 234.200 166.800 ;
        RECT 233.200 165.600 234.200 166.200 ;
        RECT 233.200 162.200 234.000 165.600 ;
        RECT 236.400 162.200 237.200 170.200 ;
        RECT 238.000 169.600 242.000 170.200 ;
        RECT 238.000 162.200 238.800 169.600 ;
        RECT 241.200 162.200 242.000 169.600 ;
        RECT 242.800 162.200 243.600 173.700 ;
        RECT 246.000 173.600 248.600 174.400 ;
        RECT 250.000 173.800 251.600 174.400 ;
        RECT 250.800 173.600 251.600 173.800 ;
        RECT 246.000 170.200 246.800 170.400 ;
        RECT 248.000 170.200 248.600 173.600 ;
        RECT 249.200 171.600 250.000 173.200 ;
        RECT 246.000 169.600 247.400 170.200 ;
        RECT 248.000 169.600 249.000 170.200 ;
        RECT 246.800 168.400 247.400 169.600 ;
        RECT 246.800 167.600 247.600 168.400 ;
        RECT 248.200 162.200 249.000 169.600 ;
        RECT 252.400 168.800 253.200 170.400 ;
        RECT 254.000 162.200 254.800 175.800 ;
        RECT 257.200 175.600 258.000 176.400 ;
        RECT 258.800 175.800 259.600 179.800 ;
        RECT 255.600 173.600 256.400 175.200 ;
        RECT 257.200 172.200 258.000 172.400 ;
        RECT 259.000 172.200 259.600 175.800 ;
        RECT 264.800 174.400 265.600 179.800 ;
        RECT 270.200 176.400 271.000 177.200 ;
        RECT 270.000 175.600 270.800 176.400 ;
        RECT 271.600 175.800 272.400 179.800 ;
        RECT 282.800 176.000 283.600 179.800 ;
        RECT 286.000 176.000 286.800 179.800 ;
        RECT 282.800 175.800 286.800 176.000 ;
        RECT 287.600 175.800 288.400 179.800 ;
        RECT 290.800 177.800 291.600 179.800 ;
        RECT 260.400 172.800 261.200 174.400 ;
        RECT 264.800 174.200 266.000 174.400 ;
        RECT 263.800 173.600 266.000 174.200 ;
        RECT 262.000 172.200 262.800 172.400 ;
        RECT 257.200 171.600 259.600 172.200 ;
        RECT 261.200 171.600 262.800 172.200 ;
        RECT 257.400 170.200 258.000 171.600 ;
        RECT 261.200 171.200 262.000 171.600 ;
        RECT 263.800 170.400 264.400 173.600 ;
        RECT 266.000 171.600 267.600 172.400 ;
        RECT 270.000 172.200 270.800 172.400 ;
        RECT 271.800 172.200 272.400 175.800 ;
        RECT 283.000 175.400 286.600 175.800 ;
        RECT 283.600 174.400 284.400 174.800 ;
        RECT 287.600 174.400 288.200 175.800 ;
        RECT 289.200 175.600 290.000 177.200 ;
        RECT 291.000 176.400 291.600 177.800 ;
        RECT 290.800 175.600 291.600 176.400 ;
        RECT 295.600 176.000 296.400 179.800 ;
        RECT 291.000 174.400 291.600 175.600 ;
        RECT 273.200 172.800 274.000 174.400 ;
        RECT 282.800 173.800 284.400 174.400 ;
        RECT 282.800 173.600 283.600 173.800 ;
        RECT 285.800 173.600 288.400 174.400 ;
        RECT 290.800 173.600 291.600 174.400 ;
        RECT 274.800 172.300 275.600 172.400 ;
        RECT 281.200 172.300 282.000 172.400 ;
        RECT 274.800 172.200 282.000 172.300 ;
        RECT 270.000 171.600 272.400 172.200 ;
        RECT 274.000 171.700 282.000 172.200 ;
        RECT 274.000 171.600 275.600 171.700 ;
        RECT 281.200 171.600 282.000 171.700 ;
        RECT 284.400 171.600 285.200 173.200 ;
        RECT 257.200 162.200 258.000 170.200 ;
        RECT 258.800 169.600 262.800 170.200 ;
        RECT 263.600 169.600 264.400 170.400 ;
        RECT 268.400 169.600 269.200 171.200 ;
        RECT 270.200 170.200 270.800 171.600 ;
        RECT 274.000 171.200 274.800 171.600 ;
        RECT 285.800 170.200 286.400 173.600 ;
        RECT 287.600 170.200 288.400 170.400 ;
        RECT 291.000 170.200 291.600 173.600 ;
        RECT 295.400 175.200 296.400 176.000 ;
        RECT 292.400 172.300 293.200 172.400 ;
        RECT 295.400 172.300 296.200 175.200 ;
        RECT 297.200 174.600 298.000 179.800 ;
        RECT 303.600 176.600 304.400 179.800 ;
        RECT 305.200 177.000 306.000 179.800 ;
        RECT 306.800 177.000 307.600 179.800 ;
        RECT 308.400 177.000 309.200 179.800 ;
        RECT 310.000 177.000 310.800 179.800 ;
        RECT 313.200 177.000 314.000 179.800 ;
        RECT 316.400 177.000 317.200 179.800 ;
        RECT 318.000 177.000 318.800 179.800 ;
        RECT 319.600 177.000 320.400 179.800 ;
        RECT 302.000 175.800 304.400 176.600 ;
        RECT 321.200 176.600 322.000 179.800 ;
        RECT 302.000 175.200 302.800 175.800 ;
        RECT 292.400 171.700 296.200 172.300 ;
        RECT 292.400 170.800 293.200 171.700 ;
        RECT 295.400 170.800 296.200 171.700 ;
        RECT 296.800 174.000 298.000 174.600 ;
        RECT 301.000 174.600 302.800 175.200 ;
        RECT 306.800 175.600 307.800 176.400 ;
        RECT 310.800 175.600 312.400 176.400 ;
        RECT 313.200 175.800 317.800 176.400 ;
        RECT 321.200 175.800 323.800 176.600 ;
        RECT 313.200 175.600 314.000 175.800 ;
        RECT 296.800 172.000 297.400 174.000 ;
        RECT 301.000 173.400 301.800 174.600 ;
        RECT 298.000 172.600 301.800 173.400 ;
        RECT 306.800 172.800 307.600 175.600 ;
        RECT 313.200 174.800 314.000 175.000 ;
        RECT 309.600 174.200 314.000 174.800 ;
        RECT 309.600 174.000 310.400 174.200 ;
        RECT 314.800 173.600 315.600 175.200 ;
        RECT 317.000 173.400 317.800 175.800 ;
        RECT 323.000 175.200 323.800 175.800 ;
        RECT 323.000 174.400 326.000 175.200 ;
        RECT 327.600 173.800 328.400 179.800 ;
        RECT 329.800 176.400 330.600 179.800 ;
        RECT 329.800 175.800 331.600 176.400 ;
        RECT 310.000 172.600 313.200 173.400 ;
        RECT 317.000 172.600 319.000 173.400 ;
        RECT 319.600 173.000 328.400 173.800 ;
        RECT 303.600 172.000 304.400 172.600 ;
        RECT 321.200 172.000 322.000 172.400 ;
        RECT 324.400 172.000 325.200 172.400 ;
        RECT 326.200 172.000 327.000 172.200 ;
        RECT 296.800 171.400 297.600 172.000 ;
        RECT 303.600 171.400 327.000 172.000 ;
        RECT 258.800 162.200 259.600 169.600 ;
        RECT 262.000 162.200 262.800 169.600 ;
        RECT 263.800 167.000 264.400 169.600 ;
        RECT 265.200 167.600 266.000 169.200 ;
        RECT 263.800 166.400 267.400 167.000 ;
        RECT 263.800 166.200 264.400 166.400 ;
        RECT 263.600 162.200 264.400 166.200 ;
        RECT 266.800 166.200 267.400 166.400 ;
        RECT 266.800 162.200 267.600 166.200 ;
        RECT 270.000 162.200 270.800 170.200 ;
        RECT 271.600 169.600 275.600 170.200 ;
        RECT 271.600 162.200 272.400 169.600 ;
        RECT 274.800 162.200 275.600 169.600 ;
        RECT 285.400 169.600 286.400 170.200 ;
        RECT 287.000 169.600 288.400 170.200 ;
        RECT 285.400 162.200 286.200 169.600 ;
        RECT 287.000 168.400 287.600 169.600 ;
        RECT 290.800 169.400 292.600 170.200 ;
        RECT 295.400 170.000 296.400 170.800 ;
        RECT 286.800 167.600 287.600 168.400 ;
        RECT 291.800 162.200 292.600 169.400 ;
        RECT 295.600 162.200 296.400 170.000 ;
        RECT 297.000 169.600 297.600 171.400 ;
        RECT 297.000 169.000 306.000 169.600 ;
        RECT 297.000 167.400 297.600 169.000 ;
        RECT 305.200 168.800 306.000 169.000 ;
        RECT 308.400 169.000 317.000 169.600 ;
        RECT 308.400 168.800 309.200 169.000 ;
        RECT 300.200 167.600 302.800 168.400 ;
        RECT 297.000 166.800 299.600 167.400 ;
        RECT 298.800 162.200 299.600 166.800 ;
        RECT 302.000 162.200 302.800 167.600 ;
        RECT 303.400 166.800 307.600 167.600 ;
        RECT 305.200 162.200 306.000 165.000 ;
        RECT 306.800 162.200 307.600 165.000 ;
        RECT 308.400 162.200 309.200 165.000 ;
        RECT 310.000 162.200 310.800 168.400 ;
        RECT 313.200 167.600 315.800 168.400 ;
        RECT 316.400 168.200 317.000 169.000 ;
        RECT 318.000 169.400 318.800 169.600 ;
        RECT 318.000 169.000 323.400 169.400 ;
        RECT 318.000 168.800 324.200 169.000 ;
        RECT 322.800 168.200 324.200 168.800 ;
        RECT 316.400 167.600 322.200 168.200 ;
        RECT 325.200 168.000 326.800 168.800 ;
        RECT 325.200 167.600 325.800 168.000 ;
        RECT 313.200 162.200 314.000 167.000 ;
        RECT 316.400 162.200 317.200 167.000 ;
        RECT 321.600 166.800 325.800 167.600 ;
        RECT 327.600 167.400 328.400 173.000 ;
        RECT 329.200 168.800 330.000 170.400 ;
        RECT 326.400 166.800 328.400 167.400 ;
        RECT 318.000 162.200 318.800 165.000 ;
        RECT 319.600 162.200 320.400 165.000 ;
        RECT 322.800 162.200 323.600 166.800 ;
        RECT 326.400 166.200 327.000 166.800 ;
        RECT 326.000 165.600 327.000 166.200 ;
        RECT 326.000 162.200 326.800 165.600 ;
        RECT 330.800 162.200 331.600 175.800 ;
        RECT 334.000 175.600 334.800 177.200 ;
        RECT 332.400 173.600 333.200 175.200 ;
        RECT 335.600 174.300 336.400 179.800 ;
        RECT 337.200 176.000 338.000 179.800 ;
        RECT 340.400 176.000 341.200 179.800 ;
        RECT 337.200 175.800 341.200 176.000 ;
        RECT 342.000 175.800 342.800 179.800 ;
        RECT 343.600 175.800 344.400 179.800 ;
        RECT 345.200 176.000 346.000 179.800 ;
        RECT 348.400 176.000 349.200 179.800 ;
        RECT 345.200 175.800 349.200 176.000 ;
        RECT 337.400 175.400 341.000 175.800 ;
        RECT 338.000 174.400 338.800 174.800 ;
        RECT 342.000 174.400 342.600 175.800 ;
        RECT 343.800 174.400 344.400 175.800 ;
        RECT 345.400 175.400 349.000 175.800 ;
        RECT 350.000 175.200 350.800 179.800 ;
        RECT 347.600 174.400 348.400 174.800 ;
        RECT 350.000 174.600 352.200 175.200 ;
        RECT 337.200 174.300 338.800 174.400 ;
        RECT 335.600 173.800 338.800 174.300 ;
        RECT 335.600 173.700 338.000 173.800 ;
        RECT 335.600 162.200 336.400 173.700 ;
        RECT 337.200 173.600 338.000 173.700 ;
        RECT 340.200 173.600 342.800 174.400 ;
        RECT 343.600 173.600 346.200 174.400 ;
        RECT 347.600 173.800 349.200 174.400 ;
        RECT 348.400 173.600 349.200 173.800 ;
        RECT 338.800 171.600 339.600 173.200 ;
        RECT 340.200 170.200 340.800 173.600 ;
        RECT 345.600 172.300 346.200 173.600 ;
        RECT 342.100 171.700 346.200 172.300 ;
        RECT 342.100 170.400 342.700 171.700 ;
        RECT 342.000 170.200 342.800 170.400 ;
        RECT 339.800 169.600 340.800 170.200 ;
        RECT 341.400 169.600 342.800 170.200 ;
        RECT 343.600 170.200 344.400 170.400 ;
        RECT 345.600 170.200 346.200 171.700 ;
        RECT 351.600 171.600 352.200 174.600 ;
        RECT 353.200 172.400 354.000 179.800 ;
        RECT 351.600 170.800 352.800 171.600 ;
        RECT 351.600 170.200 352.200 170.800 ;
        RECT 353.400 170.200 354.000 172.400 ;
        RECT 343.600 169.600 345.000 170.200 ;
        RECT 345.600 169.600 346.600 170.200 ;
        RECT 339.800 162.200 340.600 169.600 ;
        RECT 341.400 168.400 342.000 169.600 ;
        RECT 341.200 167.600 342.000 168.400 ;
        RECT 344.400 168.400 345.000 169.600 ;
        RECT 344.400 167.600 345.200 168.400 ;
        RECT 345.800 162.200 346.600 169.600 ;
        RECT 350.000 169.600 352.200 170.200 ;
        RECT 350.000 162.200 350.800 169.600 ;
        RECT 353.200 162.200 354.000 170.200 ;
        RECT 354.800 174.300 355.600 179.800 ;
        RECT 356.400 175.600 357.200 177.200 ;
        RECT 358.000 176.000 358.800 179.800 ;
        RECT 361.200 176.000 362.000 179.800 ;
        RECT 358.000 175.800 362.000 176.000 ;
        RECT 362.800 175.800 363.600 179.800 ;
        RECT 358.200 175.400 361.800 175.800 ;
        RECT 358.800 174.400 359.600 174.800 ;
        RECT 362.800 174.400 363.400 175.800 ;
        RECT 358.000 174.300 359.600 174.400 ;
        RECT 354.800 173.800 359.600 174.300 ;
        RECT 354.800 173.700 358.800 173.800 ;
        RECT 354.800 162.200 355.600 173.700 ;
        RECT 358.000 173.600 358.800 173.700 ;
        RECT 361.000 173.600 363.600 174.400 ;
        RECT 364.400 173.800 365.200 179.800 ;
        RECT 370.800 176.600 371.600 179.800 ;
        RECT 372.400 177.000 373.200 179.800 ;
        RECT 374.000 177.000 374.800 179.800 ;
        RECT 375.600 177.000 376.400 179.800 ;
        RECT 378.800 177.000 379.600 179.800 ;
        RECT 382.000 177.000 382.800 179.800 ;
        RECT 383.600 177.000 384.400 179.800 ;
        RECT 385.200 177.000 386.000 179.800 ;
        RECT 386.800 177.000 387.600 179.800 ;
        RECT 369.000 175.800 371.600 176.600 ;
        RECT 388.400 176.600 389.200 179.800 ;
        RECT 375.000 175.800 379.600 176.400 ;
        RECT 369.000 175.200 369.800 175.800 ;
        RECT 366.800 174.400 369.800 175.200 ;
        RECT 359.600 171.600 360.400 173.200 ;
        RECT 361.000 170.200 361.600 173.600 ;
        RECT 364.400 173.000 373.200 173.800 ;
        RECT 375.000 173.400 375.800 175.800 ;
        RECT 378.800 175.600 379.600 175.800 ;
        RECT 380.400 175.600 382.000 176.400 ;
        RECT 385.000 175.600 386.000 176.400 ;
        RECT 388.400 175.800 390.800 176.600 ;
        RECT 377.200 173.600 378.000 175.200 ;
        RECT 378.800 174.800 379.600 175.000 ;
        RECT 378.800 174.200 383.200 174.800 ;
        RECT 382.400 174.000 383.200 174.200 ;
        RECT 362.800 170.200 363.600 170.400 ;
        RECT 360.600 169.600 361.600 170.200 ;
        RECT 362.200 169.600 363.600 170.200 ;
        RECT 360.600 162.200 361.400 169.600 ;
        RECT 362.200 168.400 362.800 169.600 ;
        RECT 362.000 167.600 362.800 168.400 ;
        RECT 364.400 167.400 365.200 173.000 ;
        RECT 373.800 172.600 375.800 173.400 ;
        RECT 379.600 172.600 382.800 173.400 ;
        RECT 385.200 172.800 386.000 175.600 ;
        RECT 390.000 175.200 390.800 175.800 ;
        RECT 390.000 174.600 391.800 175.200 ;
        RECT 391.000 173.400 391.800 174.600 ;
        RECT 394.800 174.600 395.600 179.800 ;
        RECT 396.400 176.000 397.200 179.800 ;
        RECT 396.400 175.200 397.400 176.000 ;
        RECT 394.800 174.000 396.000 174.600 ;
        RECT 391.000 172.600 394.800 173.400 ;
        RECT 365.800 172.000 366.600 172.200 ;
        RECT 370.800 172.000 371.600 172.400 ;
        RECT 388.400 172.000 389.200 172.600 ;
        RECT 395.400 172.000 396.000 174.000 ;
        RECT 365.800 171.400 389.200 172.000 ;
        RECT 395.200 171.400 396.000 172.000 ;
        RECT 395.200 169.600 395.800 171.400 ;
        RECT 396.600 170.800 397.400 175.200 ;
        RECT 400.800 174.200 401.600 179.800 ;
        RECT 374.000 169.400 374.800 169.600 ;
        RECT 369.400 169.000 374.800 169.400 ;
        RECT 368.600 168.800 374.800 169.000 ;
        RECT 375.800 169.000 384.400 169.600 ;
        RECT 366.000 168.000 367.600 168.800 ;
        RECT 368.600 168.200 370.000 168.800 ;
        RECT 375.800 168.200 376.400 169.000 ;
        RECT 383.600 168.800 384.400 169.000 ;
        RECT 386.800 169.000 395.800 169.600 ;
        RECT 386.800 168.800 387.600 169.000 ;
        RECT 367.000 167.600 367.600 168.000 ;
        RECT 370.600 167.600 376.400 168.200 ;
        RECT 377.000 167.600 379.600 168.400 ;
        RECT 364.400 166.800 366.400 167.400 ;
        RECT 367.000 166.800 371.200 167.600 ;
        RECT 365.800 166.200 366.400 166.800 ;
        RECT 365.800 165.600 366.800 166.200 ;
        RECT 366.000 162.200 366.800 165.600 ;
        RECT 369.200 162.200 370.000 166.800 ;
        RECT 372.400 162.200 373.200 165.000 ;
        RECT 374.000 162.200 374.800 165.000 ;
        RECT 375.600 162.200 376.400 167.000 ;
        RECT 378.800 162.200 379.600 167.000 ;
        RECT 382.000 162.200 382.800 168.400 ;
        RECT 390.000 167.600 392.600 168.400 ;
        RECT 385.200 166.800 389.400 167.600 ;
        RECT 383.600 162.200 384.400 165.000 ;
        RECT 385.200 162.200 386.000 165.000 ;
        RECT 386.800 162.200 387.600 165.000 ;
        RECT 390.000 162.200 390.800 167.600 ;
        RECT 395.200 167.400 395.800 169.000 ;
        RECT 393.200 166.800 395.800 167.400 ;
        RECT 396.400 170.000 397.400 170.800 ;
        RECT 399.800 173.800 401.600 174.200 ;
        RECT 407.600 177.800 408.400 179.800 ;
        RECT 407.600 174.400 408.200 177.800 ;
        RECT 409.200 175.600 410.000 177.200 ;
        RECT 410.800 176.300 411.600 176.400 ;
        RECT 418.800 176.300 419.600 179.800 ;
        RECT 410.800 175.700 419.600 176.300 ;
        RECT 410.800 175.600 411.600 175.700 ;
        RECT 418.600 175.200 419.600 175.700 ;
        RECT 399.800 173.600 401.400 173.800 ;
        RECT 407.600 173.600 408.400 174.400 ;
        RECT 399.800 170.400 400.400 173.600 ;
        RECT 402.000 171.600 403.600 172.400 ;
        RECT 393.200 162.200 394.000 166.800 ;
        RECT 396.400 162.200 397.200 170.000 ;
        RECT 399.600 169.600 400.400 170.400 ;
        RECT 402.800 170.300 403.600 170.400 ;
        RECT 404.400 170.300 405.200 171.200 ;
        RECT 406.000 170.800 406.800 172.400 ;
        RECT 402.800 169.700 405.200 170.300 ;
        RECT 407.600 170.200 408.200 173.600 ;
        RECT 418.600 170.800 419.400 175.200 ;
        RECT 420.400 174.600 421.200 179.800 ;
        RECT 426.800 176.600 427.600 179.800 ;
        RECT 428.400 177.000 429.200 179.800 ;
        RECT 430.000 177.000 430.800 179.800 ;
        RECT 431.600 177.000 432.400 179.800 ;
        RECT 433.200 177.000 434.000 179.800 ;
        RECT 436.400 177.000 437.200 179.800 ;
        RECT 439.600 177.000 440.400 179.800 ;
        RECT 441.200 177.000 442.000 179.800 ;
        RECT 442.800 177.000 443.600 179.800 ;
        RECT 425.200 175.800 427.600 176.600 ;
        RECT 444.400 176.600 445.200 179.800 ;
        RECT 425.200 175.200 426.000 175.800 ;
        RECT 420.000 174.000 421.200 174.600 ;
        RECT 424.200 174.600 426.000 175.200 ;
        RECT 430.000 175.600 431.000 176.400 ;
        RECT 434.000 175.600 435.600 176.400 ;
        RECT 436.400 175.800 441.000 176.400 ;
        RECT 444.400 175.800 447.000 176.600 ;
        RECT 436.400 175.600 437.200 175.800 ;
        RECT 420.000 172.000 420.600 174.000 ;
        RECT 424.200 173.400 425.000 174.600 ;
        RECT 421.200 172.600 425.000 173.400 ;
        RECT 430.000 172.800 430.800 175.600 ;
        RECT 436.400 174.800 437.200 175.000 ;
        RECT 432.800 174.200 437.200 174.800 ;
        RECT 432.800 174.000 433.600 174.200 ;
        RECT 438.000 173.600 438.800 175.200 ;
        RECT 440.200 173.400 441.000 175.800 ;
        RECT 446.200 175.200 447.000 175.800 ;
        RECT 446.200 174.400 449.200 175.200 ;
        RECT 450.800 173.800 451.600 179.800 ;
        RECT 433.200 172.600 436.400 173.400 ;
        RECT 440.200 172.600 442.200 173.400 ;
        RECT 442.800 173.000 451.600 173.800 ;
        RECT 426.800 172.000 427.600 172.600 ;
        RECT 444.400 172.000 445.200 172.400 ;
        RECT 447.600 172.000 448.400 172.400 ;
        RECT 449.400 172.000 450.200 172.200 ;
        RECT 420.000 171.400 420.800 172.000 ;
        RECT 426.800 171.400 450.200 172.000 ;
        RECT 402.800 169.600 403.600 169.700 ;
        RECT 404.400 169.600 405.200 169.700 ;
        RECT 399.800 167.000 400.400 169.600 ;
        RECT 406.600 169.400 408.400 170.200 ;
        RECT 418.600 170.000 419.600 170.800 ;
        RECT 401.200 168.300 402.000 169.200 ;
        RECT 404.400 168.300 405.200 168.400 ;
        RECT 401.200 167.700 405.200 168.300 ;
        RECT 401.200 167.600 402.000 167.700 ;
        RECT 404.400 167.600 405.200 167.700 ;
        RECT 399.800 166.400 403.400 167.000 ;
        RECT 399.800 166.200 400.400 166.400 ;
        RECT 399.600 162.200 400.400 166.200 ;
        RECT 402.800 166.200 403.400 166.400 ;
        RECT 402.800 162.200 403.600 166.200 ;
        RECT 406.600 164.400 407.400 169.400 ;
        RECT 406.600 163.600 408.400 164.400 ;
        RECT 406.600 162.200 407.400 163.600 ;
        RECT 418.800 162.200 419.600 170.000 ;
        RECT 420.200 169.600 420.800 171.400 ;
        RECT 420.200 169.000 429.200 169.600 ;
        RECT 420.200 167.400 420.800 169.000 ;
        RECT 428.400 168.800 429.200 169.000 ;
        RECT 431.600 169.000 440.200 169.600 ;
        RECT 431.600 168.800 432.400 169.000 ;
        RECT 423.400 167.600 426.000 168.400 ;
        RECT 420.200 166.800 422.800 167.400 ;
        RECT 422.000 162.200 422.800 166.800 ;
        RECT 425.200 162.200 426.000 167.600 ;
        RECT 426.600 166.800 430.800 167.600 ;
        RECT 428.400 162.200 429.200 165.000 ;
        RECT 430.000 162.200 430.800 165.000 ;
        RECT 431.600 162.200 432.400 165.000 ;
        RECT 433.200 162.200 434.000 168.400 ;
        RECT 436.400 167.600 439.000 168.400 ;
        RECT 439.600 168.200 440.200 169.000 ;
        RECT 441.200 169.400 442.000 169.600 ;
        RECT 441.200 169.000 446.600 169.400 ;
        RECT 441.200 168.800 447.400 169.000 ;
        RECT 446.000 168.200 447.400 168.800 ;
        RECT 439.600 167.600 445.400 168.200 ;
        RECT 448.400 168.000 450.000 168.800 ;
        RECT 448.400 167.600 449.000 168.000 ;
        RECT 436.400 162.200 437.200 167.000 ;
        RECT 439.600 162.200 440.400 167.000 ;
        RECT 444.800 166.800 449.000 167.600 ;
        RECT 450.800 167.400 451.600 173.000 ;
        RECT 454.000 177.800 454.800 179.800 ;
        RECT 454.000 174.400 454.600 177.800 ;
        RECT 455.600 175.600 456.400 177.200 ;
        RECT 454.000 173.600 454.800 174.400 ;
        RECT 458.800 174.300 459.600 179.800 ;
        RECT 463.600 177.600 464.400 179.800 ;
        RECT 463.600 174.400 464.200 177.600 ;
        RECT 460.400 174.300 461.200 174.400 ;
        RECT 458.800 173.700 461.200 174.300 ;
        RECT 452.400 170.800 453.200 172.400 ;
        RECT 454.000 170.200 454.600 173.600 ;
        RECT 455.600 172.300 456.400 172.400 ;
        RECT 458.800 172.300 459.600 173.700 ;
        RECT 460.400 173.600 461.200 173.700 ;
        RECT 463.600 173.600 464.400 174.400 ;
        RECT 468.000 174.200 468.800 179.800 ;
        RECT 474.400 178.400 475.200 179.800 ;
        RECT 474.400 177.600 475.600 178.400 ;
        RECT 474.400 174.200 475.200 177.600 ;
        RECT 467.000 173.800 468.800 174.200 ;
        RECT 473.400 173.800 475.200 174.200 ;
        RECT 467.000 173.600 468.600 173.800 ;
        RECT 473.400 173.600 475.000 173.800 ;
        RECT 455.600 171.700 459.600 172.300 ;
        RECT 455.600 171.600 456.400 171.700 ;
        RECT 449.600 166.800 451.600 167.400 ;
        RECT 453.000 169.400 454.800 170.200 ;
        RECT 441.200 162.200 442.000 165.000 ;
        RECT 442.800 162.200 443.600 165.000 ;
        RECT 446.000 162.200 446.800 166.800 ;
        RECT 449.600 166.200 450.200 166.800 ;
        RECT 449.200 165.600 450.200 166.200 ;
        RECT 449.200 162.200 450.000 165.600 ;
        RECT 453.000 164.400 453.800 169.400 ;
        RECT 453.000 163.600 454.800 164.400 ;
        RECT 453.000 162.200 453.800 163.600 ;
        RECT 458.800 162.200 459.600 171.700 ;
        RECT 463.600 170.200 464.200 173.600 ;
        RECT 467.000 170.400 467.600 173.600 ;
        RECT 469.200 171.600 470.800 172.400 ;
        RECT 473.400 170.400 474.000 173.600 ;
        RECT 462.600 169.400 464.400 170.200 ;
        RECT 466.800 169.600 467.600 170.400 ;
        RECT 473.200 169.600 474.000 170.400 ;
        RECT 462.600 162.200 463.400 169.400 ;
        RECT 467.000 167.000 467.600 169.600 ;
        RECT 468.400 167.600 469.200 169.200 ;
        RECT 473.400 167.000 474.000 169.600 ;
        RECT 474.800 167.600 475.600 169.200 ;
        RECT 467.000 166.400 470.600 167.000 ;
        RECT 466.800 162.200 467.600 166.400 ;
        RECT 470.000 166.200 470.600 166.400 ;
        RECT 473.400 166.400 477.000 167.000 ;
        RECT 473.400 166.200 474.000 166.400 ;
        RECT 470.000 162.200 470.800 166.200 ;
        RECT 473.200 162.200 474.000 166.200 ;
        RECT 476.400 166.200 477.000 166.400 ;
        RECT 476.400 162.200 477.200 166.200 ;
        RECT 479.600 162.200 480.400 179.800 ;
        RECT 486.400 178.400 487.200 179.800 ;
        RECT 486.400 177.600 488.400 178.400 ;
        RECT 486.400 174.200 487.200 177.600 ;
        RECT 486.400 173.800 488.200 174.200 ;
        RECT 486.600 173.600 488.200 173.800 ;
        RECT 484.400 171.600 486.000 172.400 ;
        RECT 487.600 170.400 488.200 173.600 ;
        RECT 487.600 169.600 488.400 170.400 ;
        RECT 486.000 167.600 486.800 169.200 ;
        RECT 487.600 167.000 488.200 169.600 ;
        RECT 484.600 166.400 488.200 167.000 ;
        RECT 484.600 166.200 485.200 166.400 ;
        RECT 484.400 162.200 485.200 166.200 ;
        RECT 487.600 166.200 488.200 166.400 ;
        RECT 487.600 162.200 488.400 166.200 ;
        RECT 489.200 162.200 490.000 179.800 ;
        RECT 493.600 174.200 494.400 179.800 ;
        RECT 492.600 173.800 494.400 174.200 ;
        RECT 492.600 173.600 494.200 173.800 ;
        RECT 498.800 173.600 499.600 175.200 ;
        RECT 500.400 174.300 501.200 179.800 ;
        RECT 502.200 176.400 503.000 177.200 ;
        RECT 502.000 175.600 502.800 176.400 ;
        RECT 503.600 175.800 504.400 179.800 ;
        RECT 511.000 178.400 511.800 179.800 ;
        RECT 511.000 177.600 512.400 178.400 ;
        RECT 511.000 176.400 511.800 177.600 ;
        RECT 502.000 174.300 502.800 174.400 ;
        RECT 500.400 173.700 502.800 174.300 ;
        RECT 492.600 170.400 493.200 173.600 ;
        RECT 492.400 169.600 493.200 170.400 ;
        RECT 492.600 167.000 493.200 169.600 ;
        RECT 494.000 167.600 494.800 169.200 ;
        RECT 492.600 166.400 496.200 167.000 ;
        RECT 492.600 166.200 493.200 166.400 ;
        RECT 492.400 162.200 493.200 166.200 ;
        RECT 495.600 166.200 496.200 166.400 ;
        RECT 495.600 162.200 496.400 166.200 ;
        RECT 500.400 162.200 501.200 173.700 ;
        RECT 502.000 173.600 502.800 173.700 ;
        RECT 502.000 172.200 502.800 172.400 ;
        RECT 503.800 172.200 504.400 175.800 ;
        RECT 510.000 175.800 511.800 176.400 ;
        RECT 514.800 176.000 515.600 179.800 ;
        RECT 505.200 172.800 506.000 174.400 ;
        RECT 508.400 173.600 509.200 175.200 ;
        RECT 506.800 172.200 507.600 172.400 ;
        RECT 502.000 171.600 504.400 172.200 ;
        RECT 506.000 171.600 507.600 172.200 ;
        RECT 502.200 170.200 502.800 171.600 ;
        RECT 506.000 171.200 506.800 171.600 ;
        RECT 502.000 162.200 502.800 170.200 ;
        RECT 503.600 169.600 507.600 170.200 ;
        RECT 503.600 162.200 504.400 169.600 ;
        RECT 506.800 162.200 507.600 169.600 ;
        RECT 510.000 162.200 510.800 175.800 ;
        RECT 514.600 175.200 515.600 176.000 ;
        RECT 514.600 170.800 515.400 175.200 ;
        RECT 516.400 174.600 517.200 179.800 ;
        RECT 522.800 176.600 523.600 179.800 ;
        RECT 524.400 177.000 525.200 179.800 ;
        RECT 526.000 177.000 526.800 179.800 ;
        RECT 527.600 177.000 528.400 179.800 ;
        RECT 529.200 177.000 530.000 179.800 ;
        RECT 532.400 177.000 533.200 179.800 ;
        RECT 535.600 177.000 536.400 179.800 ;
        RECT 537.200 177.000 538.000 179.800 ;
        RECT 538.800 177.000 539.600 179.800 ;
        RECT 521.200 175.800 523.600 176.600 ;
        RECT 540.400 176.600 541.200 179.800 ;
        RECT 521.200 175.200 522.000 175.800 ;
        RECT 516.000 174.000 517.200 174.600 ;
        RECT 520.200 174.600 522.000 175.200 ;
        RECT 526.000 175.600 527.000 176.400 ;
        RECT 530.000 175.600 531.600 176.400 ;
        RECT 532.400 175.800 537.000 176.400 ;
        RECT 540.400 175.800 543.000 176.600 ;
        RECT 532.400 175.600 533.200 175.800 ;
        RECT 516.000 172.000 516.600 174.000 ;
        RECT 520.200 173.400 521.000 174.600 ;
        RECT 522.800 173.600 523.600 174.400 ;
        RECT 517.200 172.600 521.000 173.400 ;
        RECT 522.900 172.600 523.500 173.600 ;
        RECT 526.000 172.800 526.800 175.600 ;
        RECT 532.400 174.800 533.200 175.000 ;
        RECT 528.800 174.200 533.200 174.800 ;
        RECT 528.800 174.000 529.600 174.200 ;
        RECT 534.000 173.600 534.800 175.200 ;
        RECT 536.200 173.400 537.000 175.800 ;
        RECT 542.200 175.200 543.000 175.800 ;
        RECT 542.200 174.400 545.200 175.200 ;
        RECT 546.800 173.800 547.600 179.800 ;
        RECT 529.200 172.600 532.400 173.400 ;
        RECT 536.200 172.600 538.200 173.400 ;
        RECT 538.800 173.000 547.600 173.800 ;
        RECT 522.800 172.000 523.600 172.600 ;
        RECT 540.400 172.000 541.200 172.400 ;
        RECT 545.400 172.000 546.200 172.200 ;
        RECT 516.000 171.400 516.800 172.000 ;
        RECT 522.800 171.400 546.200 172.000 ;
        RECT 511.600 168.800 512.400 170.400 ;
        RECT 514.600 170.000 515.600 170.800 ;
        RECT 514.800 162.200 515.600 170.000 ;
        RECT 516.200 169.600 516.800 171.400 ;
        RECT 516.200 169.000 525.200 169.600 ;
        RECT 516.200 167.400 516.800 169.000 ;
        RECT 524.400 168.800 525.200 169.000 ;
        RECT 527.600 169.000 536.200 169.600 ;
        RECT 527.600 168.800 528.400 169.000 ;
        RECT 519.400 167.600 522.000 168.400 ;
        RECT 516.200 166.800 518.800 167.400 ;
        RECT 518.000 162.200 518.800 166.800 ;
        RECT 521.200 162.200 522.000 167.600 ;
        RECT 522.600 166.800 526.800 167.600 ;
        RECT 524.400 162.200 525.200 165.000 ;
        RECT 526.000 162.200 526.800 165.000 ;
        RECT 527.600 162.200 528.400 165.000 ;
        RECT 529.200 162.200 530.000 168.400 ;
        RECT 532.400 167.600 535.000 168.400 ;
        RECT 535.600 168.200 536.200 169.000 ;
        RECT 537.200 169.400 538.000 169.600 ;
        RECT 537.200 169.000 542.600 169.400 ;
        RECT 537.200 168.800 543.400 169.000 ;
        RECT 542.000 168.200 543.400 168.800 ;
        RECT 535.600 167.600 541.400 168.200 ;
        RECT 544.400 168.000 546.000 168.800 ;
        RECT 544.400 167.600 545.000 168.000 ;
        RECT 532.400 162.200 533.200 167.000 ;
        RECT 535.600 162.200 536.400 167.000 ;
        RECT 540.800 166.800 545.000 167.600 ;
        RECT 546.800 167.400 547.600 173.000 ;
        RECT 545.600 166.800 547.600 167.400 ;
        RECT 537.200 162.200 538.000 165.000 ;
        RECT 538.800 162.200 539.600 165.000 ;
        RECT 542.000 162.200 542.800 166.800 ;
        RECT 545.600 166.200 546.200 166.800 ;
        RECT 545.200 165.600 546.200 166.200 ;
        RECT 545.200 162.200 546.000 165.600 ;
        RECT 4.400 152.400 5.200 159.800 ;
        RECT 7.600 155.800 8.400 159.800 ;
        RECT 7.800 155.600 8.400 155.800 ;
        RECT 10.800 155.800 11.600 159.800 ;
        RECT 12.600 159.200 16.200 159.800 ;
        RECT 12.600 159.000 13.200 159.200 ;
        RECT 10.800 155.600 11.400 155.800 ;
        RECT 7.800 155.000 11.400 155.600 ;
        RECT 7.600 154.300 8.400 154.400 ;
        RECT 9.200 154.300 10.000 154.400 ;
        RECT 7.600 153.700 10.000 154.300 ;
        RECT 7.600 153.600 8.400 153.700 ;
        RECT 9.200 152.800 10.000 153.700 ;
        RECT 10.800 152.400 11.400 155.000 ;
        RECT 12.400 153.000 13.200 159.000 ;
        RECT 15.600 159.000 16.200 159.200 ;
        RECT 17.200 159.200 21.200 159.800 ;
        RECT 14.000 153.000 14.800 158.600 ;
        RECT 15.600 153.400 16.400 159.000 ;
        RECT 17.200 154.000 18.000 159.200 ;
        RECT 18.800 153.800 19.600 158.600 ;
        RECT 20.400 153.800 21.200 159.200 ;
        RECT 18.800 153.400 19.400 153.800 ;
        RECT 15.600 153.000 19.400 153.400 ;
        RECT 14.200 152.400 14.800 153.000 ;
        RECT 15.800 152.800 19.400 153.000 ;
        RECT 20.600 153.200 21.200 153.800 ;
        RECT 23.600 153.800 24.400 159.800 ;
        RECT 23.600 153.200 24.200 153.800 ;
        RECT 20.600 152.600 24.200 153.200 ;
        RECT 3.000 151.800 5.200 152.400 ;
        RECT 3.000 151.200 3.600 151.800 ;
        RECT 2.400 150.400 3.600 151.200 ;
        RECT 6.000 150.800 6.800 152.400 ;
        RECT 10.800 151.600 11.600 152.400 ;
        RECT 14.000 152.200 14.800 152.400 ;
        RECT 14.000 151.600 17.400 152.200 ;
        RECT 3.000 147.400 3.600 150.400 ;
        RECT 4.400 148.800 5.200 150.400 ;
        RECT 7.600 149.600 9.200 150.400 ;
        RECT 10.800 148.400 11.400 151.600 ;
        RECT 9.800 148.200 11.400 148.400 ;
        RECT 9.600 147.800 11.400 148.200 ;
        RECT 3.000 146.800 5.200 147.400 ;
        RECT 4.400 142.200 5.200 146.800 ;
        RECT 7.600 144.300 8.400 144.400 ;
        RECT 9.600 144.300 10.400 147.800 ;
        RECT 7.600 143.700 10.400 144.300 ;
        RECT 16.800 145.000 17.400 151.600 ;
        RECT 18.000 149.600 19.600 150.400 ;
        RECT 19.600 147.600 21.200 148.400 ;
        RECT 26.800 148.300 27.600 159.800 ;
        RECT 31.000 152.600 31.800 159.800 ;
        RECT 35.800 154.400 36.600 159.800 ;
        RECT 35.800 153.600 37.200 154.400 ;
        RECT 35.800 152.600 36.600 153.600 ;
        RECT 30.000 151.800 31.800 152.600 ;
        RECT 34.800 151.800 36.600 152.600 ;
        RECT 28.400 150.300 29.200 150.400 ;
        RECT 30.200 150.300 30.800 151.800 ;
        RECT 28.400 149.700 30.800 150.300 ;
        RECT 28.400 149.600 29.200 149.700 ;
        RECT 30.200 148.400 30.800 149.700 ;
        RECT 31.600 149.600 32.400 151.200 ;
        RECT 35.000 148.400 35.600 151.800 ;
        RECT 36.400 149.600 37.200 151.200 ;
        RECT 22.100 147.700 27.600 148.300 ;
        RECT 22.100 146.400 22.700 147.700 ;
        RECT 21.000 145.600 22.800 146.400 ;
        RECT 16.800 144.400 20.800 145.000 ;
        RECT 25.200 144.800 26.000 146.400 ;
        RECT 16.800 144.200 18.000 144.400 ;
        RECT 7.600 143.600 8.400 143.700 ;
        RECT 9.600 142.200 10.400 143.700 ;
        RECT 17.200 142.200 18.000 144.200 ;
        RECT 20.200 143.600 21.200 144.400 ;
        RECT 20.400 142.200 21.200 143.600 ;
        RECT 26.800 142.200 27.600 147.700 ;
        RECT 30.000 147.600 30.800 148.400 ;
        RECT 34.800 147.600 35.600 148.400 ;
        RECT 28.400 144.800 29.200 146.400 ;
        RECT 30.200 144.200 30.800 147.600 ;
        RECT 33.200 144.800 34.000 146.400 ;
        RECT 35.000 144.200 35.600 147.600 ;
        RECT 36.400 146.300 37.200 146.400 ;
        RECT 38.000 146.300 38.800 159.800 ;
        RECT 41.200 146.800 42.000 148.400 ;
        RECT 36.400 145.700 38.800 146.300 ;
        RECT 36.400 145.600 37.200 145.700 ;
        RECT 30.000 142.200 30.800 144.200 ;
        RECT 34.800 142.200 35.600 144.200 ;
        RECT 38.000 142.200 38.800 145.700 ;
        RECT 39.600 144.800 40.400 146.400 ;
        RECT 42.800 146.200 43.600 159.800 ;
        RECT 46.000 153.800 46.800 159.800 ;
        RECT 46.200 153.200 46.800 153.800 ;
        RECT 49.200 159.200 53.200 159.800 ;
        RECT 49.200 153.800 50.000 159.200 ;
        RECT 50.800 153.800 51.600 158.600 ;
        RECT 52.400 154.000 53.200 159.200 ;
        RECT 54.200 159.200 57.800 159.800 ;
        RECT 54.200 159.000 54.800 159.200 ;
        RECT 49.200 153.200 49.800 153.800 ;
        RECT 44.400 151.600 45.200 153.200 ;
        RECT 46.200 152.600 49.800 153.200 ;
        RECT 51.000 153.400 51.600 153.800 ;
        RECT 54.000 153.400 54.800 159.000 ;
        RECT 57.200 159.000 57.800 159.200 ;
        RECT 51.000 153.000 54.800 153.400 ;
        RECT 55.600 153.000 56.400 158.600 ;
        RECT 57.200 153.000 58.000 159.000 ;
        RECT 51.000 152.800 54.600 153.000 ;
        RECT 55.600 152.400 56.200 153.000 ;
        RECT 61.400 152.400 62.200 159.800 ;
        RECT 62.800 153.600 63.600 154.400 ;
        RECT 63.000 152.400 63.600 153.600 ;
        RECT 55.600 152.200 56.400 152.400 ;
        RECT 53.000 151.600 56.400 152.200 ;
        RECT 61.400 151.800 62.400 152.400 ;
        RECT 63.000 151.800 64.400 152.400 ;
        RECT 50.800 149.600 52.400 150.400 ;
        RECT 44.400 148.300 45.200 148.400 ;
        RECT 49.200 148.300 50.800 148.400 ;
        RECT 44.400 147.700 50.800 148.300 ;
        RECT 44.400 147.600 45.200 147.700 ;
        RECT 49.200 147.600 50.800 147.700 ;
        RECT 42.800 145.600 44.600 146.200 ;
        RECT 47.600 145.600 50.000 146.400 ;
        RECT 43.800 142.200 44.600 145.600 ;
        RECT 53.000 145.000 53.600 151.600 ;
        RECT 58.800 150.300 59.600 150.400 ;
        RECT 60.400 150.300 61.200 150.400 ;
        RECT 58.800 149.700 61.200 150.300 ;
        RECT 58.800 149.600 59.600 149.700 ;
        RECT 60.400 148.800 61.200 149.700 ;
        RECT 61.800 148.400 62.400 151.800 ;
        RECT 63.600 151.600 64.400 151.800 ;
        RECT 65.200 151.600 66.000 153.200 ;
        RECT 63.700 150.300 64.300 151.600 ;
        RECT 66.800 150.300 67.600 159.800 ;
        RECT 71.600 152.000 72.400 159.800 ;
        RECT 74.800 155.200 75.600 159.800 ;
        RECT 63.700 149.700 67.600 150.300 ;
        RECT 57.200 148.300 58.000 148.400 ;
        RECT 58.800 148.300 59.600 148.400 ;
        RECT 57.200 148.200 59.600 148.300 ;
        RECT 61.800 148.300 64.400 148.400 ;
        RECT 65.200 148.300 66.000 148.400 ;
        RECT 57.200 147.700 60.400 148.200 ;
        RECT 57.200 147.600 58.000 147.700 ;
        RECT 58.800 147.600 60.400 147.700 ;
        RECT 61.800 147.700 66.000 148.300 ;
        RECT 61.800 147.600 64.400 147.700 ;
        RECT 65.200 147.600 66.000 147.700 ;
        RECT 59.600 147.200 60.400 147.600 ;
        RECT 59.000 146.200 62.600 146.600 ;
        RECT 63.600 146.200 64.200 147.600 ;
        RECT 66.800 146.200 67.600 149.700 ;
        RECT 71.400 151.200 72.400 152.000 ;
        RECT 73.000 154.600 75.600 155.200 ;
        RECT 73.000 153.000 73.600 154.600 ;
        RECT 78.000 154.400 78.800 159.800 ;
        RECT 81.200 157.000 82.000 159.800 ;
        RECT 82.800 157.000 83.600 159.800 ;
        RECT 84.400 157.000 85.200 159.800 ;
        RECT 79.400 154.400 83.600 155.200 ;
        RECT 76.200 153.600 78.800 154.400 ;
        RECT 86.000 153.600 86.800 159.800 ;
        RECT 89.200 155.000 90.000 159.800 ;
        RECT 92.400 155.000 93.200 159.800 ;
        RECT 94.000 157.000 94.800 159.800 ;
        RECT 95.600 157.000 96.400 159.800 ;
        RECT 98.800 155.200 99.600 159.800 ;
        RECT 102.000 156.400 102.800 159.800 ;
        RECT 102.000 155.800 103.000 156.400 ;
        RECT 102.400 155.200 103.000 155.800 ;
        RECT 97.600 154.400 101.800 155.200 ;
        RECT 102.400 154.600 104.400 155.200 ;
        RECT 89.200 153.600 91.800 154.400 ;
        RECT 92.400 153.800 98.200 154.400 ;
        RECT 101.200 154.000 101.800 154.400 ;
        RECT 81.200 153.000 82.000 153.200 ;
        RECT 73.000 152.400 82.000 153.000 ;
        RECT 84.400 153.000 85.200 153.200 ;
        RECT 92.400 153.000 93.000 153.800 ;
        RECT 98.800 153.200 100.200 153.800 ;
        RECT 101.200 153.200 102.800 154.000 ;
        RECT 84.400 152.400 93.000 153.000 ;
        RECT 94.000 153.000 100.200 153.200 ;
        RECT 94.000 152.600 99.400 153.000 ;
        RECT 94.000 152.400 94.800 152.600 ;
        RECT 68.400 148.300 69.200 148.400 ;
        RECT 71.400 148.300 72.200 151.200 ;
        RECT 73.000 150.600 73.600 152.400 ;
        RECT 68.400 147.700 72.200 148.300 ;
        RECT 68.400 146.800 69.200 147.700 ;
        RECT 71.400 146.800 72.200 147.700 ;
        RECT 72.800 150.000 73.600 150.600 ;
        RECT 79.600 150.000 103.000 150.600 ;
        RECT 72.800 148.000 73.400 150.000 ;
        RECT 79.600 149.400 80.400 150.000 ;
        RECT 97.200 149.600 98.000 150.000 ;
        RECT 100.400 149.600 101.200 150.000 ;
        RECT 102.200 149.800 103.000 150.000 ;
        RECT 74.000 148.600 77.800 149.400 ;
        RECT 72.800 147.400 74.000 148.000 ;
        RECT 49.600 144.400 53.600 145.000 ;
        RECT 49.200 143.600 50.200 144.400 ;
        RECT 52.400 144.200 53.600 144.400 ;
        RECT 58.800 146.000 62.800 146.200 ;
        RECT 49.200 142.200 50.000 143.600 ;
        RECT 52.400 142.200 53.200 144.200 ;
        RECT 58.800 142.200 59.600 146.000 ;
        RECT 62.000 142.200 62.800 146.000 ;
        RECT 63.600 142.200 64.400 146.200 ;
        RECT 65.800 145.600 67.600 146.200 ;
        RECT 71.400 146.000 72.400 146.800 ;
        RECT 65.800 142.200 66.600 145.600 ;
        RECT 71.600 142.200 72.400 146.000 ;
        RECT 73.200 142.200 74.000 147.400 ;
        RECT 77.000 147.400 77.800 148.600 ;
        RECT 77.000 146.800 78.800 147.400 ;
        RECT 78.000 146.200 78.800 146.800 ;
        RECT 82.800 146.400 83.600 149.200 ;
        RECT 86.000 148.600 89.200 149.400 ;
        RECT 93.000 148.600 95.000 149.400 ;
        RECT 103.600 149.000 104.400 154.600 ;
        RECT 105.800 152.600 106.600 159.800 ;
        RECT 105.800 151.800 107.600 152.600 ;
        RECT 106.800 151.600 107.600 151.800 ;
        RECT 105.200 149.600 106.000 151.200 ;
        RECT 85.600 147.800 86.400 148.000 ;
        RECT 85.600 147.200 90.000 147.800 ;
        RECT 89.200 147.000 90.000 147.200 ;
        RECT 90.800 146.800 91.600 148.400 ;
        RECT 78.000 145.400 80.400 146.200 ;
        RECT 82.800 145.600 83.800 146.400 ;
        RECT 86.800 145.600 88.400 146.400 ;
        RECT 89.200 146.200 90.000 146.400 ;
        RECT 93.000 146.200 93.800 148.600 ;
        RECT 95.600 148.200 104.400 149.000 ;
        RECT 99.000 146.800 102.000 147.600 ;
        RECT 99.000 146.200 99.800 146.800 ;
        RECT 89.200 145.600 93.800 146.200 ;
        RECT 79.600 142.200 80.400 145.400 ;
        RECT 97.200 145.400 99.800 146.200 ;
        RECT 81.200 142.200 82.000 145.000 ;
        RECT 82.800 142.200 83.600 145.000 ;
        RECT 84.400 142.200 85.200 145.000 ;
        RECT 86.000 142.200 86.800 145.000 ;
        RECT 89.200 142.200 90.000 145.000 ;
        RECT 92.400 142.200 93.200 145.000 ;
        RECT 94.000 142.200 94.800 145.000 ;
        RECT 95.600 142.200 96.400 145.000 ;
        RECT 97.200 142.200 98.000 145.400 ;
        RECT 103.600 142.200 104.400 148.200 ;
        RECT 106.800 148.400 107.400 151.600 ;
        RECT 106.800 147.600 107.600 148.400 ;
        RECT 108.400 148.300 109.200 148.400 ;
        RECT 110.000 148.300 110.800 148.400 ;
        RECT 108.400 147.700 110.800 148.300 ;
        RECT 108.400 147.600 109.200 147.700 ;
        RECT 106.800 144.200 107.400 147.600 ;
        RECT 108.500 146.400 109.100 147.600 ;
        RECT 110.000 146.800 110.800 147.700 ;
        RECT 111.600 148.300 112.400 159.800 ;
        RECT 115.800 152.400 116.600 159.800 ;
        RECT 117.200 153.600 118.000 154.400 ;
        RECT 117.400 152.400 118.000 153.600 ;
        RECT 115.800 151.800 116.800 152.400 ;
        RECT 117.400 151.800 118.800 152.400 ;
        RECT 114.800 148.800 115.600 150.400 ;
        RECT 116.200 148.400 116.800 151.800 ;
        RECT 118.000 151.600 118.800 151.800 ;
        RECT 113.200 148.300 114.000 148.400 ;
        RECT 111.600 148.200 114.000 148.300 ;
        RECT 111.600 147.700 114.800 148.200 ;
        RECT 108.400 144.800 109.200 146.400 ;
        RECT 106.800 142.200 107.600 144.200 ;
        RECT 111.600 142.200 112.400 147.700 ;
        RECT 113.200 147.600 114.800 147.700 ;
        RECT 116.200 147.600 118.800 148.400 ;
        RECT 114.000 147.200 114.800 147.600 ;
        RECT 113.400 146.200 117.000 146.600 ;
        RECT 118.000 146.200 118.600 147.600 ;
        RECT 113.200 146.000 117.200 146.200 ;
        RECT 113.200 142.200 114.000 146.000 ;
        RECT 116.400 142.200 117.200 146.000 ;
        RECT 118.000 142.200 118.800 146.200 ;
        RECT 119.600 144.800 120.400 146.400 ;
        RECT 121.200 142.200 122.000 159.800 ;
        RECT 129.200 151.400 130.000 159.800 ;
        RECT 133.600 156.400 134.400 159.800 ;
        RECT 132.400 155.800 134.400 156.400 ;
        RECT 138.000 155.800 138.800 159.800 ;
        RECT 142.200 155.800 143.400 159.800 ;
        RECT 132.400 155.000 133.200 155.800 ;
        RECT 138.000 155.200 138.600 155.800 ;
        RECT 135.800 154.600 139.400 155.200 ;
        RECT 142.000 155.000 142.800 155.800 ;
        RECT 135.800 154.400 136.600 154.600 ;
        RECT 138.600 154.400 139.400 154.600 ;
        RECT 132.400 153.000 133.200 153.200 ;
        RECT 137.000 153.000 137.800 153.200 ;
        RECT 132.400 152.400 137.800 153.000 ;
        RECT 138.400 153.000 140.600 153.600 ;
        RECT 138.400 151.800 139.000 153.000 ;
        RECT 139.800 152.800 140.600 153.000 ;
        RECT 142.200 153.200 143.600 154.000 ;
        RECT 142.200 152.200 142.800 153.200 ;
        RECT 134.200 151.400 139.000 151.800 ;
        RECT 129.200 151.200 139.000 151.400 ;
        RECT 140.400 151.600 142.800 152.200 ;
        RECT 129.200 151.000 135.000 151.200 ;
        RECT 129.200 150.800 134.800 151.000 ;
        RECT 135.600 150.200 136.400 150.400 ;
        RECT 131.400 149.600 136.400 150.200 ;
        RECT 131.400 149.400 132.200 149.600 ;
        RECT 133.000 148.400 133.800 148.600 ;
        RECT 140.400 148.400 141.000 151.600 ;
        RECT 146.800 151.200 147.600 159.800 ;
        RECT 150.000 156.400 150.800 159.800 ;
        RECT 149.800 155.800 150.800 156.400 ;
        RECT 149.800 155.200 150.400 155.800 ;
        RECT 153.200 155.200 154.000 159.800 ;
        RECT 156.400 157.000 157.200 159.800 ;
        RECT 158.000 157.000 158.800 159.800 ;
        RECT 143.400 150.600 147.600 151.200 ;
        RECT 143.400 150.400 144.200 150.600 ;
        RECT 145.000 149.800 145.800 150.000 ;
        RECT 142.000 149.200 145.800 149.800 ;
        RECT 142.000 149.000 142.800 149.200 ;
        RECT 130.000 147.800 141.000 148.400 ;
        RECT 130.000 147.600 131.600 147.800 ;
        RECT 134.000 147.600 134.800 147.800 ;
        RECT 139.800 147.600 140.600 147.800 ;
        RECT 129.200 142.200 130.000 147.000 ;
        RECT 134.200 145.600 134.800 147.600 ;
        RECT 146.800 147.200 147.600 150.600 ;
        RECT 143.800 146.600 147.600 147.200 ;
        RECT 143.800 146.400 144.600 146.600 ;
        RECT 132.400 144.200 133.200 145.000 ;
        RECT 134.000 144.800 134.800 145.600 ;
        RECT 135.800 145.400 136.600 145.600 ;
        RECT 135.800 144.800 138.600 145.400 ;
        RECT 138.000 144.200 138.600 144.800 ;
        RECT 142.000 144.200 142.800 145.000 ;
        RECT 132.400 143.600 134.400 144.200 ;
        RECT 133.600 142.200 134.400 143.600 ;
        RECT 138.000 142.200 138.800 144.200 ;
        RECT 142.000 143.600 143.400 144.200 ;
        RECT 142.200 142.200 143.400 143.600 ;
        RECT 146.800 142.200 147.600 146.600 ;
        RECT 148.400 154.600 150.400 155.200 ;
        RECT 148.400 149.000 149.200 154.600 ;
        RECT 151.000 154.400 155.200 155.200 ;
        RECT 159.600 155.000 160.400 159.800 ;
        RECT 162.800 155.000 163.600 159.800 ;
        RECT 151.000 154.000 151.600 154.400 ;
        RECT 150.000 153.200 151.600 154.000 ;
        RECT 154.600 153.800 160.400 154.400 ;
        RECT 152.600 153.200 154.000 153.800 ;
        RECT 152.600 153.000 158.800 153.200 ;
        RECT 153.400 152.600 158.800 153.000 ;
        RECT 158.000 152.400 158.800 152.600 ;
        RECT 159.800 153.000 160.400 153.800 ;
        RECT 161.000 153.600 163.600 154.400 ;
        RECT 166.000 153.600 166.800 159.800 ;
        RECT 167.600 157.000 168.400 159.800 ;
        RECT 169.200 157.000 170.000 159.800 ;
        RECT 170.800 157.000 171.600 159.800 ;
        RECT 169.200 154.400 173.400 155.200 ;
        RECT 174.000 154.400 174.800 159.800 ;
        RECT 177.200 155.200 178.000 159.800 ;
        RECT 177.200 154.600 179.800 155.200 ;
        RECT 174.000 153.600 176.600 154.400 ;
        RECT 167.600 153.000 168.400 153.200 ;
        RECT 159.800 152.400 168.400 153.000 ;
        RECT 170.800 153.000 171.600 153.200 ;
        RECT 179.200 153.000 179.800 154.600 ;
        RECT 170.800 152.400 179.800 153.000 ;
        RECT 179.200 150.600 179.800 152.400 ;
        RECT 180.400 152.000 181.200 159.800 ;
        RECT 186.200 152.400 187.000 159.800 ;
        RECT 187.600 153.600 188.400 154.400 ;
        RECT 190.000 154.300 190.800 154.400 ;
        RECT 191.600 154.300 192.400 159.800 ;
        RECT 190.000 153.700 192.400 154.300 ;
        RECT 190.000 153.600 190.800 153.700 ;
        RECT 187.800 152.400 188.400 153.600 ;
        RECT 180.400 151.200 181.400 152.000 ;
        RECT 186.200 151.800 187.200 152.400 ;
        RECT 187.800 151.800 189.200 152.400 ;
        RECT 149.800 150.000 173.200 150.600 ;
        RECT 179.200 150.000 180.000 150.600 ;
        RECT 149.800 149.800 150.600 150.000 ;
        RECT 151.600 149.600 152.400 150.000 ;
        RECT 154.800 149.600 155.600 150.000 ;
        RECT 172.400 149.400 173.200 150.000 ;
        RECT 148.400 148.200 157.200 149.000 ;
        RECT 157.800 148.600 159.800 149.400 ;
        RECT 163.600 148.600 166.800 149.400 ;
        RECT 148.400 142.200 149.200 148.200 ;
        RECT 150.800 146.800 153.800 147.600 ;
        RECT 153.000 146.200 153.800 146.800 ;
        RECT 159.000 146.200 159.800 148.600 ;
        RECT 161.200 146.800 162.000 148.400 ;
        RECT 166.400 147.800 167.200 148.000 ;
        RECT 162.800 147.200 167.200 147.800 ;
        RECT 162.800 147.000 163.600 147.200 ;
        RECT 169.200 146.400 170.000 149.200 ;
        RECT 175.000 148.600 178.800 149.400 ;
        RECT 175.000 147.400 175.800 148.600 ;
        RECT 179.400 148.000 180.000 150.000 ;
        RECT 162.800 146.200 163.600 146.400 ;
        RECT 153.000 145.400 155.600 146.200 ;
        RECT 159.000 145.600 163.600 146.200 ;
        RECT 164.400 145.600 166.000 146.400 ;
        RECT 169.000 145.600 170.000 146.400 ;
        RECT 174.000 146.800 175.800 147.400 ;
        RECT 178.800 147.400 180.000 148.000 ;
        RECT 180.600 148.300 181.400 151.200 ;
        RECT 185.200 148.800 186.000 150.400 ;
        RECT 186.600 148.400 187.200 151.800 ;
        RECT 188.400 151.600 189.200 151.800 ;
        RECT 183.600 148.300 184.400 148.400 ;
        RECT 180.600 148.200 184.400 148.300 ;
        RECT 186.600 148.300 189.200 148.400 ;
        RECT 190.000 148.300 190.800 148.400 ;
        RECT 180.600 147.700 185.200 148.200 ;
        RECT 174.000 146.200 174.800 146.800 ;
        RECT 154.800 142.200 155.600 145.400 ;
        RECT 172.400 145.400 174.800 146.200 ;
        RECT 156.400 142.200 157.200 145.000 ;
        RECT 158.000 142.200 158.800 145.000 ;
        RECT 159.600 142.200 160.400 145.000 ;
        RECT 162.800 142.200 163.600 145.000 ;
        RECT 166.000 142.200 166.800 145.000 ;
        RECT 167.600 142.200 168.400 145.000 ;
        RECT 169.200 142.200 170.000 145.000 ;
        RECT 170.800 142.200 171.600 145.000 ;
        RECT 172.400 142.200 173.200 145.400 ;
        RECT 178.800 142.200 179.600 147.400 ;
        RECT 180.600 146.800 181.400 147.700 ;
        RECT 183.600 147.600 185.200 147.700 ;
        RECT 186.600 147.700 190.800 148.300 ;
        RECT 186.600 147.600 189.200 147.700 ;
        RECT 184.400 147.200 185.200 147.600 ;
        RECT 180.400 146.000 181.400 146.800 ;
        RECT 183.800 146.200 187.400 146.600 ;
        RECT 188.400 146.200 189.000 147.600 ;
        RECT 190.000 146.800 190.800 147.700 ;
        RECT 191.600 146.200 192.400 153.700 ;
        RECT 193.200 151.600 194.000 153.200 ;
        RECT 194.800 151.800 195.600 159.800 ;
        RECT 196.400 152.400 197.200 159.800 ;
        RECT 199.600 152.400 200.400 159.800 ;
        RECT 196.400 151.800 200.400 152.400 ;
        RECT 195.000 150.400 195.600 151.800 ;
        RECT 198.800 150.400 199.600 150.800 ;
        RECT 194.800 149.800 197.200 150.400 ;
        RECT 198.800 149.800 200.400 150.400 ;
        RECT 194.800 149.600 195.600 149.800 ;
        RECT 193.200 148.300 194.000 148.400 ;
        RECT 196.600 148.300 197.200 149.800 ;
        RECT 199.600 149.600 200.400 149.800 ;
        RECT 193.200 147.700 197.200 148.300 ;
        RECT 193.200 147.600 194.000 147.700 ;
        RECT 183.600 146.000 187.600 146.200 ;
        RECT 180.400 142.200 181.200 146.000 ;
        RECT 183.600 142.200 184.400 146.000 ;
        RECT 186.800 142.200 187.600 146.000 ;
        RECT 188.400 142.200 189.200 146.200 ;
        RECT 191.600 145.600 193.400 146.200 ;
        RECT 194.800 145.600 195.600 146.400 ;
        RECT 196.600 146.200 197.200 147.700 ;
        RECT 198.000 148.300 198.800 149.200 ;
        RECT 202.800 148.300 203.600 159.800 ;
        RECT 205.000 152.600 205.800 159.800 ;
        RECT 210.800 155.800 211.600 159.800 ;
        RECT 205.000 151.800 206.800 152.600 ;
        RECT 204.400 149.600 205.200 151.200 ;
        RECT 198.000 147.700 203.600 148.300 ;
        RECT 198.000 147.600 198.800 147.700 ;
        RECT 192.600 142.200 193.400 145.600 ;
        RECT 195.000 144.800 195.800 145.600 ;
        RECT 196.400 142.200 197.200 146.200 ;
        RECT 201.200 144.800 202.000 146.400 ;
        RECT 202.800 142.200 203.600 147.700 ;
        RECT 206.000 148.400 206.600 151.800 ;
        RECT 211.000 151.600 211.600 155.800 ;
        RECT 214.000 151.800 214.800 159.800 ;
        RECT 218.200 152.400 219.000 159.800 ;
        RECT 223.600 156.400 224.400 159.800 ;
        RECT 223.400 155.800 224.400 156.400 ;
        RECT 223.400 155.200 224.000 155.800 ;
        RECT 226.800 155.200 227.600 159.800 ;
        RECT 230.000 157.000 230.800 159.800 ;
        RECT 231.600 157.000 232.400 159.800 ;
        RECT 222.000 154.600 224.000 155.200 ;
        RECT 219.600 153.600 220.400 154.400 ;
        RECT 219.800 152.400 220.400 153.600 ;
        RECT 218.200 151.800 219.200 152.400 ;
        RECT 219.800 151.800 221.200 152.400 ;
        RECT 211.000 151.000 213.400 151.600 ;
        RECT 210.800 149.600 211.600 150.400 ;
        RECT 206.000 147.600 206.800 148.400 ;
        RECT 207.600 148.300 208.400 148.400 ;
        RECT 209.200 148.300 210.000 149.200 ;
        RECT 207.600 147.700 210.000 148.300 ;
        RECT 211.000 148.800 211.600 149.600 ;
        RECT 211.000 148.200 212.000 148.800 ;
        RECT 211.200 148.000 212.000 148.200 ;
        RECT 207.600 147.600 208.400 147.700 ;
        RECT 209.200 147.600 210.000 147.700 ;
        RECT 212.800 147.600 213.400 151.000 ;
        RECT 214.200 150.400 214.800 151.800 ;
        RECT 218.600 150.400 219.200 151.800 ;
        RECT 220.400 151.600 221.200 151.800 ;
        RECT 214.000 150.300 214.800 150.400 ;
        RECT 217.200 150.300 218.000 150.400 ;
        RECT 214.000 149.700 218.000 150.300 ;
        RECT 214.000 149.600 214.800 149.700 ;
        RECT 206.000 144.200 206.600 147.600 ;
        RECT 212.800 147.400 213.600 147.600 ;
        RECT 210.600 147.000 213.600 147.400 ;
        RECT 209.400 146.800 213.600 147.000 ;
        RECT 209.400 146.400 211.200 146.800 ;
        RECT 207.600 144.800 208.400 146.400 ;
        RECT 209.400 146.200 210.000 146.400 ;
        RECT 214.200 146.200 214.800 149.600 ;
        RECT 217.200 148.800 218.000 149.700 ;
        RECT 218.600 149.600 219.600 150.400 ;
        RECT 218.600 148.400 219.200 149.600 ;
        RECT 222.000 149.000 222.800 154.600 ;
        RECT 224.600 154.400 228.800 155.200 ;
        RECT 233.200 155.000 234.000 159.800 ;
        RECT 236.400 155.000 237.200 159.800 ;
        RECT 224.600 154.000 225.200 154.400 ;
        RECT 223.600 153.200 225.200 154.000 ;
        RECT 228.200 153.800 234.000 154.400 ;
        RECT 226.200 153.200 227.600 153.800 ;
        RECT 226.200 153.000 232.400 153.200 ;
        RECT 227.000 152.600 232.400 153.000 ;
        RECT 231.600 152.400 232.400 152.600 ;
        RECT 233.400 153.000 234.000 153.800 ;
        RECT 234.600 153.600 237.200 154.400 ;
        RECT 239.600 153.600 240.400 159.800 ;
        RECT 241.200 157.000 242.000 159.800 ;
        RECT 242.800 157.000 243.600 159.800 ;
        RECT 244.400 157.000 245.200 159.800 ;
        RECT 242.800 154.400 247.000 155.200 ;
        RECT 247.600 154.400 248.400 159.800 ;
        RECT 250.800 155.200 251.600 159.800 ;
        RECT 250.800 154.600 253.400 155.200 ;
        RECT 247.600 153.600 250.200 154.400 ;
        RECT 241.200 153.000 242.000 153.200 ;
        RECT 233.400 152.400 242.000 153.000 ;
        RECT 244.400 153.000 245.200 153.200 ;
        RECT 252.800 153.000 253.400 154.600 ;
        RECT 244.400 152.400 253.400 153.000 ;
        RECT 252.800 150.600 253.400 152.400 ;
        RECT 254.000 152.000 254.800 159.800 ;
        RECT 255.600 152.300 256.400 152.400 ;
        RECT 257.200 152.300 258.000 153.200 ;
        RECT 254.000 151.200 255.000 152.000 ;
        RECT 255.600 151.700 258.000 152.300 ;
        RECT 255.600 151.600 256.400 151.700 ;
        RECT 257.200 151.600 258.000 151.700 ;
        RECT 223.400 150.000 246.800 150.600 ;
        RECT 252.800 150.000 253.600 150.600 ;
        RECT 223.400 149.800 224.200 150.000 ;
        RECT 225.200 149.600 226.000 150.000 ;
        RECT 228.400 149.600 229.200 150.000 ;
        RECT 246.000 149.400 246.800 150.000 ;
        RECT 215.600 148.200 216.400 148.400 ;
        RECT 215.600 147.600 217.200 148.200 ;
        RECT 218.600 147.600 221.200 148.400 ;
        RECT 222.000 148.200 230.800 149.000 ;
        RECT 231.400 148.600 233.400 149.400 ;
        RECT 237.200 148.600 240.400 149.400 ;
        RECT 216.400 147.200 217.200 147.600 ;
        RECT 215.800 146.200 219.400 146.600 ;
        RECT 220.400 146.200 221.000 147.600 ;
        RECT 206.000 142.200 206.800 144.200 ;
        RECT 209.200 142.200 210.000 146.200 ;
        RECT 213.400 145.200 214.800 146.200 ;
        RECT 215.600 146.000 219.600 146.200 ;
        RECT 213.400 142.200 214.200 145.200 ;
        RECT 215.600 142.200 216.400 146.000 ;
        RECT 218.800 142.200 219.600 146.000 ;
        RECT 220.400 142.200 221.200 146.200 ;
        RECT 222.000 142.200 222.800 148.200 ;
        RECT 224.400 146.800 227.400 147.600 ;
        RECT 226.600 146.200 227.400 146.800 ;
        RECT 232.600 146.200 233.400 148.600 ;
        RECT 234.800 146.800 235.600 148.400 ;
        RECT 240.000 147.800 240.800 148.000 ;
        RECT 236.400 147.200 240.800 147.800 ;
        RECT 236.400 147.000 237.200 147.200 ;
        RECT 242.800 146.400 243.600 149.200 ;
        RECT 248.600 148.600 252.400 149.400 ;
        RECT 248.600 147.400 249.400 148.600 ;
        RECT 253.000 148.000 253.600 150.000 ;
        RECT 236.400 146.200 237.200 146.400 ;
        RECT 226.600 145.400 229.200 146.200 ;
        RECT 232.600 145.600 237.200 146.200 ;
        RECT 238.000 145.600 239.600 146.400 ;
        RECT 242.600 145.600 243.600 146.400 ;
        RECT 247.600 146.800 249.400 147.400 ;
        RECT 252.400 147.400 253.600 148.000 ;
        RECT 247.600 146.200 248.400 146.800 ;
        RECT 228.400 142.200 229.200 145.400 ;
        RECT 246.000 145.400 248.400 146.200 ;
        RECT 230.000 142.200 230.800 145.000 ;
        RECT 231.600 142.200 232.400 145.000 ;
        RECT 233.200 142.200 234.000 145.000 ;
        RECT 236.400 142.200 237.200 145.000 ;
        RECT 239.600 142.200 240.400 145.000 ;
        RECT 241.200 142.200 242.000 145.000 ;
        RECT 242.800 142.200 243.600 145.000 ;
        RECT 244.400 142.200 245.200 145.000 ;
        RECT 246.000 142.200 246.800 145.400 ;
        RECT 252.400 142.200 253.200 147.400 ;
        RECT 254.200 146.800 255.000 151.200 ;
        RECT 254.000 146.000 255.000 146.800 ;
        RECT 258.800 146.200 259.600 159.800 ;
        RECT 262.000 151.800 262.800 159.800 ;
        RECT 263.600 152.400 264.400 159.800 ;
        RECT 266.800 152.400 267.600 159.800 ;
        RECT 270.000 155.800 270.800 159.800 ;
        RECT 270.200 155.600 270.800 155.800 ;
        RECT 273.200 155.800 274.000 159.800 ;
        RECT 282.800 155.800 283.600 159.800 ;
        RECT 273.200 155.600 273.800 155.800 ;
        RECT 270.200 155.000 273.800 155.600 ;
        RECT 271.600 152.800 272.400 154.400 ;
        RECT 273.200 152.400 273.800 155.000 ;
        RECT 263.600 151.800 267.600 152.400 ;
        RECT 262.200 150.400 262.800 151.800 ;
        RECT 268.400 150.800 269.200 152.400 ;
        RECT 273.200 151.600 274.000 152.400 ;
        RECT 283.000 151.600 283.600 155.800 ;
        RECT 286.000 152.300 286.800 159.800 ;
        RECT 288.400 153.600 289.200 154.400 ;
        RECT 288.400 152.400 289.000 153.600 ;
        RECT 289.800 152.400 290.600 159.800 ;
        RECT 287.600 152.300 289.000 152.400 ;
        RECT 286.000 151.800 289.000 152.300 ;
        RECT 289.600 151.800 290.600 152.400 ;
        RECT 295.600 152.000 296.400 159.800 ;
        RECT 298.800 155.200 299.600 159.800 ;
        RECT 286.100 151.700 288.400 151.800 ;
        RECT 266.000 150.400 266.800 150.800 ;
        RECT 262.000 149.800 264.400 150.400 ;
        RECT 266.000 149.800 267.600 150.400 ;
        RECT 262.000 149.600 262.800 149.800 ;
        RECT 260.400 146.800 261.200 148.400 ;
        RECT 262.000 148.300 262.800 148.400 ;
        RECT 263.800 148.300 264.400 149.800 ;
        RECT 266.800 149.600 267.600 149.800 ;
        RECT 270.000 149.600 271.600 150.400 ;
        RECT 262.000 147.700 264.400 148.300 ;
        RECT 262.000 147.600 262.800 147.700 ;
        RECT 254.000 142.200 254.800 146.000 ;
        RECT 257.800 145.600 259.600 146.200 ;
        RECT 262.000 145.600 262.800 146.400 ;
        RECT 263.800 146.200 264.400 147.700 ;
        RECT 265.200 147.600 266.000 149.200 ;
        RECT 273.200 148.400 273.800 151.600 ;
        RECT 283.000 151.000 285.400 151.600 ;
        RECT 282.800 149.600 283.600 150.400 ;
        RECT 272.200 148.200 273.800 148.400 ;
        RECT 272.000 147.800 273.800 148.200 ;
        RECT 279.600 148.300 280.400 148.400 ;
        RECT 281.200 148.300 282.000 149.200 ;
        RECT 283.000 148.800 283.600 149.600 ;
        RECT 257.800 142.200 258.600 145.600 ;
        RECT 262.200 144.800 263.000 145.600 ;
        RECT 263.600 142.200 264.400 146.200 ;
        RECT 272.000 142.200 272.800 147.800 ;
        RECT 279.600 147.700 282.000 148.300 ;
        RECT 282.800 148.000 284.000 148.800 ;
        RECT 279.600 147.600 280.400 147.700 ;
        RECT 281.200 147.600 282.000 147.700 ;
        RECT 284.800 147.600 285.400 151.000 ;
        RECT 286.200 150.400 286.800 151.700 ;
        RECT 287.600 151.600 288.400 151.700 ;
        RECT 286.000 149.600 286.800 150.400 ;
        RECT 284.800 147.400 285.600 147.600 ;
        RECT 282.600 147.000 285.600 147.400 ;
        RECT 281.400 146.800 285.600 147.000 ;
        RECT 281.400 146.400 283.200 146.800 ;
        RECT 281.400 146.200 282.000 146.400 ;
        RECT 286.200 146.200 286.800 149.600 ;
        RECT 289.600 148.400 290.200 151.800 ;
        RECT 295.400 151.200 296.400 152.000 ;
        RECT 297.000 154.600 299.600 155.200 ;
        RECT 297.000 153.000 297.600 154.600 ;
        RECT 302.000 154.400 302.800 159.800 ;
        RECT 305.200 157.000 306.000 159.800 ;
        RECT 306.800 157.000 307.600 159.800 ;
        RECT 308.400 157.000 309.200 159.800 ;
        RECT 303.400 154.400 307.600 155.200 ;
        RECT 300.200 153.600 302.800 154.400 ;
        RECT 310.000 153.600 310.800 159.800 ;
        RECT 313.200 155.000 314.000 159.800 ;
        RECT 316.400 155.000 317.200 159.800 ;
        RECT 318.000 157.000 318.800 159.800 ;
        RECT 319.600 157.000 320.400 159.800 ;
        RECT 322.800 155.200 323.600 159.800 ;
        RECT 326.000 156.400 326.800 159.800 ;
        RECT 326.000 155.800 327.000 156.400 ;
        RECT 326.400 155.200 327.000 155.800 ;
        RECT 321.600 154.400 325.800 155.200 ;
        RECT 326.400 154.600 328.400 155.200 ;
        RECT 313.200 153.600 315.800 154.400 ;
        RECT 316.400 153.800 322.200 154.400 ;
        RECT 325.200 154.000 325.800 154.400 ;
        RECT 305.200 153.000 306.000 153.200 ;
        RECT 297.000 152.400 306.000 153.000 ;
        RECT 308.400 153.000 309.200 153.200 ;
        RECT 316.400 153.000 317.000 153.800 ;
        RECT 322.800 153.200 324.200 153.800 ;
        RECT 325.200 153.200 326.800 154.000 ;
        RECT 308.400 152.400 317.000 153.000 ;
        RECT 318.000 153.000 324.200 153.200 ;
        RECT 318.000 152.600 323.400 153.000 ;
        RECT 318.000 152.400 318.800 152.600 ;
        RECT 290.800 148.800 291.600 150.400 ;
        RECT 287.600 147.600 290.200 148.400 ;
        RECT 292.400 148.300 293.200 148.400 ;
        RECT 295.400 148.300 296.200 151.200 ;
        RECT 297.000 150.600 297.600 152.400 ;
        RECT 324.400 152.300 325.200 152.400 ;
        RECT 326.000 152.300 326.800 152.400 ;
        RECT 321.000 151.800 322.000 152.000 ;
        RECT 324.400 151.800 326.800 152.300 ;
        RECT 298.200 151.700 326.800 151.800 ;
        RECT 298.200 151.200 325.200 151.700 ;
        RECT 326.000 151.600 326.800 151.700 ;
        RECT 298.200 151.000 299.000 151.200 ;
        RECT 292.400 148.200 296.200 148.300 ;
        RECT 291.600 147.700 296.200 148.200 ;
        RECT 291.600 147.600 293.200 147.700 ;
        RECT 287.800 146.200 288.400 147.600 ;
        RECT 291.600 147.200 292.400 147.600 ;
        RECT 295.400 146.800 296.200 147.700 ;
        RECT 296.800 150.000 297.600 150.600 ;
        RECT 296.800 148.000 297.400 150.000 ;
        RECT 298.000 148.600 301.800 149.400 ;
        RECT 296.800 147.400 298.000 148.000 ;
        RECT 289.400 146.200 293.000 146.600 ;
        RECT 281.200 142.200 282.000 146.200 ;
        RECT 285.400 145.200 286.800 146.200 ;
        RECT 285.400 142.200 286.200 145.200 ;
        RECT 287.600 142.200 288.400 146.200 ;
        RECT 289.200 146.000 293.200 146.200 ;
        RECT 295.400 146.000 296.400 146.800 ;
        RECT 289.200 142.200 290.000 146.000 ;
        RECT 292.400 142.200 293.200 146.000 ;
        RECT 295.600 142.200 296.400 146.000 ;
        RECT 297.200 142.200 298.000 147.400 ;
        RECT 301.000 147.400 301.800 148.600 ;
        RECT 301.000 146.800 302.800 147.400 ;
        RECT 302.000 146.200 302.800 146.800 ;
        RECT 306.800 146.400 307.600 149.200 ;
        RECT 310.000 148.600 313.200 149.400 ;
        RECT 317.000 148.600 319.000 149.400 ;
        RECT 327.600 149.000 328.400 154.600 ;
        RECT 330.000 153.600 330.800 154.400 ;
        RECT 330.000 152.400 330.600 153.600 ;
        RECT 331.400 152.400 332.200 159.800 ;
        RECT 329.200 151.800 330.600 152.400 ;
        RECT 331.200 151.800 332.200 152.400 ;
        RECT 329.200 151.600 330.000 151.800 ;
        RECT 309.600 147.800 310.400 148.000 ;
        RECT 309.600 147.200 314.000 147.800 ;
        RECT 313.200 147.000 314.000 147.200 ;
        RECT 314.800 146.800 315.600 148.400 ;
        RECT 302.000 145.400 304.400 146.200 ;
        RECT 306.800 145.600 307.800 146.400 ;
        RECT 310.800 145.600 312.400 146.400 ;
        RECT 313.200 146.200 314.000 146.400 ;
        RECT 317.000 146.200 317.800 148.600 ;
        RECT 319.600 148.200 328.400 149.000 ;
        RECT 331.200 148.400 331.800 151.800 ;
        RECT 332.400 148.800 333.200 150.400 ;
        RECT 323.000 146.800 326.000 147.600 ;
        RECT 323.000 146.200 323.800 146.800 ;
        RECT 313.200 145.600 317.800 146.200 ;
        RECT 303.600 142.200 304.400 145.400 ;
        RECT 321.200 145.400 323.800 146.200 ;
        RECT 305.200 142.200 306.000 145.000 ;
        RECT 306.800 142.200 307.600 145.000 ;
        RECT 308.400 142.200 309.200 145.000 ;
        RECT 310.000 142.200 310.800 145.000 ;
        RECT 313.200 142.200 314.000 145.000 ;
        RECT 316.400 142.200 317.200 145.000 ;
        RECT 318.000 142.200 318.800 145.000 ;
        RECT 319.600 142.200 320.400 145.000 ;
        RECT 321.200 142.200 322.000 145.400 ;
        RECT 327.600 142.200 328.400 148.200 ;
        RECT 329.200 147.600 331.800 148.400 ;
        RECT 334.000 148.300 334.800 148.400 ;
        RECT 335.600 148.300 336.400 159.800 ;
        RECT 339.600 153.600 340.400 154.400 ;
        RECT 339.600 152.400 340.200 153.600 ;
        RECT 341.000 152.400 341.800 159.800 ;
        RECT 346.000 153.600 346.800 154.400 ;
        RECT 346.000 152.400 346.600 153.600 ;
        RECT 347.400 152.400 348.200 159.800 ;
        RECT 353.800 158.400 354.600 159.800 ;
        RECT 353.800 157.600 355.600 158.400 ;
        RECT 352.400 153.600 353.200 154.400 ;
        RECT 352.400 152.400 353.000 153.600 ;
        RECT 353.800 152.400 354.600 157.600 ;
        RECT 338.800 151.800 340.200 152.400 ;
        RECT 340.800 151.800 341.800 152.400 ;
        RECT 345.200 151.800 346.600 152.400 ;
        RECT 347.200 151.800 348.200 152.400 ;
        RECT 351.600 151.800 353.000 152.400 ;
        RECT 353.600 151.800 354.600 152.400 ;
        RECT 360.600 152.400 361.400 159.800 ;
        RECT 362.000 153.600 362.800 154.400 ;
        RECT 362.200 152.400 362.800 153.600 ;
        RECT 360.600 151.800 361.600 152.400 ;
        RECT 362.200 151.800 363.600 152.400 ;
        RECT 338.800 151.600 339.600 151.800 ;
        RECT 340.800 150.400 341.400 151.800 ;
        RECT 345.200 151.600 346.000 151.800 ;
        RECT 347.200 150.400 347.800 151.800 ;
        RECT 351.600 151.600 352.400 151.800 ;
        RECT 340.400 149.600 341.400 150.400 ;
        RECT 346.800 149.600 347.800 150.400 ;
        RECT 340.800 148.400 341.400 149.600 ;
        RECT 347.200 148.400 347.800 149.600 ;
        RECT 353.600 148.400 354.200 151.800 ;
        RECT 361.000 150.400 361.600 151.800 ;
        RECT 362.800 151.600 363.600 151.800 ;
        RECT 361.000 149.600 362.000 150.400 ;
        RECT 366.000 150.300 366.800 159.800 ;
        RECT 369.200 159.200 373.200 159.800 ;
        RECT 367.600 151.600 368.400 153.200 ;
        RECT 369.200 151.800 370.000 159.200 ;
        RECT 370.800 151.800 371.600 158.600 ;
        RECT 372.400 152.400 373.200 159.200 ;
        RECT 375.600 152.400 376.400 159.800 ;
        RECT 381.000 152.800 381.800 159.800 ;
        RECT 385.200 155.000 386.000 159.000 ;
        RECT 372.400 151.800 376.400 152.400 ;
        RECT 380.200 152.200 381.800 152.800 ;
        RECT 371.000 151.200 371.600 151.800 ;
        RECT 367.600 150.300 368.400 150.400 ;
        RECT 366.000 149.700 368.400 150.300 ;
        RECT 361.000 148.400 361.600 149.600 ;
        RECT 334.000 148.200 336.400 148.300 ;
        RECT 333.200 147.700 336.400 148.200 ;
        RECT 333.200 147.600 334.800 147.700 ;
        RECT 329.400 146.200 330.000 147.600 ;
        RECT 333.200 147.200 334.000 147.600 ;
        RECT 331.000 146.200 334.600 146.600 ;
        RECT 329.200 142.200 330.000 146.200 ;
        RECT 330.800 146.000 334.800 146.200 ;
        RECT 330.800 142.200 331.600 146.000 ;
        RECT 334.000 142.200 334.800 146.000 ;
        RECT 335.600 142.200 336.400 147.700 ;
        RECT 338.800 147.600 341.400 148.400 ;
        RECT 343.600 148.200 344.400 148.400 ;
        RECT 342.800 147.600 344.400 148.200 ;
        RECT 345.200 147.600 347.800 148.400 ;
        RECT 350.000 148.200 350.800 148.400 ;
        RECT 349.200 147.600 350.800 148.200 ;
        RECT 351.600 147.600 354.200 148.400 ;
        RECT 356.400 148.300 357.200 148.400 ;
        RECT 358.000 148.300 358.800 148.400 ;
        RECT 356.400 148.200 358.800 148.300 ;
        RECT 355.600 147.700 359.600 148.200 ;
        RECT 355.600 147.600 357.200 147.700 ;
        RECT 358.000 147.600 359.600 147.700 ;
        RECT 361.000 147.600 363.600 148.400 ;
        RECT 337.200 144.800 338.000 146.400 ;
        RECT 339.000 146.200 339.600 147.600 ;
        RECT 342.800 147.200 343.600 147.600 ;
        RECT 340.600 146.200 344.200 146.600 ;
        RECT 345.400 146.200 346.000 147.600 ;
        RECT 349.200 147.200 350.000 147.600 ;
        RECT 347.000 146.200 350.600 146.600 ;
        RECT 351.800 146.200 352.400 147.600 ;
        RECT 355.600 147.200 356.400 147.600 ;
        RECT 358.800 147.200 359.600 147.600 ;
        RECT 353.400 146.200 357.000 146.600 ;
        RECT 358.200 146.200 361.800 146.600 ;
        RECT 362.800 146.200 363.400 147.600 ;
        RECT 366.000 146.200 366.800 149.700 ;
        RECT 367.600 149.600 368.400 149.700 ;
        RECT 369.200 149.600 370.000 151.200 ;
        RECT 371.000 150.600 373.000 151.200 ;
        RECT 372.400 150.400 373.000 150.600 ;
        RECT 374.800 150.400 375.600 150.800 ;
        RECT 372.400 149.600 373.200 150.400 ;
        RECT 374.800 149.800 376.400 150.400 ;
        RECT 375.600 149.600 376.400 149.800 ;
        RECT 378.800 149.600 379.600 151.200 ;
        RECT 371.000 148.800 371.800 149.600 ;
        RECT 371.000 148.400 371.600 148.800 ;
        RECT 370.800 147.600 371.600 148.400 ;
        RECT 372.400 146.200 373.000 149.600 ;
        RECT 374.000 147.600 374.800 149.200 ;
        RECT 380.200 148.400 380.800 152.200 ;
        RECT 385.400 151.600 386.000 155.000 ;
        RECT 382.200 151.000 386.000 151.600 ;
        RECT 382.200 149.000 382.800 151.000 ;
        RECT 377.200 148.300 378.000 148.400 ;
        RECT 378.800 148.300 380.800 148.400 ;
        RECT 377.200 147.700 380.800 148.300 ;
        RECT 381.400 148.200 382.800 149.000 ;
        RECT 383.600 148.800 384.400 150.400 ;
        RECT 385.200 148.800 386.000 150.400 ;
        RECT 377.200 147.600 378.000 147.700 ;
        RECT 378.800 147.600 380.800 147.700 ;
        RECT 380.200 147.000 380.800 147.600 ;
        RECT 381.800 147.800 382.800 148.200 ;
        RECT 381.800 147.200 386.000 147.800 ;
        RECT 380.200 146.600 381.000 147.000 ;
        RECT 338.800 142.200 339.600 146.200 ;
        RECT 340.400 146.000 344.400 146.200 ;
        RECT 340.400 142.200 341.200 146.000 ;
        RECT 343.600 142.200 344.400 146.000 ;
        RECT 345.200 142.200 346.000 146.200 ;
        RECT 346.800 146.000 350.800 146.200 ;
        RECT 346.800 142.200 347.600 146.000 ;
        RECT 350.000 142.200 350.800 146.000 ;
        RECT 351.600 142.200 352.400 146.200 ;
        RECT 353.200 146.000 357.200 146.200 ;
        RECT 353.200 142.200 354.000 146.000 ;
        RECT 356.400 142.200 357.200 146.000 ;
        RECT 358.000 146.000 362.000 146.200 ;
        RECT 358.000 142.200 358.800 146.000 ;
        RECT 361.200 142.200 362.000 146.000 ;
        RECT 362.800 142.200 363.600 146.200 ;
        RECT 366.000 145.600 367.800 146.200 ;
        RECT 367.000 142.200 367.800 145.600 ;
        RECT 371.800 142.200 373.400 146.200 ;
        RECT 380.200 146.000 381.800 146.600 ;
        RECT 381.000 143.000 381.800 146.000 ;
        RECT 385.400 145.000 386.000 147.200 ;
        RECT 385.200 143.000 386.000 145.000 ;
        RECT 386.800 142.200 387.600 159.800 ;
        RECT 388.400 152.300 389.200 152.400 ;
        RECT 390.000 152.300 390.800 159.800 ;
        RECT 388.400 151.800 390.800 152.300 ;
        RECT 393.200 155.800 394.000 159.800 ;
        RECT 396.400 155.800 397.200 159.800 ;
        RECT 388.400 151.700 390.700 151.800 ;
        RECT 388.400 151.600 389.200 151.700 ;
        RECT 390.000 150.400 390.600 151.700 ;
        RECT 393.200 151.600 393.800 155.800 ;
        RECT 396.600 155.600 397.200 155.800 ;
        RECT 399.600 155.800 400.400 159.800 ;
        RECT 402.800 155.800 403.600 159.800 ;
        RECT 399.600 155.600 400.200 155.800 ;
        RECT 396.600 155.000 400.200 155.600 ;
        RECT 403.000 155.600 403.600 155.800 ;
        RECT 406.000 155.800 406.800 159.800 ;
        RECT 406.000 155.600 406.600 155.800 ;
        RECT 403.000 155.000 406.600 155.600 ;
        RECT 396.600 152.400 397.200 155.000 ;
        RECT 398.000 152.800 398.800 154.400 ;
        RECT 403.000 152.400 403.600 155.000 ;
        RECT 404.400 152.800 405.200 154.400 ;
        RECT 410.000 153.600 410.800 154.400 ;
        RECT 410.000 152.400 410.600 153.600 ;
        RECT 411.400 152.400 412.200 159.800 ;
        RECT 396.400 151.600 397.200 152.400 ;
        RECT 391.400 151.000 393.800 151.600 ;
        RECT 390.000 149.600 390.800 150.400 ;
        RECT 388.400 144.800 389.200 146.400 ;
        RECT 390.000 146.200 390.600 149.600 ;
        RECT 391.400 147.600 392.000 151.000 ;
        RECT 393.200 149.600 394.000 150.400 ;
        RECT 393.200 148.800 393.800 149.600 ;
        RECT 392.800 148.200 393.800 148.800 ;
        RECT 392.800 148.000 393.600 148.200 ;
        RECT 394.800 147.600 395.600 149.200 ;
        RECT 396.600 148.400 397.200 151.600 ;
        RECT 401.200 150.800 402.000 152.400 ;
        RECT 402.800 151.600 403.600 152.400 ;
        RECT 398.800 149.600 400.400 150.400 ;
        RECT 403.000 148.400 403.600 151.600 ;
        RECT 407.600 150.800 408.400 152.400 ;
        RECT 409.200 151.800 410.600 152.400 ;
        RECT 411.200 151.800 412.200 152.400 ;
        RECT 409.200 151.600 410.000 151.800 ;
        RECT 411.200 150.400 411.800 151.800 ;
        RECT 405.200 149.600 406.800 150.400 ;
        RECT 410.800 149.600 411.800 150.400 ;
        RECT 411.200 148.400 411.800 149.600 ;
        RECT 412.400 148.800 413.200 150.400 ;
        RECT 396.600 148.200 398.200 148.400 ;
        RECT 403.000 148.200 404.600 148.400 ;
        RECT 396.600 147.800 398.400 148.200 ;
        RECT 403.000 147.800 404.800 148.200 ;
        RECT 391.200 147.400 392.000 147.600 ;
        RECT 391.200 147.000 394.200 147.400 ;
        RECT 391.200 146.800 395.400 147.000 ;
        RECT 393.600 146.400 395.400 146.800 ;
        RECT 394.800 146.200 395.400 146.400 ;
        RECT 390.000 145.200 391.400 146.200 ;
        RECT 390.600 142.200 391.400 145.200 ;
        RECT 394.800 142.200 395.600 146.200 ;
        RECT 397.600 142.200 398.400 147.800 ;
        RECT 404.000 144.400 404.800 147.800 ;
        RECT 409.200 147.600 411.800 148.400 ;
        RECT 414.000 148.300 414.800 148.400 ;
        RECT 417.200 148.300 418.000 159.800 ;
        RECT 418.800 155.000 419.600 159.000 ;
        RECT 418.800 151.600 419.400 155.000 ;
        RECT 423.000 152.800 423.800 159.800 ;
        RECT 423.000 152.200 424.600 152.800 ;
        RECT 423.600 151.600 424.600 152.200 ;
        RECT 418.800 151.000 422.600 151.600 ;
        RECT 418.800 148.800 419.600 150.400 ;
        RECT 420.400 148.800 421.200 150.400 ;
        RECT 422.000 149.000 422.600 151.000 ;
        RECT 414.000 148.200 418.000 148.300 ;
        RECT 413.200 147.700 418.000 148.200 ;
        RECT 422.000 148.200 423.400 149.000 ;
        RECT 424.000 148.400 424.600 151.600 ;
        RECT 434.800 151.400 435.600 159.800 ;
        RECT 439.200 156.400 440.000 159.800 ;
        RECT 438.000 155.800 440.000 156.400 ;
        RECT 443.600 155.800 444.400 159.800 ;
        RECT 447.800 155.800 449.000 159.800 ;
        RECT 438.000 155.000 438.800 155.800 ;
        RECT 443.600 155.200 444.200 155.800 ;
        RECT 441.400 154.600 445.000 155.200 ;
        RECT 447.600 155.000 448.400 155.800 ;
        RECT 441.400 154.400 442.200 154.600 ;
        RECT 444.200 154.400 445.000 154.600 ;
        RECT 438.000 153.000 438.800 153.200 ;
        RECT 442.600 153.000 443.400 153.200 ;
        RECT 438.000 152.400 443.400 153.000 ;
        RECT 444.000 153.000 446.200 153.600 ;
        RECT 444.000 151.800 444.600 153.000 ;
        RECT 445.400 152.800 446.200 153.000 ;
        RECT 447.800 153.200 449.200 154.000 ;
        RECT 447.800 152.200 448.400 153.200 ;
        RECT 439.800 151.400 444.600 151.800 ;
        RECT 434.800 151.200 444.600 151.400 ;
        RECT 446.000 151.600 448.400 152.200 ;
        RECT 425.200 149.600 426.000 151.200 ;
        RECT 434.800 151.000 440.600 151.200 ;
        RECT 434.800 150.800 440.400 151.000 ;
        RECT 441.200 150.300 442.000 150.400 ;
        RECT 444.400 150.300 445.200 150.400 ;
        RECT 441.200 150.200 445.200 150.300 ;
        RECT 437.000 149.700 445.200 150.200 ;
        RECT 437.000 149.600 442.000 149.700 ;
        RECT 444.400 149.600 445.200 149.700 ;
        RECT 437.000 149.400 437.800 149.600 ;
        RECT 438.600 148.400 439.400 148.600 ;
        RECT 446.000 148.400 446.600 151.600 ;
        RECT 452.400 151.200 453.200 159.800 ;
        RECT 454.000 155.800 454.800 159.800 ;
        RECT 454.200 155.600 454.800 155.800 ;
        RECT 457.200 155.800 458.000 159.800 ;
        RECT 462.000 155.800 462.800 159.800 ;
        RECT 457.200 155.600 457.800 155.800 ;
        RECT 454.200 155.000 457.800 155.600 ;
        RECT 462.200 155.600 462.800 155.800 ;
        RECT 465.200 155.800 466.000 159.800 ;
        RECT 465.200 155.600 465.800 155.800 ;
        RECT 462.200 155.000 465.800 155.600 ;
        RECT 454.200 152.400 454.800 155.000 ;
        RECT 455.600 152.800 456.400 154.400 ;
        RECT 457.200 154.300 458.000 154.400 ;
        RECT 463.600 154.300 464.400 154.400 ;
        RECT 457.200 153.700 464.400 154.300 ;
        RECT 457.200 153.600 458.000 153.700 ;
        RECT 463.600 152.800 464.400 153.700 ;
        RECT 454.000 151.600 454.800 152.400 ;
        RECT 449.000 150.600 453.200 151.200 ;
        RECT 449.000 150.400 449.800 150.600 ;
        RECT 450.600 149.800 451.400 150.000 ;
        RECT 447.600 149.200 451.400 149.800 ;
        RECT 447.600 149.000 448.400 149.200 ;
        RECT 422.000 147.800 423.000 148.200 ;
        RECT 413.200 147.600 414.800 147.700 ;
        RECT 409.400 146.200 410.000 147.600 ;
        RECT 413.200 147.200 414.000 147.600 ;
        RECT 411.000 146.200 414.600 146.600 ;
        RECT 404.000 143.600 405.200 144.400 ;
        RECT 404.000 142.200 404.800 143.600 ;
        RECT 409.200 142.200 410.000 146.200 ;
        RECT 410.800 146.000 414.800 146.200 ;
        RECT 410.800 142.200 411.600 146.000 ;
        RECT 414.000 142.200 414.800 146.000 ;
        RECT 415.600 144.800 416.400 146.400 ;
        RECT 417.200 142.200 418.000 147.700 ;
        RECT 418.800 147.200 423.000 147.800 ;
        RECT 424.000 147.600 426.000 148.400 ;
        RECT 426.800 148.300 427.600 148.400 ;
        RECT 435.600 148.300 446.600 148.400 ;
        RECT 426.800 147.800 446.600 148.300 ;
        RECT 426.800 147.700 437.200 147.800 ;
        RECT 426.800 147.600 427.600 147.700 ;
        RECT 435.600 147.600 437.200 147.700 ;
        RECT 418.800 145.000 419.400 147.200 ;
        RECT 424.000 147.000 424.600 147.600 ;
        RECT 423.800 146.600 424.600 147.000 ;
        RECT 423.000 146.000 424.600 146.600 ;
        RECT 418.800 143.000 419.600 145.000 ;
        RECT 423.000 143.000 423.800 146.000 ;
        RECT 434.800 142.200 435.600 147.000 ;
        RECT 439.800 145.600 440.400 147.800 ;
        RECT 445.400 147.600 446.200 147.800 ;
        RECT 452.400 147.200 453.200 150.600 ;
        RECT 454.200 148.400 454.800 151.600 ;
        RECT 465.200 152.400 465.800 155.000 ;
        RECT 466.800 153.800 467.600 159.800 ;
        RECT 467.000 153.200 467.600 153.800 ;
        RECT 470.000 159.200 474.000 159.800 ;
        RECT 470.000 153.800 470.800 159.200 ;
        RECT 471.600 153.800 472.400 158.600 ;
        RECT 473.200 154.000 474.000 159.200 ;
        RECT 475.000 159.200 478.600 159.800 ;
        RECT 475.000 159.000 475.600 159.200 ;
        RECT 470.000 153.200 470.600 153.800 ;
        RECT 467.000 152.600 470.600 153.200 ;
        RECT 471.800 153.400 472.400 153.800 ;
        RECT 474.800 153.400 475.600 159.000 ;
        RECT 478.000 159.000 478.600 159.200 ;
        RECT 471.800 153.000 475.600 153.400 ;
        RECT 476.400 153.000 477.200 158.600 ;
        RECT 478.000 153.000 478.800 159.000 ;
        RECT 471.800 152.800 475.400 153.000 ;
        RECT 476.400 152.400 477.000 153.000 ;
        RECT 483.400 152.800 484.200 159.800 ;
        RECT 487.600 155.000 488.400 159.000 ;
        RECT 465.200 151.600 466.000 152.400 ;
        RECT 476.400 152.200 477.200 152.400 ;
        RECT 473.800 151.600 477.200 152.200 ;
        RECT 482.600 152.200 484.200 152.800 ;
        RECT 456.400 149.600 458.000 150.400 ;
        RECT 465.200 148.400 465.800 151.600 ;
        RECT 471.600 149.600 473.200 150.400 ;
        RECT 454.200 148.200 455.800 148.400 ;
        RECT 464.200 148.200 465.800 148.400 ;
        RECT 454.200 147.800 456.000 148.200 ;
        RECT 449.400 146.600 453.200 147.200 ;
        RECT 449.400 146.400 450.200 146.600 ;
        RECT 438.000 144.200 438.800 145.000 ;
        RECT 439.600 144.800 440.400 145.600 ;
        RECT 441.400 145.400 442.200 145.600 ;
        RECT 441.400 144.800 444.200 145.400 ;
        RECT 443.600 144.200 444.200 144.800 ;
        RECT 447.600 144.200 448.400 145.000 ;
        RECT 438.000 143.600 440.000 144.200 ;
        RECT 439.200 142.200 440.000 143.600 ;
        RECT 443.600 142.200 444.400 144.200 ;
        RECT 447.600 143.600 449.000 144.200 ;
        RECT 447.800 142.200 449.000 143.600 ;
        RECT 452.400 142.200 453.200 146.600 ;
        RECT 455.200 146.400 456.000 147.800 ;
        RECT 454.000 145.600 456.000 146.400 ;
        RECT 455.200 142.200 456.000 145.600 ;
        RECT 464.000 147.800 465.800 148.200 ;
        RECT 464.000 142.200 464.800 147.800 ;
        RECT 473.800 145.000 474.400 151.600 ;
        RECT 481.200 149.600 482.000 151.200 ;
        RECT 482.600 148.400 483.200 152.200 ;
        RECT 487.800 151.600 488.400 155.000 ;
        RECT 484.600 151.000 488.400 151.600 ;
        RECT 484.600 149.000 485.200 151.000 ;
        RECT 481.200 147.600 483.200 148.400 ;
        RECT 483.800 148.200 485.200 149.000 ;
        RECT 486.000 148.800 486.800 150.400 ;
        RECT 487.600 148.800 488.400 150.400 ;
        RECT 482.600 147.000 483.200 147.600 ;
        RECT 484.200 147.800 485.200 148.200 ;
        RECT 484.200 147.200 488.400 147.800 ;
        RECT 482.600 146.600 483.400 147.000 ;
        RECT 482.600 146.000 484.200 146.600 ;
        RECT 470.400 144.400 474.400 145.000 ;
        RECT 483.400 144.400 484.200 146.000 ;
        RECT 487.800 145.000 488.400 147.200 ;
        RECT 470.000 143.600 471.000 144.400 ;
        RECT 473.200 144.200 474.400 144.400 ;
        RECT 470.000 142.200 470.800 143.600 ;
        RECT 473.200 142.200 474.000 144.200 ;
        RECT 482.800 143.600 484.200 144.400 ;
        RECT 483.400 143.000 484.200 143.600 ;
        RECT 487.600 143.000 488.400 145.000 ;
        RECT 489.200 142.200 490.000 159.800 ;
        RECT 495.000 158.400 497.000 159.800 ;
        RECT 495.000 157.600 498.000 158.400 ;
        RECT 495.000 151.800 497.000 157.600 ;
        RECT 504.200 152.800 505.000 159.800 ;
        RECT 508.400 155.000 509.200 159.000 ;
        RECT 503.400 152.200 505.000 152.800 ;
        RECT 492.400 147.600 493.200 149.200 ;
        RECT 494.000 148.800 494.800 150.400 ;
        RECT 495.800 148.400 496.400 151.800 ;
        RECT 497.200 148.800 498.000 150.400 ;
        RECT 502.000 149.600 502.800 151.200 ;
        RECT 503.400 148.400 504.000 152.200 ;
        RECT 508.600 151.600 509.200 155.000 ;
        RECT 505.400 151.000 509.200 151.600 ;
        RECT 505.400 149.000 506.000 151.000 ;
        RECT 495.600 148.200 496.400 148.400 ;
        RECT 498.800 148.200 499.600 148.400 ;
        RECT 494.000 147.600 496.400 148.200 ;
        RECT 498.000 147.600 499.600 148.200 ;
        RECT 502.000 147.600 504.000 148.400 ;
        RECT 504.600 148.200 506.000 149.000 ;
        RECT 506.800 148.800 507.600 150.400 ;
        RECT 508.400 148.800 509.200 150.400 ;
        RECT 490.800 144.800 491.600 146.400 ;
        RECT 494.000 146.200 494.600 147.600 ;
        RECT 498.000 147.200 498.800 147.600 ;
        RECT 503.400 147.000 504.000 147.600 ;
        RECT 505.000 147.800 506.000 148.200 ;
        RECT 505.000 147.200 509.200 147.800 ;
        RECT 503.400 146.600 504.200 147.000 ;
        RECT 495.800 146.200 499.400 146.600 ;
        RECT 492.400 142.800 493.200 146.200 ;
        RECT 494.000 143.400 494.800 146.200 ;
        RECT 495.600 146.000 499.600 146.200 ;
        RECT 503.400 146.000 505.000 146.600 ;
        RECT 495.600 142.800 496.400 146.000 ;
        RECT 492.400 142.200 496.400 142.800 ;
        RECT 498.800 142.200 499.600 146.000 ;
        RECT 504.200 144.400 505.000 146.000 ;
        RECT 508.600 145.000 509.200 147.200 ;
        RECT 503.600 143.600 505.000 144.400 ;
        RECT 504.200 143.000 505.000 143.600 ;
        RECT 508.400 143.000 509.200 145.000 ;
        RECT 510.000 142.200 510.800 159.800 ;
        RECT 511.600 154.300 512.400 154.400 ;
        RECT 513.200 154.300 514.000 159.800 ;
        RECT 511.600 153.700 514.000 154.300 ;
        RECT 511.600 153.600 512.400 153.700 ;
        RECT 511.600 144.800 512.400 146.400 ;
        RECT 513.200 142.200 514.000 153.700 ;
        RECT 516.400 155.000 517.200 159.000 ;
        RECT 520.600 158.400 521.400 159.800 ;
        RECT 520.600 157.600 522.000 158.400 ;
        RECT 516.400 151.600 517.000 155.000 ;
        RECT 520.600 152.800 521.400 157.600 ;
        RECT 520.600 152.200 522.200 152.800 ;
        RECT 516.400 151.000 520.200 151.600 ;
        RECT 516.400 148.800 517.200 150.400 ;
        RECT 518.000 148.800 518.800 150.400 ;
        RECT 519.600 149.000 520.200 151.000 ;
        RECT 519.600 148.200 521.000 149.000 ;
        RECT 521.600 148.400 522.200 152.200 ;
        RECT 526.000 151.400 526.800 159.800 ;
        RECT 530.400 156.400 531.200 159.800 ;
        RECT 529.200 155.800 531.200 156.400 ;
        RECT 534.800 155.800 535.600 159.800 ;
        RECT 539.000 155.800 540.200 159.800 ;
        RECT 529.200 155.000 530.000 155.800 ;
        RECT 534.800 155.200 535.400 155.800 ;
        RECT 532.600 154.600 536.200 155.200 ;
        RECT 538.800 155.000 539.600 155.800 ;
        RECT 532.600 154.400 533.400 154.600 ;
        RECT 535.400 154.400 536.200 154.600 ;
        RECT 529.200 153.000 530.000 153.200 ;
        RECT 533.800 153.000 534.600 153.200 ;
        RECT 529.200 152.400 534.600 153.000 ;
        RECT 535.200 153.000 537.400 153.600 ;
        RECT 535.200 151.800 535.800 153.000 ;
        RECT 536.600 152.800 537.400 153.000 ;
        RECT 539.000 153.200 540.400 154.000 ;
        RECT 539.000 152.200 539.600 153.200 ;
        RECT 531.000 151.400 535.800 151.800 ;
        RECT 526.000 151.200 535.800 151.400 ;
        RECT 537.200 151.600 539.600 152.200 ;
        RECT 522.800 150.300 523.600 151.200 ;
        RECT 526.000 151.000 531.800 151.200 ;
        RECT 526.000 150.800 531.600 151.000 ;
        RECT 524.400 150.300 525.200 150.400 ;
        RECT 522.800 149.700 525.200 150.300 ;
        RECT 532.400 150.200 533.200 150.400 ;
        RECT 522.800 149.600 523.600 149.700 ;
        RECT 524.400 149.600 525.200 149.700 ;
        RECT 528.200 149.600 533.200 150.200 ;
        RECT 528.200 149.400 529.000 149.600 ;
        RECT 530.800 149.400 531.600 149.600 ;
        RECT 529.800 148.400 530.600 148.600 ;
        RECT 537.200 148.400 537.800 151.600 ;
        RECT 543.600 151.200 544.400 159.800 ;
        RECT 545.200 152.400 546.000 159.800 ;
        RECT 545.200 151.800 547.400 152.400 ;
        RECT 540.200 150.600 544.400 151.200 ;
        RECT 540.200 150.400 541.000 150.600 ;
        RECT 541.800 149.800 542.600 150.000 ;
        RECT 538.800 149.200 542.600 149.800 ;
        RECT 538.800 149.000 539.600 149.200 ;
        RECT 519.600 147.800 520.600 148.200 ;
        RECT 516.400 147.200 520.600 147.800 ;
        RECT 521.600 147.600 523.600 148.400 ;
        RECT 526.800 147.800 537.800 148.400 ;
        RECT 526.800 147.600 528.400 147.800 ;
        RECT 514.800 144.800 515.600 146.400 ;
        RECT 516.400 145.000 517.000 147.200 ;
        RECT 521.600 147.000 522.200 147.600 ;
        RECT 521.400 146.600 522.200 147.000 ;
        RECT 520.600 146.000 522.200 146.600 ;
        RECT 516.400 143.000 517.200 145.000 ;
        RECT 520.600 143.000 521.400 146.000 ;
        RECT 526.000 142.200 526.800 147.000 ;
        RECT 531.000 145.600 531.600 147.800 ;
        RECT 532.400 147.600 533.200 147.800 ;
        RECT 536.600 147.600 537.400 147.800 ;
        RECT 543.600 147.200 544.400 150.600 ;
        RECT 546.800 151.200 547.400 151.800 ;
        RECT 546.800 150.400 548.000 151.200 ;
        RECT 545.200 148.800 546.000 150.400 ;
        RECT 546.800 147.400 547.400 150.400 ;
        RECT 540.600 146.600 544.400 147.200 ;
        RECT 540.600 146.400 541.400 146.600 ;
        RECT 529.200 144.200 530.000 145.000 ;
        RECT 530.800 144.800 531.600 145.600 ;
        RECT 532.600 145.400 533.400 145.600 ;
        RECT 532.600 144.800 535.400 145.400 ;
        RECT 534.800 144.200 535.400 144.800 ;
        RECT 538.800 144.200 539.600 145.000 ;
        RECT 529.200 143.600 531.200 144.200 ;
        RECT 530.400 142.200 531.200 143.600 ;
        RECT 534.800 142.200 535.600 144.200 ;
        RECT 538.800 143.600 540.200 144.200 ;
        RECT 539.000 142.200 540.200 143.600 ;
        RECT 543.600 142.200 544.400 146.600 ;
        RECT 545.200 146.800 547.400 147.400 ;
        RECT 545.200 142.200 546.000 146.800 ;
        RECT 1.200 122.200 2.000 139.800 ;
        RECT 4.400 135.600 5.200 137.200 ;
        RECT 2.800 133.600 3.600 135.200 ;
        RECT 6.000 122.200 6.800 139.800 ;
        RECT 8.200 136.400 9.000 139.800 ;
        RECT 14.000 137.800 14.800 139.800 ;
        RECT 8.200 135.800 10.000 136.400 ;
        RECT 7.600 128.800 8.400 130.400 ;
        RECT 9.200 122.200 10.000 135.800 ;
        RECT 12.400 135.600 13.200 137.200 ;
        RECT 10.800 134.300 11.600 135.200 ;
        RECT 12.500 134.300 13.100 135.600 ;
        RECT 14.200 134.400 14.800 137.800 ;
        RECT 17.200 136.000 18.000 139.800 ;
        RECT 20.400 136.000 21.200 139.800 ;
        RECT 17.200 135.800 21.200 136.000 ;
        RECT 22.000 135.800 22.800 139.800 ;
        RECT 17.400 135.400 21.000 135.800 ;
        RECT 18.000 134.400 18.800 134.800 ;
        RECT 22.000 134.400 22.600 135.800 ;
        RECT 10.800 133.700 13.100 134.300 ;
        RECT 14.000 134.300 14.800 134.400 ;
        RECT 17.200 134.300 18.800 134.400 ;
        RECT 14.000 133.800 18.800 134.300 ;
        RECT 14.000 133.700 18.000 133.800 ;
        RECT 10.800 133.600 11.600 133.700 ;
        RECT 14.000 133.600 14.800 133.700 ;
        RECT 17.200 133.600 18.000 133.700 ;
        RECT 20.200 133.600 22.800 134.400 ;
        RECT 24.800 134.200 25.600 139.800 ;
        RECT 31.200 134.200 32.000 139.800 ;
        RECT 36.400 136.000 37.200 139.800 ;
        RECT 39.600 136.000 40.400 139.800 ;
        RECT 36.400 135.800 40.400 136.000 ;
        RECT 41.200 135.800 42.000 139.800 ;
        RECT 36.600 135.400 40.200 135.800 ;
        RECT 37.200 134.400 38.000 134.800 ;
        RECT 41.200 134.400 41.800 135.800 ;
        RECT 23.800 133.800 25.600 134.200 ;
        RECT 30.200 133.800 32.000 134.200 ;
        RECT 36.400 133.800 38.000 134.400 ;
        RECT 23.800 133.600 25.400 133.800 ;
        RECT 30.200 133.600 31.800 133.800 ;
        RECT 36.400 133.600 37.200 133.800 ;
        RECT 39.400 133.600 42.000 134.400 ;
        RECT 44.000 134.200 44.800 139.800 ;
        RECT 50.800 136.000 51.600 139.800 ;
        RECT 43.000 133.800 44.800 134.200 ;
        RECT 50.600 135.200 51.600 136.000 ;
        RECT 43.000 133.600 44.600 133.800 ;
        RECT 14.200 130.200 14.800 133.600 ;
        RECT 15.600 130.800 16.400 132.400 ;
        RECT 18.800 131.600 19.600 133.200 ;
        RECT 20.200 130.200 20.800 133.600 ;
        RECT 23.800 130.400 24.400 133.600 ;
        RECT 26.000 131.600 27.600 132.400 ;
        RECT 22.000 130.200 22.800 130.400 ;
        RECT 14.000 129.400 15.800 130.200 ;
        RECT 15.000 122.200 15.800 129.400 ;
        RECT 19.800 129.600 20.800 130.200 ;
        RECT 21.400 129.600 22.800 130.200 ;
        RECT 23.600 129.600 24.400 130.400 ;
        RECT 28.400 129.600 29.200 131.200 ;
        RECT 30.200 130.400 30.800 133.600 ;
        RECT 32.400 131.600 34.000 132.400 ;
        RECT 38.000 131.600 38.800 133.200 ;
        RECT 30.000 129.600 30.800 130.400 ;
        RECT 34.800 129.600 35.600 131.200 ;
        RECT 39.400 130.200 40.000 133.600 ;
        RECT 43.000 130.400 43.600 133.600 ;
        RECT 45.200 131.600 46.800 132.400 ;
        RECT 41.200 130.200 42.000 130.400 ;
        RECT 39.000 129.600 40.000 130.200 ;
        RECT 40.600 129.600 42.000 130.200 ;
        RECT 42.800 129.600 43.600 130.400 ;
        RECT 47.600 129.600 48.400 131.200 ;
        RECT 50.600 130.800 51.400 135.200 ;
        RECT 52.400 134.600 53.200 139.800 ;
        RECT 58.800 136.600 59.600 139.800 ;
        RECT 60.400 137.000 61.200 139.800 ;
        RECT 62.000 137.000 62.800 139.800 ;
        RECT 63.600 137.000 64.400 139.800 ;
        RECT 65.200 137.000 66.000 139.800 ;
        RECT 68.400 137.000 69.200 139.800 ;
        RECT 71.600 137.000 72.400 139.800 ;
        RECT 73.200 137.000 74.000 139.800 ;
        RECT 74.800 137.000 75.600 139.800 ;
        RECT 57.200 135.800 59.600 136.600 ;
        RECT 76.400 136.600 77.200 139.800 ;
        RECT 57.200 135.200 58.000 135.800 ;
        RECT 52.000 134.000 53.200 134.600 ;
        RECT 56.200 134.600 58.000 135.200 ;
        RECT 62.000 135.600 63.000 136.400 ;
        RECT 66.000 135.600 67.600 136.400 ;
        RECT 68.400 135.800 73.000 136.400 ;
        RECT 76.400 135.800 79.000 136.600 ;
        RECT 68.400 135.600 69.200 135.800 ;
        RECT 52.000 132.000 52.600 134.000 ;
        RECT 56.200 133.400 57.000 134.600 ;
        RECT 53.200 132.600 57.000 133.400 ;
        RECT 62.000 132.800 62.800 135.600 ;
        RECT 68.400 134.800 69.200 135.000 ;
        RECT 64.800 134.200 69.200 134.800 ;
        RECT 64.800 134.000 65.600 134.200 ;
        RECT 70.000 133.600 70.800 135.200 ;
        RECT 72.200 133.400 73.000 135.800 ;
        RECT 78.200 135.200 79.000 135.800 ;
        RECT 78.200 134.400 81.200 135.200 ;
        RECT 82.800 133.800 83.600 139.800 ;
        RECT 86.000 137.800 86.800 139.800 ;
        RECT 84.400 135.600 85.200 137.200 ;
        RECT 86.200 134.400 86.800 137.800 ;
        RECT 65.200 132.600 68.400 133.400 ;
        RECT 72.200 132.600 74.200 133.400 ;
        RECT 74.800 133.000 83.600 133.800 ;
        RECT 86.000 133.600 86.800 134.400 ;
        RECT 58.800 132.000 59.600 132.600 ;
        RECT 70.000 132.000 70.800 132.400 ;
        RECT 76.400 132.000 77.200 132.400 ;
        RECT 79.600 132.000 80.400 132.400 ;
        RECT 81.400 132.000 82.200 132.200 ;
        RECT 52.000 131.400 52.800 132.000 ;
        RECT 58.800 131.400 82.200 132.000 ;
        RECT 50.600 130.000 51.600 130.800 ;
        RECT 19.800 122.200 20.600 129.600 ;
        RECT 21.400 128.400 22.000 129.600 ;
        RECT 21.200 127.600 22.000 128.400 ;
        RECT 23.800 127.000 24.400 129.600 ;
        RECT 25.200 127.600 26.000 129.200 ;
        RECT 30.200 127.000 30.800 129.600 ;
        RECT 31.600 127.600 32.400 129.200 ;
        RECT 23.800 126.400 27.400 127.000 ;
        RECT 23.800 126.200 24.400 126.400 ;
        RECT 23.600 122.200 24.400 126.200 ;
        RECT 26.800 126.200 27.400 126.400 ;
        RECT 30.200 126.400 33.800 127.000 ;
        RECT 30.200 126.200 30.800 126.400 ;
        RECT 26.800 122.200 27.600 126.200 ;
        RECT 30.000 122.200 30.800 126.200 ;
        RECT 33.200 122.200 34.000 126.400 ;
        RECT 39.000 122.200 39.800 129.600 ;
        RECT 40.600 128.400 41.200 129.600 ;
        RECT 40.400 127.600 41.200 128.400 ;
        RECT 43.000 127.000 43.600 129.600 ;
        RECT 44.400 128.300 45.200 129.200 ;
        RECT 49.200 128.300 50.000 128.400 ;
        RECT 44.400 127.700 50.000 128.300 ;
        RECT 44.400 127.600 45.200 127.700 ;
        RECT 49.200 127.600 50.000 127.700 ;
        RECT 43.000 126.400 46.600 127.000 ;
        RECT 43.000 126.200 43.600 126.400 ;
        RECT 42.800 122.200 43.600 126.200 ;
        RECT 46.000 126.200 46.600 126.400 ;
        RECT 46.000 122.200 46.800 126.200 ;
        RECT 50.800 122.200 51.600 130.000 ;
        RECT 52.200 129.600 52.800 131.400 ;
        RECT 52.200 129.000 61.200 129.600 ;
        RECT 52.200 127.400 52.800 129.000 ;
        RECT 60.400 128.800 61.200 129.000 ;
        RECT 63.600 129.000 72.200 129.600 ;
        RECT 63.600 128.800 64.400 129.000 ;
        RECT 55.400 127.600 58.000 128.400 ;
        RECT 52.200 126.800 54.800 127.400 ;
        RECT 54.000 122.200 54.800 126.800 ;
        RECT 57.200 122.200 58.000 127.600 ;
        RECT 58.600 126.800 62.800 127.600 ;
        RECT 60.400 122.200 61.200 125.000 ;
        RECT 62.000 122.200 62.800 125.000 ;
        RECT 63.600 122.200 64.400 125.000 ;
        RECT 65.200 122.200 66.000 128.400 ;
        RECT 68.400 127.600 71.000 128.400 ;
        RECT 71.600 128.200 72.200 129.000 ;
        RECT 73.200 129.400 74.000 129.600 ;
        RECT 73.200 129.000 78.600 129.400 ;
        RECT 73.200 128.800 79.400 129.000 ;
        RECT 78.000 128.200 79.400 128.800 ;
        RECT 71.600 127.600 77.400 128.200 ;
        RECT 80.400 128.000 82.000 128.800 ;
        RECT 80.400 127.600 81.000 128.000 ;
        RECT 68.400 122.200 69.200 127.000 ;
        RECT 71.600 122.200 72.400 127.000 ;
        RECT 76.800 126.800 81.000 127.600 ;
        RECT 82.800 127.400 83.600 133.000 ;
        RECT 86.200 130.400 86.800 133.600 ;
        RECT 87.600 132.300 88.400 132.400 ;
        RECT 89.200 132.300 90.000 139.800 ;
        RECT 95.600 135.800 96.400 139.800 ;
        RECT 97.000 136.400 97.800 137.200 ;
        RECT 90.800 133.600 91.600 135.200 ;
        RECT 94.000 132.800 94.800 134.400 ;
        RECT 87.600 131.700 90.000 132.300 ;
        RECT 87.600 130.800 88.400 131.700 ;
        RECT 86.000 130.200 86.800 130.400 ;
        RECT 86.000 129.400 87.800 130.200 ;
        RECT 81.600 126.800 83.600 127.400 ;
        RECT 73.200 122.200 74.000 125.000 ;
        RECT 74.800 122.200 75.600 125.000 ;
        RECT 78.000 122.200 78.800 126.800 ;
        RECT 81.600 126.200 82.200 126.800 ;
        RECT 81.200 125.600 82.200 126.200 ;
        RECT 81.200 122.200 82.000 125.600 ;
        RECT 87.000 122.200 87.800 129.400 ;
        RECT 89.200 122.200 90.000 131.700 ;
        RECT 92.400 132.200 93.200 132.400 ;
        RECT 95.600 132.200 96.200 135.800 ;
        RECT 97.200 135.600 98.000 136.400 ;
        RECT 98.800 133.800 99.600 139.800 ;
        RECT 105.200 136.600 106.000 139.800 ;
        RECT 106.800 137.000 107.600 139.800 ;
        RECT 108.400 137.000 109.200 139.800 ;
        RECT 110.000 137.000 110.800 139.800 ;
        RECT 113.200 137.000 114.000 139.800 ;
        RECT 116.400 137.000 117.200 139.800 ;
        RECT 118.000 137.000 118.800 139.800 ;
        RECT 119.600 137.000 120.400 139.800 ;
        RECT 121.200 137.000 122.000 139.800 ;
        RECT 103.400 135.800 106.000 136.600 ;
        RECT 122.800 136.600 123.600 139.800 ;
        RECT 109.400 135.800 114.000 136.400 ;
        RECT 103.400 135.200 104.200 135.800 ;
        RECT 101.200 134.400 104.200 135.200 ;
        RECT 98.800 133.000 107.600 133.800 ;
        RECT 109.400 133.400 110.200 135.800 ;
        RECT 113.200 135.600 114.000 135.800 ;
        RECT 114.800 135.600 116.400 136.400 ;
        RECT 119.400 135.600 120.400 136.400 ;
        RECT 122.800 135.800 125.200 136.600 ;
        RECT 111.600 133.600 112.400 135.200 ;
        RECT 113.200 134.800 114.000 135.000 ;
        RECT 113.200 134.200 117.600 134.800 ;
        RECT 116.800 134.000 117.600 134.200 ;
        RECT 97.200 132.200 98.000 132.400 ;
        RECT 92.400 131.600 94.000 132.200 ;
        RECT 95.600 131.600 98.000 132.200 ;
        RECT 93.200 131.200 94.000 131.600 ;
        RECT 97.200 130.200 97.800 131.600 ;
        RECT 92.400 129.600 96.400 130.200 ;
        RECT 92.400 122.200 93.200 129.600 ;
        RECT 95.600 122.200 96.400 129.600 ;
        RECT 97.200 122.200 98.000 130.200 ;
        RECT 98.800 127.400 99.600 133.000 ;
        RECT 108.200 132.600 110.200 133.400 ;
        RECT 114.000 132.600 117.200 133.400 ;
        RECT 119.600 132.800 120.400 135.600 ;
        RECT 124.400 135.200 125.200 135.800 ;
        RECT 124.400 134.600 126.200 135.200 ;
        RECT 125.400 133.400 126.200 134.600 ;
        RECT 129.200 134.600 130.000 139.800 ;
        RECT 130.800 136.000 131.600 139.800 ;
        RECT 130.800 135.200 131.800 136.000 ;
        RECT 129.200 134.000 130.400 134.600 ;
        RECT 125.400 132.600 129.200 133.400 ;
        RECT 100.400 132.200 101.200 132.400 ;
        RECT 100.200 132.000 101.200 132.200 ;
        RECT 105.200 132.000 106.000 132.400 ;
        RECT 122.800 132.000 123.600 132.600 ;
        RECT 129.800 132.000 130.400 134.000 ;
        RECT 100.200 131.400 123.600 132.000 ;
        RECT 129.600 131.400 130.400 132.000 ;
        RECT 129.600 129.600 130.200 131.400 ;
        RECT 131.000 130.800 131.800 135.200 ;
        RECT 108.400 129.400 109.200 129.600 ;
        RECT 103.800 129.000 109.200 129.400 ;
        RECT 103.000 128.800 109.200 129.000 ;
        RECT 110.200 129.000 118.800 129.600 ;
        RECT 100.400 128.000 102.000 128.800 ;
        RECT 103.000 128.200 104.400 128.800 ;
        RECT 110.200 128.200 110.800 129.000 ;
        RECT 118.000 128.800 118.800 129.000 ;
        RECT 121.200 129.000 130.200 129.600 ;
        RECT 121.200 128.800 122.000 129.000 ;
        RECT 101.400 127.600 102.000 128.000 ;
        RECT 105.000 127.600 110.800 128.200 ;
        RECT 111.400 127.600 114.000 128.400 ;
        RECT 98.800 126.800 100.800 127.400 ;
        RECT 101.400 126.800 105.600 127.600 ;
        RECT 100.200 126.200 100.800 126.800 ;
        RECT 100.200 125.600 101.200 126.200 ;
        RECT 100.400 122.200 101.200 125.600 ;
        RECT 103.600 122.200 104.400 126.800 ;
        RECT 106.800 122.200 107.600 125.000 ;
        RECT 108.400 122.200 109.200 125.000 ;
        RECT 110.000 122.200 110.800 127.000 ;
        RECT 113.200 122.200 114.000 127.000 ;
        RECT 116.400 122.200 117.200 128.400 ;
        RECT 124.400 127.600 127.000 128.400 ;
        RECT 119.600 126.800 123.800 127.600 ;
        RECT 118.000 122.200 118.800 125.000 ;
        RECT 119.600 122.200 120.400 125.000 ;
        RECT 121.200 122.200 122.000 125.000 ;
        RECT 124.400 122.200 125.200 127.600 ;
        RECT 129.600 127.400 130.200 129.000 ;
        RECT 127.600 126.800 130.200 127.400 ;
        RECT 130.800 130.000 131.800 130.800 ;
        RECT 127.600 122.200 128.400 126.800 ;
        RECT 130.800 122.200 131.600 130.000 ;
        RECT 137.200 124.300 138.000 124.400 ;
        RECT 140.400 124.300 141.200 139.800 ;
        RECT 142.000 135.600 142.800 137.200 ;
        RECT 143.600 136.000 144.400 139.800 ;
        RECT 146.800 136.000 147.600 139.800 ;
        RECT 143.600 135.800 147.600 136.000 ;
        RECT 148.400 135.800 149.200 139.800 ;
        RECT 150.000 135.800 150.800 139.800 ;
        RECT 154.200 138.400 155.000 139.800 ;
        RECT 154.200 137.600 155.600 138.400 ;
        RECT 154.200 136.800 155.000 137.600 ;
        RECT 157.000 136.800 157.800 139.800 ;
        RECT 154.200 135.800 155.600 136.800 ;
        RECT 143.800 135.400 147.400 135.800 ;
        RECT 144.400 134.400 145.200 134.800 ;
        RECT 148.400 134.400 149.000 135.800 ;
        RECT 150.200 135.600 150.800 135.800 ;
        RECT 150.200 135.200 152.000 135.600 ;
        RECT 150.200 135.000 154.400 135.200 ;
        RECT 151.400 134.600 154.400 135.000 ;
        RECT 153.600 134.400 154.400 134.600 ;
        RECT 143.600 133.800 145.200 134.400 ;
        RECT 146.600 134.300 149.200 134.400 ;
        RECT 150.000 134.300 150.800 134.400 ;
        RECT 143.600 133.600 144.400 133.800 ;
        RECT 146.600 133.700 150.800 134.300 ;
        RECT 152.000 133.800 152.800 134.000 ;
        RECT 146.600 133.600 149.200 133.700 ;
        RECT 145.200 131.600 146.000 133.200 ;
        RECT 146.600 130.200 147.200 133.600 ;
        RECT 150.000 132.800 150.800 133.700 ;
        RECT 151.800 133.200 152.800 133.800 ;
        RECT 151.800 132.400 152.400 133.200 ;
        RECT 151.600 131.600 152.400 132.400 ;
        RECT 153.600 131.000 154.200 134.400 ;
        RECT 155.000 132.400 155.600 135.800 ;
        RECT 154.800 131.600 155.600 132.400 ;
        RECT 151.800 130.400 154.200 131.000 ;
        RECT 148.400 130.300 149.200 130.400 ;
        RECT 150.000 130.300 150.800 130.400 ;
        RECT 148.400 130.200 150.800 130.300 ;
        RECT 137.200 123.700 141.200 124.300 ;
        RECT 137.200 123.600 138.000 123.700 ;
        RECT 140.400 122.200 141.200 123.700 ;
        RECT 146.200 129.600 147.200 130.200 ;
        RECT 147.800 129.700 150.800 130.200 ;
        RECT 147.800 129.600 149.200 129.700 ;
        RECT 150.000 129.600 150.800 129.700 ;
        RECT 146.200 122.200 147.000 129.600 ;
        RECT 147.800 128.400 148.400 129.600 ;
        RECT 147.600 127.600 148.400 128.400 ;
        RECT 151.800 126.200 152.400 130.400 ;
        RECT 155.000 130.200 155.600 131.600 ;
        RECT 151.600 122.200 152.400 126.200 ;
        RECT 154.800 122.200 155.600 130.200 ;
        RECT 156.400 135.800 157.800 136.800 ;
        RECT 161.200 135.800 162.000 139.800 ;
        RECT 164.400 137.800 165.200 139.800 ;
        RECT 156.400 132.400 157.000 135.800 ;
        RECT 161.200 135.600 161.800 135.800 ;
        RECT 160.000 135.200 161.800 135.600 ;
        RECT 157.600 135.000 161.800 135.200 ;
        RECT 157.600 134.600 160.600 135.000 ;
        RECT 157.600 134.400 158.400 134.600 ;
        RECT 164.400 134.400 165.000 137.800 ;
        RECT 166.000 135.600 166.800 137.200 ;
        RECT 167.600 136.000 168.400 139.800 ;
        RECT 170.800 136.000 171.600 139.800 ;
        RECT 167.600 135.800 171.600 136.000 ;
        RECT 172.400 135.800 173.200 139.800 ;
        RECT 174.600 138.400 175.400 139.800 ;
        RECT 174.600 137.600 176.400 138.400 ;
        RECT 174.600 136.400 175.400 137.600 ;
        RECT 174.600 135.800 176.400 136.400 ;
        RECT 167.800 135.400 171.400 135.800 ;
        RECT 168.400 134.400 169.200 134.800 ;
        RECT 172.400 134.400 173.000 135.800 ;
        RECT 156.400 131.600 157.200 132.400 ;
        RECT 156.400 130.400 157.000 131.600 ;
        RECT 157.800 131.000 158.400 134.400 ;
        RECT 159.200 133.800 160.000 134.000 ;
        RECT 159.200 133.200 160.200 133.800 ;
        RECT 159.600 132.400 160.200 133.200 ;
        RECT 161.200 132.800 162.000 134.400 ;
        RECT 164.400 134.300 165.200 134.400 ;
        RECT 167.600 134.300 169.200 134.400 ;
        RECT 164.400 133.800 169.200 134.300 ;
        RECT 164.400 133.700 168.400 133.800 ;
        RECT 164.400 133.600 165.200 133.700 ;
        RECT 167.600 133.600 168.400 133.700 ;
        RECT 170.600 133.600 173.200 134.400 ;
        RECT 159.600 131.600 160.400 132.400 ;
        RECT 157.800 130.400 160.200 131.000 ;
        RECT 162.800 130.800 163.600 132.400 ;
        RECT 156.400 122.200 157.200 130.400 ;
        RECT 159.600 126.200 160.200 130.400 ;
        RECT 164.400 130.200 165.000 133.600 ;
        RECT 169.200 131.600 170.000 133.200 ;
        RECT 170.600 130.200 171.200 133.600 ;
        RECT 172.400 132.300 173.200 132.400 ;
        RECT 172.400 131.700 174.700 132.300 ;
        RECT 172.400 131.600 173.200 131.700 ;
        RECT 174.100 130.400 174.700 131.700 ;
        RECT 172.400 130.200 173.200 130.400 ;
        RECT 163.400 129.400 165.200 130.200 ;
        RECT 170.200 129.600 171.200 130.200 ;
        RECT 171.800 129.600 173.200 130.200 ;
        RECT 159.600 122.200 160.400 126.200 ;
        RECT 163.400 122.200 164.200 129.400 ;
        RECT 170.200 122.200 171.000 129.600 ;
        RECT 171.800 128.400 172.400 129.600 ;
        RECT 174.000 128.800 174.800 130.400 ;
        RECT 171.600 127.600 172.400 128.400 ;
        RECT 175.600 122.200 176.400 135.800 ;
        RECT 177.200 134.300 178.000 135.200 ;
        RECT 178.800 134.300 179.600 139.800 ;
        RECT 180.400 136.300 181.200 137.200 ;
        RECT 182.000 136.300 182.800 136.400 ;
        RECT 180.400 135.700 182.800 136.300 ;
        RECT 183.600 136.000 184.400 139.800 ;
        RECT 180.400 135.600 181.200 135.700 ;
        RECT 182.000 135.600 182.800 135.700 ;
        RECT 177.200 133.700 179.600 134.300 ;
        RECT 177.200 133.600 178.000 133.700 ;
        RECT 178.800 122.200 179.600 133.700 ;
        RECT 183.400 135.200 184.400 136.000 ;
        RECT 183.400 130.800 184.200 135.200 ;
        RECT 185.200 134.600 186.000 139.800 ;
        RECT 191.600 136.600 192.400 139.800 ;
        RECT 193.200 137.000 194.000 139.800 ;
        RECT 194.800 137.000 195.600 139.800 ;
        RECT 196.400 137.000 197.200 139.800 ;
        RECT 198.000 137.000 198.800 139.800 ;
        RECT 201.200 137.000 202.000 139.800 ;
        RECT 204.400 137.000 205.200 139.800 ;
        RECT 206.000 137.000 206.800 139.800 ;
        RECT 207.600 137.000 208.400 139.800 ;
        RECT 190.000 135.800 192.400 136.600 ;
        RECT 209.200 136.600 210.000 139.800 ;
        RECT 190.000 135.200 190.800 135.800 ;
        RECT 184.800 134.000 186.000 134.600 ;
        RECT 189.000 134.600 190.800 135.200 ;
        RECT 194.800 135.600 195.800 136.400 ;
        RECT 198.800 135.600 200.400 136.400 ;
        RECT 201.200 135.800 205.800 136.400 ;
        RECT 209.200 135.800 211.800 136.600 ;
        RECT 201.200 135.600 202.000 135.800 ;
        RECT 184.800 132.000 185.400 134.000 ;
        RECT 189.000 133.400 189.800 134.600 ;
        RECT 186.000 132.600 189.800 133.400 ;
        RECT 194.800 132.800 195.600 135.600 ;
        RECT 201.200 134.800 202.000 135.000 ;
        RECT 197.600 134.200 202.000 134.800 ;
        RECT 197.600 134.000 198.400 134.200 ;
        RECT 202.800 133.600 203.600 135.200 ;
        RECT 205.000 133.400 205.800 135.800 ;
        RECT 211.000 135.200 211.800 135.800 ;
        RECT 211.000 134.400 214.000 135.200 ;
        RECT 215.600 133.800 216.400 139.800 ;
        RECT 218.800 137.800 219.600 139.800 ;
        RECT 217.200 135.600 218.000 137.200 ;
        RECT 219.000 134.400 219.600 137.800 ;
        RECT 222.000 135.800 222.800 139.800 ;
        RECT 223.600 136.000 224.400 139.800 ;
        RECT 226.800 136.000 227.600 139.800 ;
        RECT 223.600 135.800 227.600 136.000 ;
        RECT 228.400 136.000 229.200 139.800 ;
        RECT 231.600 136.000 232.400 139.800 ;
        RECT 228.400 135.800 232.400 136.000 ;
        RECT 233.200 135.800 234.000 139.800 ;
        RECT 222.200 134.400 222.800 135.800 ;
        RECT 223.800 135.400 227.400 135.800 ;
        RECT 228.600 135.400 232.200 135.800 ;
        RECT 226.000 134.400 226.800 134.800 ;
        RECT 229.200 134.400 230.000 134.800 ;
        RECT 233.200 134.400 233.800 135.800 ;
        RECT 198.000 132.600 201.200 133.400 ;
        RECT 205.000 132.600 207.000 133.400 ;
        RECT 207.600 133.000 216.400 133.800 ;
        RECT 218.800 133.600 219.600 134.400 ;
        RECT 222.000 133.600 224.600 134.400 ;
        RECT 226.000 133.800 227.600 134.400 ;
        RECT 226.800 133.600 227.600 133.800 ;
        RECT 228.400 133.800 230.000 134.400 ;
        RECT 228.400 133.600 229.200 133.800 ;
        RECT 231.400 133.600 234.000 134.400 ;
        RECT 236.000 134.200 236.800 139.800 ;
        RECT 235.000 133.800 236.800 134.200 ;
        RECT 235.000 133.600 236.600 133.800 ;
        RECT 191.600 132.000 192.400 132.600 ;
        RECT 209.200 132.000 210.000 132.400 ;
        RECT 210.800 132.000 211.600 132.400 ;
        RECT 214.200 132.000 215.000 132.200 ;
        RECT 184.800 131.400 185.600 132.000 ;
        RECT 191.600 131.400 215.000 132.000 ;
        RECT 183.400 130.000 184.400 130.800 ;
        RECT 183.600 122.200 184.400 130.000 ;
        RECT 185.000 129.600 185.600 131.400 ;
        RECT 185.000 129.000 194.000 129.600 ;
        RECT 185.000 127.400 185.600 129.000 ;
        RECT 193.200 128.800 194.000 129.000 ;
        RECT 196.400 129.000 205.000 129.600 ;
        RECT 196.400 128.800 197.200 129.000 ;
        RECT 188.200 127.600 190.800 128.400 ;
        RECT 185.000 126.800 187.600 127.400 ;
        RECT 186.800 122.200 187.600 126.800 ;
        RECT 190.000 122.200 190.800 127.600 ;
        RECT 191.400 126.800 195.600 127.600 ;
        RECT 193.200 122.200 194.000 125.000 ;
        RECT 194.800 122.200 195.600 125.000 ;
        RECT 196.400 122.200 197.200 125.000 ;
        RECT 198.000 122.200 198.800 128.400 ;
        RECT 201.200 127.600 203.800 128.400 ;
        RECT 204.400 128.200 205.000 129.000 ;
        RECT 206.000 129.400 206.800 129.600 ;
        RECT 206.000 129.000 211.400 129.400 ;
        RECT 206.000 128.800 212.200 129.000 ;
        RECT 210.800 128.200 212.200 128.800 ;
        RECT 204.400 127.600 210.200 128.200 ;
        RECT 213.200 128.000 214.800 128.800 ;
        RECT 213.200 127.600 213.800 128.000 ;
        RECT 201.200 122.200 202.000 127.000 ;
        RECT 204.400 122.200 205.200 127.000 ;
        RECT 209.600 126.800 213.800 127.600 ;
        RECT 215.600 127.400 216.400 133.000 ;
        RECT 219.000 130.200 219.600 133.600 ;
        RECT 220.400 132.300 221.200 132.400 ;
        RECT 224.000 132.300 224.600 133.600 ;
        RECT 220.400 131.700 224.600 132.300 ;
        RECT 220.400 130.800 221.200 131.700 ;
        RECT 222.000 130.200 222.800 130.400 ;
        RECT 224.000 130.200 224.600 131.700 ;
        RECT 225.200 132.300 226.000 133.200 ;
        RECT 226.800 132.300 227.600 132.400 ;
        RECT 230.000 132.300 230.800 133.200 ;
        RECT 225.200 131.700 230.800 132.300 ;
        RECT 225.200 131.600 226.000 131.700 ;
        RECT 226.800 131.600 227.600 131.700 ;
        RECT 230.000 131.600 230.800 131.700 ;
        RECT 231.400 132.400 232.000 133.600 ;
        RECT 231.400 131.600 232.400 132.400 ;
        RECT 233.200 132.300 234.000 132.400 ;
        RECT 235.000 132.300 235.600 133.600 ;
        RECT 233.200 131.700 235.600 132.300 ;
        RECT 233.200 131.600 234.000 131.700 ;
        RECT 231.400 130.200 232.000 131.600 ;
        RECT 235.000 130.400 235.600 131.700 ;
        RECT 237.200 131.600 238.800 132.400 ;
        RECT 233.200 130.200 234.000 130.400 ;
        RECT 218.800 129.400 220.600 130.200 ;
        RECT 222.000 129.600 223.400 130.200 ;
        RECT 224.000 129.600 225.000 130.200 ;
        RECT 214.400 126.800 216.400 127.400 ;
        RECT 206.000 122.200 206.800 125.000 ;
        RECT 207.600 122.200 208.400 125.000 ;
        RECT 210.800 122.200 211.600 126.800 ;
        RECT 214.400 126.200 215.000 126.800 ;
        RECT 214.000 125.600 215.000 126.200 ;
        RECT 214.000 122.200 214.800 125.600 ;
        RECT 219.800 122.200 220.600 129.400 ;
        RECT 222.800 128.400 223.400 129.600 ;
        RECT 222.800 127.600 223.600 128.400 ;
        RECT 224.200 122.200 225.000 129.600 ;
        RECT 231.000 129.600 232.000 130.200 ;
        RECT 232.600 129.600 234.000 130.200 ;
        RECT 234.800 129.600 235.600 130.400 ;
        RECT 239.600 130.300 240.400 131.200 ;
        RECT 241.200 130.300 242.000 139.800 ;
        RECT 242.800 135.600 243.600 137.200 ;
        RECT 245.000 136.400 245.800 139.800 ;
        RECT 250.800 137.600 251.600 139.800 ;
        RECT 255.600 137.800 256.400 139.800 ;
        RECT 245.000 135.800 246.800 136.400 ;
        RECT 244.400 130.300 245.200 130.400 ;
        RECT 239.600 129.700 245.200 130.300 ;
        RECT 239.600 129.600 240.400 129.700 ;
        RECT 231.000 122.200 231.800 129.600 ;
        RECT 232.600 128.400 233.200 129.600 ;
        RECT 232.400 127.600 233.200 128.400 ;
        RECT 235.000 127.000 235.600 129.600 ;
        RECT 236.400 127.600 237.200 129.200 ;
        RECT 235.000 126.400 238.600 127.000 ;
        RECT 235.000 126.200 235.600 126.400 ;
        RECT 234.800 122.200 235.600 126.200 ;
        RECT 238.000 126.200 238.600 126.400 ;
        RECT 238.000 122.200 238.800 126.200 ;
        RECT 241.200 122.200 242.000 129.700 ;
        RECT 244.400 128.800 245.200 129.700 ;
        RECT 246.000 122.200 246.800 135.800 ;
        RECT 247.600 134.300 248.400 135.200 ;
        RECT 250.800 134.400 251.400 137.600 ;
        RECT 252.400 135.600 253.200 137.200 ;
        RECT 254.000 135.600 254.800 137.200 ;
        RECT 255.800 134.400 256.400 137.800 ;
        RECT 258.800 136.000 259.600 139.800 ;
        RECT 262.000 136.000 262.800 139.800 ;
        RECT 258.800 135.800 262.800 136.000 ;
        RECT 263.600 138.300 264.400 139.800 ;
        RECT 265.200 138.300 266.000 138.400 ;
        RECT 263.600 137.700 266.000 138.300 ;
        RECT 263.600 135.800 264.400 137.700 ;
        RECT 265.200 137.600 266.000 137.700 ;
        RECT 273.200 136.000 274.000 139.800 ;
        RECT 259.000 135.400 262.600 135.800 ;
        RECT 259.600 134.400 260.400 134.800 ;
        RECT 263.600 134.400 264.200 135.800 ;
        RECT 273.000 135.200 274.000 136.000 ;
        RECT 249.200 134.300 250.000 134.400 ;
        RECT 247.600 133.700 250.000 134.300 ;
        RECT 247.600 133.600 248.400 133.700 ;
        RECT 249.200 133.600 250.000 133.700 ;
        RECT 250.800 133.600 251.600 134.400 ;
        RECT 252.400 134.300 253.200 134.400 ;
        RECT 255.600 134.300 256.400 134.400 ;
        RECT 252.400 133.700 256.400 134.300 ;
        RECT 252.400 133.600 253.200 133.700 ;
        RECT 255.600 133.600 256.400 133.700 ;
        RECT 258.800 133.800 260.400 134.400 ;
        RECT 258.800 133.600 259.600 133.800 ;
        RECT 261.800 133.600 264.400 134.400 ;
        RECT 249.200 130.800 250.000 132.400 ;
        RECT 250.800 130.200 251.400 133.600 ;
        RECT 255.800 130.200 256.400 133.600 ;
        RECT 257.200 132.300 258.000 132.400 ;
        RECT 258.900 132.300 259.500 133.600 ;
        RECT 257.200 131.700 259.500 132.300 ;
        RECT 257.200 130.800 258.000 131.700 ;
        RECT 260.400 131.600 261.200 133.200 ;
        RECT 261.800 130.200 262.400 133.600 ;
        RECT 273.000 130.800 273.800 135.200 ;
        RECT 274.800 134.600 275.600 139.800 ;
        RECT 281.200 136.600 282.000 139.800 ;
        RECT 282.800 137.000 283.600 139.800 ;
        RECT 284.400 137.000 285.200 139.800 ;
        RECT 286.000 137.000 286.800 139.800 ;
        RECT 287.600 137.000 288.400 139.800 ;
        RECT 290.800 137.000 291.600 139.800 ;
        RECT 294.000 137.000 294.800 139.800 ;
        RECT 295.600 137.000 296.400 139.800 ;
        RECT 297.200 137.000 298.000 139.800 ;
        RECT 279.600 135.800 282.000 136.600 ;
        RECT 298.800 136.600 299.600 139.800 ;
        RECT 279.600 135.200 280.400 135.800 ;
        RECT 274.400 134.000 275.600 134.600 ;
        RECT 278.600 134.600 280.400 135.200 ;
        RECT 284.400 135.600 285.400 136.400 ;
        RECT 288.400 135.600 290.000 136.400 ;
        RECT 290.800 135.800 295.400 136.400 ;
        RECT 298.800 135.800 301.400 136.600 ;
        RECT 290.800 135.600 291.600 135.800 ;
        RECT 274.400 132.000 275.000 134.000 ;
        RECT 278.600 133.400 279.400 134.600 ;
        RECT 275.600 132.600 279.400 133.400 ;
        RECT 284.400 132.800 285.200 135.600 ;
        RECT 290.800 134.800 291.600 135.000 ;
        RECT 287.200 134.200 291.600 134.800 ;
        RECT 287.200 134.000 288.000 134.200 ;
        RECT 292.400 133.600 293.200 135.200 ;
        RECT 294.600 133.400 295.400 135.800 ;
        RECT 300.600 135.200 301.400 135.800 ;
        RECT 300.600 134.400 303.600 135.200 ;
        RECT 305.200 133.800 306.000 139.800 ;
        RECT 306.800 135.800 307.600 139.800 ;
        RECT 308.400 136.000 309.200 139.800 ;
        RECT 311.600 136.000 312.400 139.800 ;
        RECT 308.400 135.800 312.400 136.000 ;
        RECT 307.000 134.400 307.600 135.800 ;
        RECT 308.600 135.400 312.200 135.800 ;
        RECT 310.800 134.400 311.600 134.800 ;
        RECT 287.600 132.600 290.800 133.400 ;
        RECT 294.600 132.600 296.600 133.400 ;
        RECT 297.200 133.000 306.000 133.800 ;
        RECT 306.800 133.600 309.400 134.400 ;
        RECT 310.800 134.300 312.400 134.400 ;
        RECT 313.200 134.300 314.000 139.800 ;
        RECT 314.800 135.600 315.600 137.200 ;
        RECT 316.400 135.800 317.200 139.800 ;
        RECT 318.000 136.000 318.800 139.800 ;
        RECT 321.200 136.000 322.000 139.800 ;
        RECT 318.000 135.800 322.000 136.000 ;
        RECT 316.600 134.400 317.200 135.800 ;
        RECT 318.200 135.400 321.800 135.800 ;
        RECT 320.400 134.400 321.200 134.800 ;
        RECT 310.800 133.800 314.000 134.300 ;
        RECT 311.600 133.700 314.000 133.800 ;
        RECT 311.600 133.600 312.400 133.700 ;
        RECT 274.400 131.400 275.200 132.000 ;
        RECT 263.600 130.200 264.400 130.400 ;
        RECT 249.800 129.400 251.600 130.200 ;
        RECT 255.600 129.400 257.400 130.200 ;
        RECT 249.800 124.400 250.600 129.400 ;
        RECT 249.800 123.600 251.600 124.400 ;
        RECT 249.800 122.200 250.600 123.600 ;
        RECT 256.600 122.200 257.400 129.400 ;
        RECT 261.400 129.600 262.400 130.200 ;
        RECT 263.000 129.600 264.400 130.200 ;
        RECT 273.000 130.000 274.000 130.800 ;
        RECT 261.400 122.200 262.200 129.600 ;
        RECT 263.000 128.400 263.600 129.600 ;
        RECT 262.800 127.600 263.600 128.400 ;
        RECT 273.200 122.200 274.000 130.000 ;
        RECT 274.600 129.600 275.200 131.400 ;
        RECT 275.800 130.800 276.600 131.000 ;
        RECT 275.800 130.300 302.800 130.800 ;
        RECT 303.600 130.300 304.400 130.400 ;
        RECT 275.800 130.200 304.400 130.300 ;
        RECT 298.600 130.000 299.400 130.200 ;
        RECT 302.000 129.700 304.400 130.200 ;
        RECT 302.000 129.600 302.800 129.700 ;
        RECT 303.600 129.600 304.400 129.700 ;
        RECT 274.600 129.000 283.600 129.600 ;
        RECT 274.600 127.400 275.200 129.000 ;
        RECT 282.800 128.800 283.600 129.000 ;
        RECT 286.000 129.000 294.600 129.600 ;
        RECT 286.000 128.800 286.800 129.000 ;
        RECT 277.800 127.600 280.400 128.400 ;
        RECT 274.600 126.800 277.200 127.400 ;
        RECT 276.400 122.200 277.200 126.800 ;
        RECT 279.600 122.200 280.400 127.600 ;
        RECT 281.000 126.800 285.200 127.600 ;
        RECT 282.800 122.200 283.600 125.000 ;
        RECT 284.400 122.200 285.200 125.000 ;
        RECT 286.000 122.200 286.800 125.000 ;
        RECT 287.600 122.200 288.400 128.400 ;
        RECT 290.800 127.600 293.400 128.400 ;
        RECT 294.000 128.200 294.600 129.000 ;
        RECT 295.600 129.400 296.400 129.600 ;
        RECT 295.600 129.000 301.000 129.400 ;
        RECT 295.600 128.800 301.800 129.000 ;
        RECT 300.400 128.200 301.800 128.800 ;
        RECT 294.000 127.600 299.800 128.200 ;
        RECT 302.800 128.000 304.400 128.800 ;
        RECT 302.800 127.600 303.400 128.000 ;
        RECT 290.800 122.200 291.600 127.000 ;
        RECT 294.000 122.200 294.800 127.000 ;
        RECT 299.200 126.800 303.400 127.600 ;
        RECT 305.200 127.400 306.000 133.000 ;
        RECT 306.800 130.200 307.600 130.400 ;
        RECT 308.800 130.200 309.400 133.600 ;
        RECT 310.000 131.600 310.800 133.200 ;
        RECT 306.800 129.600 308.200 130.200 ;
        RECT 308.800 129.600 309.800 130.200 ;
        RECT 307.600 128.400 308.200 129.600 ;
        RECT 307.600 127.600 308.400 128.400 ;
        RECT 304.000 126.800 306.000 127.400 ;
        RECT 295.600 122.200 296.400 125.000 ;
        RECT 297.200 122.200 298.000 125.000 ;
        RECT 300.400 122.200 301.200 126.800 ;
        RECT 304.000 126.200 304.600 126.800 ;
        RECT 303.600 125.600 304.600 126.200 ;
        RECT 303.600 122.200 304.400 125.600 ;
        RECT 309.000 122.200 309.800 129.600 ;
        RECT 313.200 122.200 314.000 133.700 ;
        RECT 316.400 133.600 319.000 134.400 ;
        RECT 320.400 133.800 322.000 134.400 ;
        RECT 321.200 133.600 322.000 133.800 ;
        RECT 322.800 133.800 323.600 139.800 ;
        RECT 329.200 136.600 330.000 139.800 ;
        RECT 330.800 137.000 331.600 139.800 ;
        RECT 332.400 137.000 333.200 139.800 ;
        RECT 334.000 137.000 334.800 139.800 ;
        RECT 337.200 137.000 338.000 139.800 ;
        RECT 340.400 137.000 341.200 139.800 ;
        RECT 342.000 137.000 342.800 139.800 ;
        RECT 343.600 137.000 344.400 139.800 ;
        RECT 345.200 137.000 346.000 139.800 ;
        RECT 327.400 135.800 330.000 136.600 ;
        RECT 346.800 136.600 347.600 139.800 ;
        RECT 333.400 135.800 338.000 136.400 ;
        RECT 327.400 135.200 328.200 135.800 ;
        RECT 325.200 134.400 328.200 135.200 ;
        RECT 314.800 130.300 315.600 130.400 ;
        RECT 316.400 130.300 317.200 130.400 ;
        RECT 314.800 130.200 317.200 130.300 ;
        RECT 318.400 130.200 319.000 133.600 ;
        RECT 322.800 133.000 331.600 133.800 ;
        RECT 333.400 133.400 334.200 135.800 ;
        RECT 337.200 135.600 338.000 135.800 ;
        RECT 338.800 135.600 340.400 136.400 ;
        RECT 343.400 135.600 344.400 136.400 ;
        RECT 346.800 135.800 349.200 136.600 ;
        RECT 335.600 133.600 336.400 135.200 ;
        RECT 337.200 134.800 338.000 135.000 ;
        RECT 337.200 134.200 341.600 134.800 ;
        RECT 340.800 134.000 341.600 134.200 ;
        RECT 314.800 129.700 317.800 130.200 ;
        RECT 314.800 129.600 315.600 129.700 ;
        RECT 316.400 129.600 317.800 129.700 ;
        RECT 318.400 129.600 319.400 130.200 ;
        RECT 317.200 128.400 317.800 129.600 ;
        RECT 317.200 127.600 318.000 128.400 ;
        RECT 318.600 122.200 319.400 129.600 ;
        RECT 322.800 127.400 323.600 133.000 ;
        RECT 332.200 132.600 334.200 133.400 ;
        RECT 338.000 132.600 341.200 133.400 ;
        RECT 343.600 132.800 344.400 135.600 ;
        RECT 348.400 135.200 349.200 135.800 ;
        RECT 348.400 134.600 350.200 135.200 ;
        RECT 349.400 133.400 350.200 134.600 ;
        RECT 353.200 134.600 354.000 139.800 ;
        RECT 354.800 136.300 355.600 139.800 ;
        RECT 356.400 136.300 357.200 136.400 ;
        RECT 354.800 135.700 357.200 136.300 ;
        RECT 354.800 135.200 355.800 135.700 ;
        RECT 356.400 135.600 357.200 135.700 ;
        RECT 353.200 134.000 354.400 134.600 ;
        RECT 349.400 132.600 353.200 133.400 ;
        RECT 324.200 132.000 325.000 132.200 ;
        RECT 326.000 132.000 326.800 132.400 ;
        RECT 329.200 132.000 330.000 132.400 ;
        RECT 346.800 132.000 347.600 132.600 ;
        RECT 353.800 132.000 354.400 134.000 ;
        RECT 324.200 131.400 347.600 132.000 ;
        RECT 353.600 131.400 354.400 132.000 ;
        RECT 353.600 129.600 354.200 131.400 ;
        RECT 355.000 130.800 355.800 135.200 ;
        RECT 332.400 129.400 333.200 129.600 ;
        RECT 327.800 129.000 333.200 129.400 ;
        RECT 327.000 128.800 333.200 129.000 ;
        RECT 334.200 129.000 342.800 129.600 ;
        RECT 324.400 128.000 326.000 128.800 ;
        RECT 327.000 128.200 328.400 128.800 ;
        RECT 334.200 128.200 334.800 129.000 ;
        RECT 342.000 128.800 342.800 129.000 ;
        RECT 345.200 129.000 354.200 129.600 ;
        RECT 345.200 128.800 346.000 129.000 ;
        RECT 325.400 127.600 326.000 128.000 ;
        RECT 329.000 127.600 334.800 128.200 ;
        RECT 335.400 127.600 338.000 128.400 ;
        RECT 322.800 126.800 324.800 127.400 ;
        RECT 325.400 126.800 329.600 127.600 ;
        RECT 324.200 126.200 324.800 126.800 ;
        RECT 324.200 125.600 325.200 126.200 ;
        RECT 324.400 122.200 325.200 125.600 ;
        RECT 327.600 122.200 328.400 126.800 ;
        RECT 330.800 122.200 331.600 125.000 ;
        RECT 332.400 122.200 333.200 125.000 ;
        RECT 334.000 122.200 334.800 127.000 ;
        RECT 337.200 122.200 338.000 127.000 ;
        RECT 340.400 122.200 341.200 128.400 ;
        RECT 348.400 127.600 351.000 128.400 ;
        RECT 343.600 126.800 347.800 127.600 ;
        RECT 342.000 122.200 342.800 125.000 ;
        RECT 343.600 122.200 344.400 125.000 ;
        RECT 345.200 122.200 346.000 125.000 ;
        RECT 348.400 122.200 349.200 127.600 ;
        RECT 353.600 127.400 354.200 129.000 ;
        RECT 351.600 126.800 354.200 127.400 ;
        RECT 354.800 130.000 355.800 130.800 ;
        RECT 359.600 134.300 360.400 139.800 ;
        RECT 361.200 135.600 362.000 137.200 ;
        RECT 361.200 134.300 362.000 134.400 ;
        RECT 359.600 133.700 362.000 134.300 ;
        RECT 351.600 122.200 352.400 126.800 ;
        RECT 354.800 122.200 355.600 130.000 ;
        RECT 359.600 122.200 360.400 133.700 ;
        RECT 361.200 133.600 362.000 133.700 ;
        RECT 362.800 122.200 363.600 139.800 ;
        RECT 364.400 139.200 368.400 139.800 ;
        RECT 364.400 135.800 365.200 139.200 ;
        RECT 366.000 135.800 366.800 138.600 ;
        RECT 367.600 136.000 368.400 139.200 ;
        RECT 370.800 136.000 371.600 139.800 ;
        RECT 367.600 135.800 371.600 136.000 ;
        RECT 375.600 135.800 376.400 139.800 ;
        RECT 380.400 137.800 381.200 139.800 ;
        RECT 377.000 136.400 377.800 137.200 ;
        RECT 366.000 134.400 366.600 135.800 ;
        RECT 367.800 135.400 371.400 135.800 ;
        RECT 370.000 134.400 370.800 134.800 ;
        RECT 364.400 132.800 365.200 134.400 ;
        RECT 366.000 133.800 368.400 134.400 ;
        RECT 370.000 133.800 371.600 134.400 ;
        RECT 367.600 133.600 368.400 133.800 ;
        RECT 370.800 133.600 371.600 133.800 ;
        RECT 366.000 131.600 366.800 133.200 ;
        RECT 367.800 132.400 368.400 133.600 ;
        RECT 367.600 131.600 368.400 132.400 ;
        RECT 369.200 131.600 370.000 133.200 ;
        RECT 374.000 132.800 374.800 134.400 ;
        RECT 372.400 132.200 373.200 132.400 ;
        RECT 375.600 132.200 376.200 135.800 ;
        RECT 377.200 135.600 378.000 136.400 ;
        RECT 378.800 135.600 379.600 137.200 ;
        RECT 377.300 134.300 377.900 135.600 ;
        RECT 380.600 134.400 381.200 137.800 ;
        RECT 386.600 135.800 388.200 139.800 ;
        RECT 380.400 134.300 381.200 134.400 ;
        RECT 377.300 133.700 381.200 134.300 ;
        RECT 380.400 133.600 381.200 133.700 ;
        RECT 382.000 134.300 382.800 134.400 ;
        RECT 385.200 134.300 386.000 134.400 ;
        RECT 382.000 133.700 386.000 134.300 ;
        RECT 382.000 133.600 382.800 133.700 ;
        RECT 377.200 132.200 378.000 132.400 ;
        RECT 372.400 131.600 374.000 132.200 ;
        RECT 375.600 131.600 378.000 132.200 ;
        RECT 367.800 130.200 368.400 131.600 ;
        RECT 373.200 131.200 374.000 131.600 ;
        RECT 377.200 130.200 377.800 131.600 ;
        RECT 380.600 130.200 381.200 133.600 ;
        RECT 385.200 132.800 386.000 133.700 ;
        RECT 387.000 132.400 387.600 135.800 ;
        RECT 388.400 134.300 389.200 134.400 ;
        RECT 391.600 134.300 392.400 139.800 ;
        RECT 393.200 135.600 394.000 137.200 ;
        RECT 396.400 136.000 397.200 139.800 ;
        RECT 388.400 133.700 392.400 134.300 ;
        RECT 388.400 133.600 389.200 133.700 ;
        RECT 388.400 133.200 389.000 133.600 ;
        RECT 388.200 132.400 389.000 133.200 ;
        RECT 382.000 130.800 382.800 132.400 ;
        RECT 383.600 132.200 384.400 132.400 ;
        RECT 383.600 131.600 385.200 132.200 ;
        RECT 386.800 131.600 387.600 132.400 ;
        RECT 384.400 131.200 385.200 131.600 ;
        RECT 387.000 131.400 387.600 131.600 ;
        RECT 387.000 130.800 389.000 131.400 ;
        RECT 390.000 130.800 390.800 132.400 ;
        RECT 388.400 130.200 389.000 130.800 ;
        RECT 367.000 122.200 369.000 130.200 ;
        RECT 372.400 129.600 376.400 130.200 ;
        RECT 372.400 122.200 373.200 129.600 ;
        RECT 375.600 122.200 376.400 129.600 ;
        RECT 377.200 122.200 378.000 130.200 ;
        RECT 380.400 129.400 382.200 130.200 ;
        RECT 381.400 122.200 382.200 129.400 ;
        RECT 383.600 129.600 387.600 130.200 ;
        RECT 383.600 122.200 384.400 129.600 ;
        RECT 386.800 122.800 387.600 129.600 ;
        RECT 388.400 123.400 389.200 130.200 ;
        RECT 390.000 122.800 390.800 130.200 ;
        RECT 386.800 122.200 390.800 122.800 ;
        RECT 391.600 122.200 392.400 133.700 ;
        RECT 396.200 135.200 397.200 136.000 ;
        RECT 396.200 130.800 397.000 135.200 ;
        RECT 398.000 134.600 398.800 139.800 ;
        RECT 404.400 136.600 405.200 139.800 ;
        RECT 406.000 137.000 406.800 139.800 ;
        RECT 407.600 137.000 408.400 139.800 ;
        RECT 409.200 137.000 410.000 139.800 ;
        RECT 410.800 137.000 411.600 139.800 ;
        RECT 414.000 137.000 414.800 139.800 ;
        RECT 417.200 137.000 418.000 139.800 ;
        RECT 418.800 137.000 419.600 139.800 ;
        RECT 420.400 137.000 421.200 139.800 ;
        RECT 402.800 135.800 405.200 136.600 ;
        RECT 422.000 136.600 422.800 139.800 ;
        RECT 402.800 135.200 403.600 135.800 ;
        RECT 397.600 134.000 398.800 134.600 ;
        RECT 401.800 134.600 403.600 135.200 ;
        RECT 407.600 135.600 408.600 136.400 ;
        RECT 411.600 135.600 413.200 136.400 ;
        RECT 414.000 135.800 418.600 136.400 ;
        RECT 422.000 135.800 424.600 136.600 ;
        RECT 414.000 135.600 414.800 135.800 ;
        RECT 397.600 132.000 398.200 134.000 ;
        RECT 401.800 133.400 402.600 134.600 ;
        RECT 398.800 132.600 402.600 133.400 ;
        RECT 407.600 132.800 408.400 135.600 ;
        RECT 414.000 134.800 414.800 135.000 ;
        RECT 410.400 134.200 414.800 134.800 ;
        RECT 410.400 134.000 411.200 134.200 ;
        RECT 415.600 133.600 416.400 135.200 ;
        RECT 417.800 133.400 418.600 135.800 ;
        RECT 423.800 135.200 424.600 135.800 ;
        RECT 423.800 134.400 426.800 135.200 ;
        RECT 428.400 133.800 429.200 139.800 ;
        RECT 438.000 137.800 438.800 139.800 ;
        RECT 436.400 135.600 437.200 137.200 ;
        RECT 438.200 134.400 438.800 137.800 ;
        RECT 444.400 135.800 445.200 139.800 ;
        RECT 451.200 138.400 452.000 139.800 ;
        RECT 450.800 137.600 452.000 138.400 ;
        RECT 445.800 136.400 446.600 137.200 ;
        RECT 410.800 132.600 414.000 133.400 ;
        RECT 417.800 132.600 419.800 133.400 ;
        RECT 420.400 133.000 429.200 133.800 ;
        RECT 438.000 133.600 438.800 134.400 ;
        RECT 404.400 132.000 405.200 132.600 ;
        RECT 422.000 132.000 422.800 132.400 ;
        RECT 425.200 132.000 426.000 132.400 ;
        RECT 427.000 132.000 427.800 132.200 ;
        RECT 397.600 131.400 398.400 132.000 ;
        RECT 404.400 131.400 427.800 132.000 ;
        RECT 396.200 130.000 397.200 130.800 ;
        RECT 396.400 122.200 397.200 130.000 ;
        RECT 397.800 129.600 398.400 131.400 ;
        RECT 397.800 129.000 406.800 129.600 ;
        RECT 397.800 127.400 398.400 129.000 ;
        RECT 406.000 128.800 406.800 129.000 ;
        RECT 409.200 129.000 417.800 129.600 ;
        RECT 409.200 128.800 410.000 129.000 ;
        RECT 401.000 127.600 403.600 128.400 ;
        RECT 397.800 126.800 400.400 127.400 ;
        RECT 399.600 122.200 400.400 126.800 ;
        RECT 402.800 122.200 403.600 127.600 ;
        RECT 404.200 126.800 408.400 127.600 ;
        RECT 406.000 122.200 406.800 125.000 ;
        RECT 407.600 122.200 408.400 125.000 ;
        RECT 409.200 122.200 410.000 125.000 ;
        RECT 410.800 122.200 411.600 128.400 ;
        RECT 414.000 127.600 416.600 128.400 ;
        RECT 417.200 128.200 417.800 129.000 ;
        RECT 418.800 129.400 419.600 129.600 ;
        RECT 418.800 129.000 424.200 129.400 ;
        RECT 418.800 128.800 425.000 129.000 ;
        RECT 423.600 128.200 425.000 128.800 ;
        RECT 417.200 127.600 423.000 128.200 ;
        RECT 426.000 128.000 427.600 128.800 ;
        RECT 426.000 127.600 426.600 128.000 ;
        RECT 414.000 122.200 414.800 127.000 ;
        RECT 417.200 122.200 418.000 127.000 ;
        RECT 422.400 126.800 426.600 127.600 ;
        RECT 428.400 127.400 429.200 133.000 ;
        RECT 434.800 132.300 435.600 132.400 ;
        RECT 438.200 132.300 438.800 133.600 ;
        RECT 442.800 132.800 443.600 134.400 ;
        RECT 434.800 131.700 438.800 132.300 ;
        RECT 434.800 131.600 435.600 131.700 ;
        RECT 438.200 130.200 438.800 131.700 ;
        RECT 439.600 130.800 440.400 132.400 ;
        RECT 441.200 132.200 442.000 132.400 ;
        RECT 444.400 132.200 445.000 135.800 ;
        RECT 446.000 135.600 446.800 136.400 ;
        RECT 451.200 134.200 452.000 137.600 ;
        RECT 454.000 136.000 454.800 139.800 ;
        RECT 457.200 139.200 461.200 139.800 ;
        RECT 457.200 136.000 458.000 139.200 ;
        RECT 454.000 135.800 458.000 136.000 ;
        RECT 458.800 135.800 459.600 138.600 ;
        RECT 460.400 135.800 461.200 139.200 ;
        RECT 454.200 135.400 457.800 135.800 ;
        RECT 454.800 134.400 455.600 134.800 ;
        RECT 459.000 134.400 459.600 135.800 ;
        RECT 451.200 133.800 453.000 134.200 ;
        RECT 451.400 133.600 453.000 133.800 ;
        RECT 454.000 133.800 455.600 134.400 ;
        RECT 457.200 133.800 459.600 134.400 ;
        RECT 460.400 134.300 461.200 134.400 ;
        RECT 462.000 134.300 462.800 139.800 ;
        RECT 463.600 135.600 464.400 137.200 ;
        RECT 454.000 133.600 454.800 133.800 ;
        RECT 457.200 133.600 458.000 133.800 ;
        RECT 460.400 133.700 462.800 134.300 ;
        RECT 446.000 132.200 446.800 132.400 ;
        RECT 441.200 131.600 442.800 132.200 ;
        RECT 444.400 131.600 446.800 132.200 ;
        RECT 449.200 131.600 450.800 132.400 ;
        RECT 442.000 131.200 442.800 131.600 ;
        RECT 446.000 130.200 446.600 131.600 ;
        RECT 438.000 129.400 439.800 130.200 ;
        RECT 427.200 126.800 429.200 127.400 ;
        RECT 418.800 122.200 419.600 125.000 ;
        RECT 420.400 122.200 421.200 125.000 ;
        RECT 423.600 122.200 424.400 126.800 ;
        RECT 427.200 126.200 427.800 126.800 ;
        RECT 426.800 125.600 427.800 126.200 ;
        RECT 426.800 122.200 427.600 125.600 ;
        RECT 439.000 122.200 439.800 129.400 ;
        RECT 441.200 129.600 445.200 130.200 ;
        RECT 441.200 122.200 442.000 129.600 ;
        RECT 444.400 122.200 445.200 129.600 ;
        RECT 446.000 128.300 446.800 130.200 ;
        RECT 447.600 129.600 448.400 131.200 ;
        RECT 452.400 130.400 453.000 133.600 ;
        RECT 455.600 131.600 456.400 133.200 ;
        RECT 452.400 129.600 453.200 130.400 ;
        RECT 457.200 130.200 457.800 133.600 ;
        RECT 458.800 131.600 459.600 133.200 ;
        RECT 460.400 132.800 461.200 133.700 ;
        RECT 450.800 128.300 451.600 129.200 ;
        RECT 446.000 127.700 451.600 128.300 ;
        RECT 446.000 122.200 446.800 127.700 ;
        RECT 450.800 127.600 451.600 127.700 ;
        RECT 452.400 127.000 453.000 129.600 ;
        RECT 449.400 126.400 453.000 127.000 ;
        RECT 449.400 126.200 450.000 126.400 ;
        RECT 449.200 122.200 450.000 126.200 ;
        RECT 452.400 126.200 453.000 126.400 ;
        RECT 452.400 122.200 453.200 126.200 ;
        RECT 456.600 122.200 458.600 130.200 ;
        RECT 462.000 122.200 462.800 133.700 ;
        RECT 465.200 133.800 466.000 139.800 ;
        RECT 471.600 136.600 472.400 139.800 ;
        RECT 473.200 137.000 474.000 139.800 ;
        RECT 474.800 137.000 475.600 139.800 ;
        RECT 476.400 137.000 477.200 139.800 ;
        RECT 479.600 137.000 480.400 139.800 ;
        RECT 482.800 137.000 483.600 139.800 ;
        RECT 484.400 137.000 485.200 139.800 ;
        RECT 486.000 137.000 486.800 139.800 ;
        RECT 487.600 137.000 488.400 139.800 ;
        RECT 469.800 135.800 472.400 136.600 ;
        RECT 489.200 136.600 490.000 139.800 ;
        RECT 475.800 135.800 480.400 136.400 ;
        RECT 469.800 135.200 470.600 135.800 ;
        RECT 467.600 134.400 470.600 135.200 ;
        RECT 465.200 133.000 474.000 133.800 ;
        RECT 475.800 133.400 476.600 135.800 ;
        RECT 479.600 135.600 480.400 135.800 ;
        RECT 481.200 135.600 482.800 136.400 ;
        RECT 485.800 135.600 486.800 136.400 ;
        RECT 489.200 135.800 491.600 136.600 ;
        RECT 478.000 133.600 478.800 135.200 ;
        RECT 479.600 134.800 480.400 135.000 ;
        RECT 479.600 134.200 484.000 134.800 ;
        RECT 483.200 134.000 484.000 134.200 ;
        RECT 465.200 127.400 466.000 133.000 ;
        RECT 474.600 132.600 476.600 133.400 ;
        RECT 480.400 132.600 483.600 133.400 ;
        RECT 486.000 132.800 486.800 135.600 ;
        RECT 490.800 135.200 491.600 135.800 ;
        RECT 490.800 134.600 492.600 135.200 ;
        RECT 491.800 133.400 492.600 134.600 ;
        RECT 495.600 134.600 496.400 139.800 ;
        RECT 497.200 136.000 498.000 139.800 ;
        RECT 500.400 137.000 501.200 139.000 ;
        RECT 497.200 135.200 498.200 136.000 ;
        RECT 495.600 134.000 496.800 134.600 ;
        RECT 491.800 132.600 495.600 133.400 ;
        RECT 466.600 132.000 467.400 132.200 ;
        RECT 470.000 132.000 470.800 132.400 ;
        RECT 471.600 132.000 472.400 132.400 ;
        RECT 489.200 132.000 490.000 132.600 ;
        RECT 496.200 132.000 496.800 134.000 ;
        RECT 466.600 131.400 490.000 132.000 ;
        RECT 496.000 131.400 496.800 132.000 ;
        RECT 496.000 129.600 496.600 131.400 ;
        RECT 497.400 130.800 498.200 135.200 ;
        RECT 500.400 134.800 501.000 137.000 ;
        RECT 504.600 136.000 505.400 139.000 ;
        RECT 512.600 136.400 513.400 139.800 ;
        RECT 504.600 135.400 506.200 136.000 ;
        RECT 505.400 135.000 506.200 135.400 ;
        RECT 511.600 135.800 513.400 136.400 ;
        RECT 514.800 136.300 515.600 136.400 ;
        RECT 516.400 136.300 517.200 139.800 ;
        RECT 500.400 134.200 504.600 134.800 ;
        RECT 503.600 133.800 504.600 134.200 ;
        RECT 505.600 134.400 506.200 135.000 ;
        RECT 500.400 131.600 501.200 133.200 ;
        RECT 502.000 131.600 502.800 133.200 ;
        RECT 503.600 133.000 505.000 133.800 ;
        RECT 505.600 133.600 507.600 134.400 ;
        RECT 510.000 133.600 510.800 135.200 ;
        RECT 503.600 131.000 504.200 133.000 ;
        RECT 474.800 129.400 475.600 129.600 ;
        RECT 470.200 129.000 475.600 129.400 ;
        RECT 469.400 128.800 475.600 129.000 ;
        RECT 476.600 129.000 485.200 129.600 ;
        RECT 466.800 128.000 468.400 128.800 ;
        RECT 469.400 128.200 470.800 128.800 ;
        RECT 476.600 128.200 477.200 129.000 ;
        RECT 484.400 128.800 485.200 129.000 ;
        RECT 487.600 129.000 496.600 129.600 ;
        RECT 487.600 128.800 488.400 129.000 ;
        RECT 467.800 127.600 468.400 128.000 ;
        RECT 471.400 127.600 477.200 128.200 ;
        RECT 477.800 127.600 480.400 128.400 ;
        RECT 465.200 126.800 467.200 127.400 ;
        RECT 467.800 126.800 472.000 127.600 ;
        RECT 466.600 126.200 467.200 126.800 ;
        RECT 466.600 125.600 467.600 126.200 ;
        RECT 466.800 122.200 467.600 125.600 ;
        RECT 470.000 122.200 470.800 126.800 ;
        RECT 473.200 122.200 474.000 125.000 ;
        RECT 474.800 122.200 475.600 125.000 ;
        RECT 476.400 122.200 477.200 127.000 ;
        RECT 479.600 122.200 480.400 127.000 ;
        RECT 482.800 122.200 483.600 128.400 ;
        RECT 490.800 127.600 493.400 128.400 ;
        RECT 486.000 126.800 490.200 127.600 ;
        RECT 484.400 122.200 485.200 125.000 ;
        RECT 486.000 122.200 486.800 125.000 ;
        RECT 487.600 122.200 488.400 125.000 ;
        RECT 490.800 122.200 491.600 127.600 ;
        RECT 496.000 127.400 496.600 129.000 ;
        RECT 494.000 126.800 496.600 127.400 ;
        RECT 497.200 130.000 498.200 130.800 ;
        RECT 500.400 130.400 504.200 131.000 ;
        RECT 494.000 122.200 494.800 126.800 ;
        RECT 497.200 122.200 498.000 130.000 ;
        RECT 500.400 127.000 501.000 130.400 ;
        RECT 505.600 129.800 506.200 133.600 ;
        RECT 506.800 130.800 507.600 132.400 ;
        RECT 504.600 129.200 506.200 129.800 ;
        RECT 500.400 123.000 501.200 127.000 ;
        RECT 504.600 124.400 505.400 129.200 ;
        RECT 510.000 128.300 510.800 128.400 ;
        RECT 511.600 128.300 512.400 135.800 ;
        RECT 514.800 135.700 517.200 136.300 ;
        RECT 514.800 135.600 515.600 135.700 ;
        RECT 516.200 135.200 517.200 135.700 ;
        RECT 516.200 130.800 517.000 135.200 ;
        RECT 518.000 134.600 518.800 139.800 ;
        RECT 524.400 136.600 525.200 139.800 ;
        RECT 526.000 137.000 526.800 139.800 ;
        RECT 527.600 137.000 528.400 139.800 ;
        RECT 529.200 137.000 530.000 139.800 ;
        RECT 530.800 137.000 531.600 139.800 ;
        RECT 534.000 137.000 534.800 139.800 ;
        RECT 537.200 137.000 538.000 139.800 ;
        RECT 538.800 137.000 539.600 139.800 ;
        RECT 540.400 137.000 541.200 139.800 ;
        RECT 522.800 135.800 525.200 136.600 ;
        RECT 542.000 136.600 542.800 139.800 ;
        RECT 522.800 135.200 523.600 135.800 ;
        RECT 517.600 134.000 518.800 134.600 ;
        RECT 521.800 134.600 523.600 135.200 ;
        RECT 527.600 135.600 528.600 136.400 ;
        RECT 531.600 135.600 533.200 136.400 ;
        RECT 534.000 135.800 538.600 136.400 ;
        RECT 542.000 135.800 544.600 136.600 ;
        RECT 534.000 135.600 534.800 135.800 ;
        RECT 517.600 132.000 518.200 134.000 ;
        RECT 521.800 133.400 522.600 134.600 ;
        RECT 518.800 132.600 522.600 133.400 ;
        RECT 527.600 132.800 528.400 135.600 ;
        RECT 534.000 134.800 534.800 135.000 ;
        RECT 530.400 134.200 534.800 134.800 ;
        RECT 530.400 134.000 531.200 134.200 ;
        RECT 535.600 133.600 536.400 135.200 ;
        RECT 537.800 133.400 538.600 135.800 ;
        RECT 543.800 135.200 544.600 135.800 ;
        RECT 543.800 134.400 546.800 135.200 ;
        RECT 548.400 133.800 549.200 139.800 ;
        RECT 530.800 132.600 534.000 133.400 ;
        RECT 537.800 132.600 539.800 133.400 ;
        RECT 540.400 133.000 549.200 133.800 ;
        RECT 524.400 132.000 525.200 132.600 ;
        RECT 542.000 132.000 542.800 132.400 ;
        RECT 543.600 132.000 544.400 132.400 ;
        RECT 547.000 132.000 547.800 132.200 ;
        RECT 517.600 131.400 518.400 132.000 ;
        RECT 524.400 131.400 547.800 132.000 ;
        RECT 513.200 128.800 514.000 130.400 ;
        RECT 516.200 130.000 517.200 130.800 ;
        RECT 510.000 127.700 512.400 128.300 ;
        RECT 510.000 127.600 510.800 127.700 ;
        RECT 504.600 123.600 506.000 124.400 ;
        RECT 504.600 122.200 505.400 123.600 ;
        RECT 511.600 122.200 512.400 127.700 ;
        RECT 516.400 122.200 517.200 130.000 ;
        RECT 517.800 129.600 518.400 131.400 ;
        RECT 517.800 129.000 526.800 129.600 ;
        RECT 517.800 127.400 518.400 129.000 ;
        RECT 526.000 128.800 526.800 129.000 ;
        RECT 529.200 129.000 537.800 129.600 ;
        RECT 529.200 128.800 530.000 129.000 ;
        RECT 521.000 127.600 523.600 128.400 ;
        RECT 517.800 126.800 520.400 127.400 ;
        RECT 519.600 122.200 520.400 126.800 ;
        RECT 522.800 122.200 523.600 127.600 ;
        RECT 524.200 126.800 528.400 127.600 ;
        RECT 526.000 122.200 526.800 125.000 ;
        RECT 527.600 122.200 528.400 125.000 ;
        RECT 529.200 122.200 530.000 125.000 ;
        RECT 530.800 122.200 531.600 128.400 ;
        RECT 534.000 127.600 536.600 128.400 ;
        RECT 537.200 128.200 537.800 129.000 ;
        RECT 538.800 129.400 539.600 129.600 ;
        RECT 538.800 129.000 544.200 129.400 ;
        RECT 538.800 128.800 545.000 129.000 ;
        RECT 543.600 128.200 545.000 128.800 ;
        RECT 537.200 127.600 543.000 128.200 ;
        RECT 546.000 128.000 547.600 128.800 ;
        RECT 546.000 127.600 546.600 128.000 ;
        RECT 534.000 122.200 534.800 127.000 ;
        RECT 537.200 122.200 538.000 127.000 ;
        RECT 542.400 126.800 546.600 127.600 ;
        RECT 548.400 127.400 549.200 133.000 ;
        RECT 547.200 126.800 549.200 127.400 ;
        RECT 538.800 122.200 539.600 125.000 ;
        RECT 540.400 122.200 541.200 125.000 ;
        RECT 543.600 122.200 544.400 126.800 ;
        RECT 547.200 126.200 547.800 126.800 ;
        RECT 546.800 125.600 547.800 126.200 ;
        RECT 546.800 122.200 547.600 125.600 ;
        RECT 1.200 115.800 2.000 119.800 ;
        RECT 1.400 115.600 2.000 115.800 ;
        RECT 4.400 115.800 5.200 119.800 ;
        RECT 4.400 115.600 5.000 115.800 ;
        RECT 1.400 115.000 5.000 115.600 ;
        RECT 1.400 112.400 2.000 115.000 ;
        RECT 2.800 114.300 3.600 114.400 ;
        RECT 6.000 114.300 6.800 114.400 ;
        RECT 2.800 113.700 6.800 114.300 ;
        RECT 2.800 112.800 3.600 113.700 ;
        RECT 6.000 113.600 6.800 113.700 ;
        RECT 1.200 111.600 2.000 112.400 ;
        RECT 4.400 112.300 5.200 112.400 ;
        RECT 6.000 112.300 6.800 112.400 ;
        RECT 4.400 111.700 6.800 112.300 ;
        RECT 4.400 111.600 5.200 111.700 ;
        RECT 1.400 108.400 2.000 111.600 ;
        RECT 6.000 110.800 6.800 111.700 ;
        RECT 3.600 109.600 5.200 110.400 ;
        RECT 1.400 108.200 3.000 108.400 ;
        RECT 1.400 107.800 3.200 108.200 ;
        RECT 2.400 102.200 3.200 107.800 ;
        RECT 7.600 106.800 8.400 108.400 ;
        RECT 9.200 106.200 10.000 119.800 ;
        RECT 12.400 115.800 13.200 119.800 ;
        RECT 12.600 115.600 13.200 115.800 ;
        RECT 15.600 115.600 16.400 119.800 ;
        RECT 18.800 115.800 19.600 119.800 ;
        RECT 19.000 115.600 19.600 115.800 ;
        RECT 22.000 115.800 22.800 119.800 ;
        RECT 26.800 115.800 27.600 119.800 ;
        RECT 22.000 115.600 22.600 115.800 ;
        RECT 12.600 115.000 16.200 115.600 ;
        RECT 19.000 115.000 22.600 115.600 ;
        RECT 27.000 115.600 27.600 115.800 ;
        RECT 30.000 115.800 30.800 119.800 ;
        RECT 30.000 115.600 30.600 115.800 ;
        RECT 27.000 115.000 30.600 115.600 ;
        RECT 10.800 111.600 11.600 113.200 ;
        RECT 12.600 112.400 13.200 115.000 ;
        RECT 14.000 112.800 14.800 114.400 ;
        RECT 19.000 112.400 19.600 115.000 ;
        RECT 20.400 112.800 21.200 114.400 ;
        RECT 28.400 112.800 29.200 114.400 ;
        RECT 30.000 112.400 30.600 115.000 ;
        RECT 32.400 113.600 33.200 114.400 ;
        RECT 32.400 112.400 33.000 113.600 ;
        RECT 33.800 112.400 34.600 119.800 ;
        RECT 12.400 111.600 13.200 112.400 ;
        RECT 12.600 108.400 13.200 111.600 ;
        RECT 17.200 110.800 18.000 112.400 ;
        RECT 18.800 111.600 19.600 112.400 ;
        RECT 14.800 109.600 16.400 110.400 ;
        RECT 19.000 108.400 19.600 111.600 ;
        RECT 23.600 110.800 24.400 112.400 ;
        RECT 25.200 110.800 26.000 112.400 ;
        RECT 30.000 111.600 30.800 112.400 ;
        RECT 31.600 111.800 33.000 112.400 ;
        RECT 33.600 111.800 34.600 112.400 ;
        RECT 31.600 111.600 32.400 111.800 ;
        RECT 21.200 109.600 22.800 110.400 ;
        RECT 26.800 109.600 28.400 110.400 ;
        RECT 30.000 108.400 30.600 111.600 ;
        RECT 33.600 108.400 34.200 111.800 ;
        RECT 34.800 110.300 35.600 110.400 ;
        RECT 36.400 110.300 37.200 110.400 ;
        RECT 39.600 110.300 40.400 119.800 ;
        RECT 44.400 112.000 45.200 119.800 ;
        RECT 47.600 115.200 48.400 119.800 ;
        RECT 34.800 109.700 40.400 110.300 ;
        RECT 34.800 108.800 35.600 109.700 ;
        RECT 36.400 109.600 37.200 109.700 ;
        RECT 12.600 108.200 14.200 108.400 ;
        RECT 19.000 108.200 20.600 108.400 ;
        RECT 29.000 108.200 30.600 108.400 ;
        RECT 12.600 107.800 14.400 108.200 ;
        RECT 19.000 107.800 20.800 108.200 ;
        RECT 9.200 105.600 11.000 106.200 ;
        RECT 10.200 104.400 11.000 105.600 ;
        RECT 9.200 103.600 11.000 104.400 ;
        RECT 10.200 102.200 11.000 103.600 ;
        RECT 13.600 102.200 14.400 107.800 ;
        RECT 20.000 102.200 20.800 107.800 ;
        RECT 28.800 107.800 30.600 108.200 ;
        RECT 28.800 102.200 29.600 107.800 ;
        RECT 31.600 107.600 34.200 108.400 ;
        RECT 36.400 108.200 37.200 108.400 ;
        RECT 35.600 107.600 37.200 108.200 ;
        RECT 31.800 106.200 32.400 107.600 ;
        RECT 35.600 107.200 36.400 107.600 ;
        RECT 33.400 106.200 37.000 106.600 ;
        RECT 31.600 102.200 32.400 106.200 ;
        RECT 33.200 106.000 37.200 106.200 ;
        RECT 33.200 102.200 34.000 106.000 ;
        RECT 36.400 102.200 37.200 106.000 ;
        RECT 39.600 102.200 40.400 109.700 ;
        RECT 44.200 111.200 45.200 112.000 ;
        RECT 45.800 114.600 48.400 115.200 ;
        RECT 45.800 113.000 46.400 114.600 ;
        RECT 50.800 114.400 51.600 119.800 ;
        RECT 54.000 117.000 54.800 119.800 ;
        RECT 55.600 117.000 56.400 119.800 ;
        RECT 57.200 117.000 58.000 119.800 ;
        RECT 52.200 114.400 56.400 115.200 ;
        RECT 49.000 113.600 51.600 114.400 ;
        RECT 58.800 113.600 59.600 119.800 ;
        RECT 62.000 115.000 62.800 119.800 ;
        RECT 65.200 115.000 66.000 119.800 ;
        RECT 66.800 117.000 67.600 119.800 ;
        RECT 68.400 117.000 69.200 119.800 ;
        RECT 71.600 115.200 72.400 119.800 ;
        RECT 74.800 116.400 75.600 119.800 ;
        RECT 74.800 115.800 75.800 116.400 ;
        RECT 75.200 115.200 75.800 115.800 ;
        RECT 70.400 114.400 74.600 115.200 ;
        RECT 75.200 114.600 77.200 115.200 ;
        RECT 62.000 113.600 64.600 114.400 ;
        RECT 65.200 113.800 71.000 114.400 ;
        RECT 74.000 114.000 74.600 114.400 ;
        RECT 54.000 113.000 54.800 113.200 ;
        RECT 45.800 112.400 54.800 113.000 ;
        RECT 57.200 113.000 58.000 113.200 ;
        RECT 65.200 113.000 65.800 113.800 ;
        RECT 71.600 113.200 73.000 113.800 ;
        RECT 74.000 113.200 75.600 114.000 ;
        RECT 57.200 112.400 65.800 113.000 ;
        RECT 66.800 113.000 73.000 113.200 ;
        RECT 66.800 112.600 72.200 113.000 ;
        RECT 66.800 112.400 67.600 112.600 ;
        RECT 41.200 106.800 42.000 108.400 ;
        RECT 44.200 106.800 45.000 111.200 ;
        RECT 45.800 110.600 46.400 112.400 ;
        RECT 45.600 110.000 46.400 110.600 ;
        RECT 52.400 110.000 75.800 110.600 ;
        RECT 45.600 108.000 46.200 110.000 ;
        RECT 52.400 109.400 53.200 110.000 ;
        RECT 70.000 109.600 70.800 110.000 ;
        RECT 75.000 109.800 75.800 110.000 ;
        RECT 46.800 108.600 50.600 109.400 ;
        RECT 45.600 107.400 46.800 108.000 ;
        RECT 44.200 106.000 45.200 106.800 ;
        RECT 44.400 102.200 45.200 106.000 ;
        RECT 46.000 102.200 46.800 107.400 ;
        RECT 49.800 107.400 50.600 108.600 ;
        RECT 49.800 106.800 51.600 107.400 ;
        RECT 50.800 106.200 51.600 106.800 ;
        RECT 55.600 106.400 56.400 109.200 ;
        RECT 58.800 108.600 62.000 109.400 ;
        RECT 65.800 108.600 67.800 109.400 ;
        RECT 76.400 109.000 77.200 114.600 ;
        RECT 80.600 112.400 81.400 119.800 ;
        RECT 86.000 116.400 86.800 119.800 ;
        RECT 85.800 115.800 86.800 116.400 ;
        RECT 85.800 115.200 86.400 115.800 ;
        RECT 89.200 115.200 90.000 119.800 ;
        RECT 92.400 117.000 93.200 119.800 ;
        RECT 94.000 117.000 94.800 119.800 ;
        RECT 84.400 114.600 86.400 115.200 ;
        RECT 82.000 113.600 82.800 114.400 ;
        RECT 82.200 112.400 82.800 113.600 ;
        RECT 80.600 111.800 81.600 112.400 ;
        RECT 82.200 111.800 83.600 112.400 ;
        RECT 58.400 107.800 59.200 108.000 ;
        RECT 58.400 107.200 62.800 107.800 ;
        RECT 62.000 107.000 62.800 107.200 ;
        RECT 63.600 106.800 64.400 108.400 ;
        RECT 50.800 105.400 53.200 106.200 ;
        RECT 55.600 105.600 56.600 106.400 ;
        RECT 59.600 105.600 61.200 106.400 ;
        RECT 62.000 106.200 62.800 106.400 ;
        RECT 65.800 106.200 66.600 108.600 ;
        RECT 68.400 108.200 77.200 109.000 ;
        RECT 79.600 108.800 80.400 110.400 ;
        RECT 81.000 108.400 81.600 111.800 ;
        RECT 82.800 111.600 83.600 111.800 ;
        RECT 84.400 109.000 85.200 114.600 ;
        RECT 87.000 114.400 91.200 115.200 ;
        RECT 95.600 115.000 96.400 119.800 ;
        RECT 98.800 115.000 99.600 119.800 ;
        RECT 87.000 114.000 87.600 114.400 ;
        RECT 86.000 113.200 87.600 114.000 ;
        RECT 90.600 113.800 96.400 114.400 ;
        RECT 88.600 113.200 90.000 113.800 ;
        RECT 88.600 113.000 94.800 113.200 ;
        RECT 89.400 112.600 94.800 113.000 ;
        RECT 94.000 112.400 94.800 112.600 ;
        RECT 95.800 113.000 96.400 113.800 ;
        RECT 97.000 113.600 99.600 114.400 ;
        RECT 102.000 113.600 102.800 119.800 ;
        RECT 103.600 117.000 104.400 119.800 ;
        RECT 105.200 117.000 106.000 119.800 ;
        RECT 106.800 117.000 107.600 119.800 ;
        RECT 105.200 114.400 109.400 115.200 ;
        RECT 110.000 114.400 110.800 119.800 ;
        RECT 113.200 115.200 114.000 119.800 ;
        RECT 113.200 114.600 115.800 115.200 ;
        RECT 110.000 113.600 112.600 114.400 ;
        RECT 103.600 113.000 104.400 113.200 ;
        RECT 95.800 112.400 104.400 113.000 ;
        RECT 106.800 113.000 107.600 113.200 ;
        RECT 115.200 113.000 115.800 114.600 ;
        RECT 106.800 112.400 115.800 113.000 ;
        RECT 115.200 110.600 115.800 112.400 ;
        RECT 116.400 112.000 117.200 119.800 ;
        RECT 116.400 111.200 117.400 112.000 ;
        RECT 85.800 110.000 109.200 110.600 ;
        RECT 115.200 110.000 116.000 110.600 ;
        RECT 85.800 109.800 86.600 110.000 ;
        RECT 87.600 109.600 88.400 110.000 ;
        RECT 90.800 109.600 91.600 110.000 ;
        RECT 108.400 109.400 109.200 110.000 ;
        RECT 71.800 106.800 74.800 107.600 ;
        RECT 71.800 106.200 72.600 106.800 ;
        RECT 62.000 105.600 66.600 106.200 ;
        RECT 52.400 102.200 53.200 105.400 ;
        RECT 70.000 105.400 72.600 106.200 ;
        RECT 54.000 102.200 54.800 105.000 ;
        RECT 55.600 102.200 56.400 105.000 ;
        RECT 57.200 102.200 58.000 105.000 ;
        RECT 58.800 102.200 59.600 105.000 ;
        RECT 62.000 102.200 62.800 105.000 ;
        RECT 65.200 102.200 66.000 105.000 ;
        RECT 66.800 102.200 67.600 105.000 ;
        RECT 68.400 102.200 69.200 105.000 ;
        RECT 70.000 102.200 70.800 105.400 ;
        RECT 76.400 102.200 77.200 108.200 ;
        RECT 78.000 108.200 78.800 108.400 ;
        RECT 78.000 107.600 79.600 108.200 ;
        RECT 81.000 107.600 83.600 108.400 ;
        RECT 84.400 108.200 93.200 109.000 ;
        RECT 93.800 108.600 95.800 109.400 ;
        RECT 99.600 108.600 102.800 109.400 ;
        RECT 78.800 107.200 79.600 107.600 ;
        RECT 78.200 106.200 81.800 106.600 ;
        RECT 82.800 106.200 83.400 107.600 ;
        RECT 78.000 106.000 82.000 106.200 ;
        RECT 78.000 102.200 78.800 106.000 ;
        RECT 81.200 102.200 82.000 106.000 ;
        RECT 82.800 102.200 83.600 106.200 ;
        RECT 84.400 102.200 85.200 108.200 ;
        RECT 86.800 106.800 89.800 107.600 ;
        RECT 89.000 106.200 89.800 106.800 ;
        RECT 95.000 106.200 95.800 108.600 ;
        RECT 97.200 106.800 98.000 108.400 ;
        RECT 102.400 107.800 103.200 108.000 ;
        RECT 98.800 107.200 103.200 107.800 ;
        RECT 98.800 107.000 99.600 107.200 ;
        RECT 105.200 106.400 106.000 109.200 ;
        RECT 111.000 108.600 114.800 109.400 ;
        RECT 111.000 107.400 111.800 108.600 ;
        RECT 115.400 108.000 116.000 110.000 ;
        RECT 98.800 106.200 99.600 106.400 ;
        RECT 89.000 105.400 91.600 106.200 ;
        RECT 95.000 105.600 99.600 106.200 ;
        RECT 100.400 105.600 102.000 106.400 ;
        RECT 105.000 105.600 106.000 106.400 ;
        RECT 110.000 106.800 111.800 107.400 ;
        RECT 114.800 107.400 116.000 108.000 ;
        RECT 110.000 106.200 110.800 106.800 ;
        RECT 90.800 102.200 91.600 105.400 ;
        RECT 108.400 105.400 110.800 106.200 ;
        RECT 92.400 102.200 93.200 105.000 ;
        RECT 94.000 102.200 94.800 105.000 ;
        RECT 95.600 102.200 96.400 105.000 ;
        RECT 98.800 102.200 99.600 105.000 ;
        RECT 102.000 102.200 102.800 105.000 ;
        RECT 103.600 102.200 104.400 105.000 ;
        RECT 105.200 102.200 106.000 105.000 ;
        RECT 106.800 102.200 107.600 105.000 ;
        RECT 108.400 102.200 109.200 105.400 ;
        RECT 114.800 102.200 115.600 107.400 ;
        RECT 116.600 106.800 117.400 111.200 ;
        RECT 116.400 106.000 117.400 106.800 ;
        RECT 116.400 102.200 117.200 106.000 ;
        RECT 119.600 102.200 120.400 119.800 ;
        RECT 129.800 112.600 130.600 119.800 ;
        RECT 129.800 111.800 131.600 112.600 ;
        RECT 134.000 111.800 134.800 119.800 ;
        RECT 135.600 112.400 136.400 119.800 ;
        RECT 138.800 112.400 139.600 119.800 ;
        RECT 135.600 111.800 139.600 112.400 ;
        RECT 130.800 111.600 131.600 111.800 ;
        RECT 127.600 110.300 128.400 110.400 ;
        RECT 129.200 110.300 130.000 111.200 ;
        RECT 127.600 109.700 130.000 110.300 ;
        RECT 127.600 109.600 128.400 109.700 ;
        RECT 129.200 109.600 130.000 109.700 ;
        RECT 130.800 108.400 131.400 111.600 ;
        RECT 134.200 110.400 134.800 111.800 ;
        RECT 138.000 110.400 138.800 110.800 ;
        RECT 134.000 109.800 136.400 110.400 ;
        RECT 138.000 109.800 139.600 110.400 ;
        RECT 134.000 109.600 134.800 109.800 ;
        RECT 130.800 107.600 131.600 108.400 ;
        RECT 121.200 106.300 122.000 106.400 ;
        RECT 129.200 106.300 130.000 106.400 ;
        RECT 121.200 105.700 130.000 106.300 ;
        RECT 121.200 104.800 122.000 105.700 ;
        RECT 129.200 105.600 130.000 105.700 ;
        RECT 130.800 104.200 131.400 107.600 ;
        RECT 132.400 104.800 133.200 106.400 ;
        RECT 134.000 105.600 134.800 106.400 ;
        RECT 135.800 106.200 136.400 109.800 ;
        RECT 138.800 109.600 139.600 109.800 ;
        RECT 137.200 107.600 138.000 109.200 ;
        RECT 134.200 104.800 135.000 105.600 ;
        RECT 130.800 102.200 131.600 104.200 ;
        RECT 135.600 102.200 136.400 106.200 ;
        RECT 140.400 104.800 141.200 106.400 ;
        RECT 142.000 106.300 142.800 119.800 ;
        RECT 144.200 112.600 145.000 119.800 ;
        RECT 144.200 111.800 146.000 112.600 ;
        RECT 151.000 112.400 151.800 119.800 ;
        RECT 152.400 113.600 153.200 114.400 ;
        RECT 152.600 112.400 153.200 113.600 ;
        RECT 154.800 112.400 155.600 119.800 ;
        RECT 158.000 112.400 158.800 119.800 ;
        RECT 151.000 111.800 152.000 112.400 ;
        RECT 152.600 111.800 154.000 112.400 ;
        RECT 154.800 111.800 158.800 112.400 ;
        RECT 159.600 111.800 160.400 119.800 ;
        RECT 163.800 112.600 164.600 119.800 ;
        RECT 162.800 111.800 164.600 112.600 ;
        RECT 168.600 112.400 169.400 119.800 ;
        RECT 170.000 113.600 170.800 114.400 ;
        RECT 170.200 112.400 170.800 113.600 ;
        RECT 143.600 109.600 144.400 111.200 ;
        RECT 145.200 110.300 145.800 111.800 ;
        RECT 148.400 110.300 149.200 110.400 ;
        RECT 145.200 109.700 149.200 110.300 ;
        RECT 145.200 108.400 145.800 109.700 ;
        RECT 148.400 109.600 149.200 109.700 ;
        RECT 150.000 108.800 150.800 110.400 ;
        RECT 151.400 108.400 152.000 111.800 ;
        RECT 153.200 111.600 154.000 111.800 ;
        RECT 155.600 110.400 156.400 110.800 ;
        RECT 159.600 110.400 160.200 111.800 ;
        RECT 154.800 109.800 156.400 110.400 ;
        RECT 158.000 109.800 160.400 110.400 ;
        RECT 154.800 109.600 155.600 109.800 ;
        RECT 145.200 107.600 146.000 108.400 ;
        RECT 148.400 108.200 149.200 108.400 ;
        RECT 148.400 107.600 150.000 108.200 ;
        RECT 151.400 107.600 154.000 108.400 ;
        RECT 154.800 108.300 155.600 108.400 ;
        RECT 156.400 108.300 157.200 109.200 ;
        RECT 154.800 107.700 157.200 108.300 ;
        RECT 154.800 107.600 155.600 107.700 ;
        RECT 156.400 107.600 157.200 107.700 ;
        RECT 143.600 106.300 144.400 106.400 ;
        RECT 142.000 105.700 144.400 106.300 ;
        RECT 142.000 102.200 142.800 105.700 ;
        RECT 143.600 105.600 144.400 105.700 ;
        RECT 145.200 104.200 145.800 107.600 ;
        RECT 149.200 107.200 150.000 107.600 ;
        RECT 146.800 104.800 147.600 106.400 ;
        RECT 148.600 106.200 152.200 106.600 ;
        RECT 153.200 106.200 153.800 107.600 ;
        RECT 158.000 106.200 158.600 109.800 ;
        RECT 159.600 109.600 160.400 109.800 ;
        RECT 163.000 108.400 163.600 111.800 ;
        RECT 167.600 111.600 169.600 112.400 ;
        RECT 170.200 111.800 171.600 112.400 ;
        RECT 170.800 111.600 171.600 111.800 ;
        RECT 164.400 109.600 165.200 111.200 ;
        RECT 167.600 108.800 168.400 110.400 ;
        RECT 169.000 108.400 169.600 111.600 ;
        RECT 170.800 110.300 171.600 110.400 ;
        RECT 172.400 110.300 173.200 119.800 ;
        RECT 170.800 109.700 173.200 110.300 ;
        RECT 170.800 109.600 171.600 109.700 ;
        RECT 162.800 108.300 163.600 108.400 ;
        RECT 166.000 108.300 166.800 108.400 ;
        RECT 162.800 108.200 166.800 108.300 ;
        RECT 162.800 107.700 167.600 108.200 ;
        RECT 162.800 107.600 163.600 107.700 ;
        RECT 166.000 107.600 167.600 107.700 ;
        RECT 169.000 107.600 171.600 108.400 ;
        RECT 148.400 106.000 152.400 106.200 ;
        RECT 145.200 102.200 146.000 104.200 ;
        RECT 148.400 102.200 149.200 106.000 ;
        RECT 151.600 102.200 152.400 106.000 ;
        RECT 153.200 102.200 154.000 106.200 ;
        RECT 158.000 102.200 158.800 106.200 ;
        RECT 159.600 105.600 160.400 106.400 ;
        RECT 159.400 104.800 160.200 105.600 ;
        RECT 161.200 104.800 162.000 106.400 ;
        RECT 163.000 104.200 163.600 107.600 ;
        RECT 166.800 107.200 167.600 107.600 ;
        RECT 166.200 106.200 169.800 106.600 ;
        RECT 170.800 106.200 171.400 107.600 ;
        RECT 162.800 102.200 163.600 104.200 ;
        RECT 166.000 106.000 170.000 106.200 ;
        RECT 166.000 102.200 166.800 106.000 ;
        RECT 169.200 102.200 170.000 106.000 ;
        RECT 170.800 102.200 171.600 106.200 ;
        RECT 172.400 102.200 173.200 109.700 ;
        RECT 175.600 106.800 176.400 108.400 ;
        RECT 174.000 104.800 174.800 106.400 ;
        RECT 177.200 106.200 178.000 119.800 ;
        RECT 182.000 116.400 182.800 119.800 ;
        RECT 181.800 115.800 182.800 116.400 ;
        RECT 181.800 115.200 182.400 115.800 ;
        RECT 185.200 115.200 186.000 119.800 ;
        RECT 188.400 117.000 189.200 119.800 ;
        RECT 190.000 117.000 190.800 119.800 ;
        RECT 180.400 114.600 182.400 115.200 ;
        RECT 178.800 111.600 179.600 113.200 ;
        RECT 180.400 109.000 181.200 114.600 ;
        RECT 183.000 114.400 187.200 115.200 ;
        RECT 191.600 115.000 192.400 119.800 ;
        RECT 194.800 115.000 195.600 119.800 ;
        RECT 183.000 114.000 183.600 114.400 ;
        RECT 182.000 113.200 183.600 114.000 ;
        RECT 186.600 113.800 192.400 114.400 ;
        RECT 184.600 113.200 186.000 113.800 ;
        RECT 184.600 113.000 190.800 113.200 ;
        RECT 185.400 112.600 190.800 113.000 ;
        RECT 190.000 112.400 190.800 112.600 ;
        RECT 191.800 113.000 192.400 113.800 ;
        RECT 193.000 113.600 195.600 114.400 ;
        RECT 198.000 113.600 198.800 119.800 ;
        RECT 199.600 117.000 200.400 119.800 ;
        RECT 201.200 117.000 202.000 119.800 ;
        RECT 202.800 117.000 203.600 119.800 ;
        RECT 201.200 114.400 205.400 115.200 ;
        RECT 206.000 114.400 206.800 119.800 ;
        RECT 209.200 115.200 210.000 119.800 ;
        RECT 209.200 114.600 211.800 115.200 ;
        RECT 206.000 113.600 208.600 114.400 ;
        RECT 199.600 113.000 200.400 113.200 ;
        RECT 191.800 112.400 200.400 113.000 ;
        RECT 202.800 113.000 203.600 113.200 ;
        RECT 211.200 113.000 211.800 114.600 ;
        RECT 202.800 112.400 211.800 113.000 ;
        RECT 211.200 110.600 211.800 112.400 ;
        RECT 212.400 112.000 213.200 119.800 ;
        RECT 212.400 111.200 213.400 112.000 ;
        RECT 215.600 111.800 216.400 119.800 ;
        RECT 217.200 112.400 218.000 119.800 ;
        RECT 220.400 112.400 221.200 119.800 ;
        RECT 217.200 111.800 221.200 112.400 ;
        RECT 181.800 110.000 205.200 110.600 ;
        RECT 211.200 110.000 212.000 110.600 ;
        RECT 181.800 109.800 182.600 110.000 ;
        RECT 183.600 109.600 184.400 110.000 ;
        RECT 186.800 109.600 187.600 110.000 ;
        RECT 204.400 109.400 205.200 110.000 ;
        RECT 180.400 108.200 189.200 109.000 ;
        RECT 189.800 108.600 191.800 109.400 ;
        RECT 195.600 108.600 198.800 109.400 ;
        RECT 177.200 105.600 179.000 106.200 ;
        RECT 178.200 102.200 179.000 105.600 ;
        RECT 180.400 102.200 181.200 108.200 ;
        RECT 182.800 106.800 185.800 107.600 ;
        RECT 185.000 106.200 185.800 106.800 ;
        RECT 191.000 106.200 191.800 108.600 ;
        RECT 193.200 106.800 194.000 108.400 ;
        RECT 198.400 107.800 199.200 108.000 ;
        RECT 194.800 107.200 199.200 107.800 ;
        RECT 194.800 107.000 195.600 107.200 ;
        RECT 201.200 106.400 202.000 109.200 ;
        RECT 207.000 108.600 210.800 109.400 ;
        RECT 207.000 107.400 207.800 108.600 ;
        RECT 211.400 108.000 212.000 110.000 ;
        RECT 194.800 106.200 195.600 106.400 ;
        RECT 185.000 105.400 187.600 106.200 ;
        RECT 191.000 105.600 195.600 106.200 ;
        RECT 196.400 105.600 198.000 106.400 ;
        RECT 201.000 105.600 202.000 106.400 ;
        RECT 206.000 106.800 207.800 107.400 ;
        RECT 210.800 107.400 212.000 108.000 ;
        RECT 206.000 106.200 206.800 106.800 ;
        RECT 186.800 102.200 187.600 105.400 ;
        RECT 204.400 105.400 206.800 106.200 ;
        RECT 188.400 102.200 189.200 105.000 ;
        RECT 190.000 102.200 190.800 105.000 ;
        RECT 191.600 102.200 192.400 105.000 ;
        RECT 194.800 102.200 195.600 105.000 ;
        RECT 198.000 102.200 198.800 105.000 ;
        RECT 199.600 102.200 200.400 105.000 ;
        RECT 201.200 102.200 202.000 105.000 ;
        RECT 202.800 102.200 203.600 105.000 ;
        RECT 204.400 102.200 205.200 105.400 ;
        RECT 210.800 102.200 211.600 107.400 ;
        RECT 212.600 106.800 213.400 111.200 ;
        RECT 215.800 110.400 216.400 111.800 ;
        RECT 222.000 111.600 222.800 113.200 ;
        RECT 219.600 110.400 220.400 110.800 ;
        RECT 215.600 109.800 218.000 110.400 ;
        RECT 219.600 109.800 221.200 110.400 ;
        RECT 215.600 109.600 216.400 109.800 ;
        RECT 215.600 108.300 216.400 108.400 ;
        RECT 217.400 108.300 218.000 109.800 ;
        RECT 220.400 109.600 221.200 109.800 ;
        RECT 215.600 107.700 218.000 108.300 ;
        RECT 215.600 107.600 216.400 107.700 ;
        RECT 212.400 106.000 213.400 106.800 ;
        RECT 214.000 106.300 214.800 106.400 ;
        RECT 215.600 106.300 216.400 106.400 ;
        RECT 212.400 102.200 213.200 106.000 ;
        RECT 214.000 105.700 216.400 106.300 ;
        RECT 217.400 106.200 218.000 107.700 ;
        RECT 218.800 108.300 219.600 109.200 ;
        RECT 223.600 108.300 224.400 119.800 ;
        RECT 227.600 113.600 228.400 114.400 ;
        RECT 227.600 112.400 228.200 113.600 ;
        RECT 229.000 112.400 229.800 119.800 ;
        RECT 235.800 112.600 236.600 119.800 ;
        RECT 226.800 111.800 228.200 112.400 ;
        RECT 228.800 111.800 229.800 112.400 ;
        RECT 234.800 111.800 236.600 112.600 ;
        RECT 226.800 111.600 227.600 111.800 ;
        RECT 225.200 110.300 226.000 110.400 ;
        RECT 228.800 110.300 229.400 111.800 ;
        RECT 225.200 109.700 229.400 110.300 ;
        RECT 225.200 109.600 226.000 109.700 ;
        RECT 228.800 108.400 229.400 109.700 ;
        RECT 230.000 110.300 230.800 110.400 ;
        RECT 235.000 110.300 235.600 111.800 ;
        RECT 230.000 109.700 235.600 110.300 ;
        RECT 230.000 108.800 230.800 109.700 ;
        RECT 235.000 108.400 235.600 109.700 ;
        RECT 236.400 109.600 237.200 111.200 ;
        RECT 218.800 107.700 224.400 108.300 ;
        RECT 218.800 107.600 219.600 107.700 ;
        RECT 223.600 106.200 224.400 107.700 ;
        RECT 225.200 106.800 226.000 108.400 ;
        RECT 226.800 107.600 229.400 108.400 ;
        RECT 231.600 108.300 232.400 108.400 ;
        RECT 233.200 108.300 234.000 108.400 ;
        RECT 231.600 108.200 234.000 108.300 ;
        RECT 230.800 107.700 234.000 108.200 ;
        RECT 230.800 107.600 232.400 107.700 ;
        RECT 233.200 107.600 234.000 107.700 ;
        RECT 234.800 107.600 235.600 108.400 ;
        RECT 227.000 106.200 227.600 107.600 ;
        RECT 230.800 107.200 231.600 107.600 ;
        RECT 228.600 106.200 232.200 106.600 ;
        RECT 214.000 105.600 214.800 105.700 ;
        RECT 215.600 105.600 216.400 105.700 ;
        RECT 215.800 104.800 216.600 105.600 ;
        RECT 217.200 102.200 218.000 106.200 ;
        RECT 222.600 105.600 224.400 106.200 ;
        RECT 222.600 102.200 223.400 105.600 ;
        RECT 226.800 102.200 227.600 106.200 ;
        RECT 228.400 106.000 232.400 106.200 ;
        RECT 228.400 102.200 229.200 106.000 ;
        RECT 231.600 102.200 232.400 106.000 ;
        RECT 233.200 104.800 234.000 106.400 ;
        RECT 235.000 104.200 235.600 107.600 ;
        RECT 236.400 106.300 237.200 106.400 ;
        RECT 238.000 106.300 238.800 119.800 ;
        RECT 241.200 111.200 242.000 119.800 ;
        RECT 245.400 112.400 246.200 119.800 ;
        RECT 248.400 113.600 249.200 114.400 ;
        RECT 248.400 112.400 249.000 113.600 ;
        RECT 249.800 112.400 250.600 119.800 ;
        RECT 245.400 111.800 246.800 112.400 ;
        RECT 241.200 110.800 245.200 111.200 ;
        RECT 241.200 110.600 245.400 110.800 ;
        RECT 244.600 110.000 245.400 110.600 ;
        RECT 246.200 110.400 246.800 111.800 ;
        RECT 247.600 111.800 249.000 112.400 ;
        RECT 249.600 111.800 250.600 112.400 ;
        RECT 256.600 112.400 257.400 119.800 ;
        RECT 258.000 113.600 258.800 114.400 ;
        RECT 258.200 112.400 258.800 113.600 ;
        RECT 260.400 112.400 261.200 119.800 ;
        RECT 263.600 112.400 264.400 119.800 ;
        RECT 256.600 111.800 257.600 112.400 ;
        RECT 258.200 111.800 259.600 112.400 ;
        RECT 260.400 111.800 264.400 112.400 ;
        RECT 265.200 111.800 266.000 119.800 ;
        RECT 274.800 112.000 275.600 119.800 ;
        RECT 278.000 115.200 278.800 119.800 ;
        RECT 247.600 111.600 248.400 111.800 ;
        RECT 243.200 108.400 244.000 109.200 ;
        RECT 242.800 107.600 243.800 108.400 ;
        RECT 244.800 107.000 245.400 110.000 ;
        RECT 246.000 109.600 246.800 110.400 ;
        RECT 246.200 108.400 246.800 109.600 ;
        RECT 249.600 108.400 250.200 111.800 ;
        RECT 250.800 108.800 251.600 110.400 ;
        RECT 252.400 110.300 253.200 110.400 ;
        RECT 255.600 110.300 256.400 110.400 ;
        RECT 252.400 109.700 256.400 110.300 ;
        RECT 252.400 109.600 253.200 109.700 ;
        RECT 255.600 108.800 256.400 109.700 ;
        RECT 257.000 110.300 257.600 111.800 ;
        RECT 258.800 111.600 259.600 111.800 ;
        RECT 261.200 110.400 262.000 110.800 ;
        RECT 265.200 110.400 265.800 111.800 ;
        RECT 274.600 111.200 275.600 112.000 ;
        RECT 276.200 114.600 278.800 115.200 ;
        RECT 276.200 113.000 276.800 114.600 ;
        RECT 281.200 114.400 282.000 119.800 ;
        RECT 284.400 117.000 285.200 119.800 ;
        RECT 286.000 117.000 286.800 119.800 ;
        RECT 287.600 117.000 288.400 119.800 ;
        RECT 282.600 114.400 286.800 115.200 ;
        RECT 279.400 113.600 282.000 114.400 ;
        RECT 289.200 113.600 290.000 119.800 ;
        RECT 292.400 115.000 293.200 119.800 ;
        RECT 295.600 115.000 296.400 119.800 ;
        RECT 297.200 117.000 298.000 119.800 ;
        RECT 298.800 117.000 299.600 119.800 ;
        RECT 302.000 115.200 302.800 119.800 ;
        RECT 305.200 116.400 306.000 119.800 ;
        RECT 305.200 115.800 306.200 116.400 ;
        RECT 305.600 115.200 306.200 115.800 ;
        RECT 300.800 114.400 305.000 115.200 ;
        RECT 305.600 114.600 307.600 115.200 ;
        RECT 292.400 113.600 295.000 114.400 ;
        RECT 295.600 113.800 301.400 114.400 ;
        RECT 304.400 114.000 305.000 114.400 ;
        RECT 284.400 113.000 285.200 113.200 ;
        RECT 276.200 112.400 285.200 113.000 ;
        RECT 287.600 113.000 288.400 113.200 ;
        RECT 295.600 113.000 296.200 113.800 ;
        RECT 302.000 113.200 303.400 113.800 ;
        RECT 304.400 113.200 306.000 114.000 ;
        RECT 287.600 112.400 296.200 113.000 ;
        RECT 297.200 113.000 303.400 113.200 ;
        RECT 297.200 112.600 302.600 113.000 ;
        RECT 297.200 112.400 298.000 112.600 ;
        RECT 260.400 110.300 262.000 110.400 ;
        RECT 257.000 109.800 262.000 110.300 ;
        RECT 263.600 109.800 266.000 110.400 ;
        RECT 257.000 109.700 261.200 109.800 ;
        RECT 257.000 108.400 257.600 109.700 ;
        RECT 260.400 109.600 261.200 109.700 ;
        RECT 246.000 107.600 246.800 108.400 ;
        RECT 247.600 107.600 250.200 108.400 ;
        RECT 252.400 108.200 253.200 108.400 ;
        RECT 251.600 107.600 253.200 108.200 ;
        RECT 254.000 108.200 254.800 108.400 ;
        RECT 254.000 107.600 255.600 108.200 ;
        RECT 257.000 107.600 259.600 108.400 ;
        RECT 262.000 107.600 262.800 109.200 ;
        RECT 243.000 106.400 245.400 107.000 ;
        RECT 236.400 105.700 238.800 106.300 ;
        RECT 236.400 105.600 237.200 105.700 ;
        RECT 234.800 102.200 235.600 104.200 ;
        RECT 238.000 102.200 238.800 105.700 ;
        RECT 239.600 104.800 240.400 106.400 ;
        RECT 241.200 104.800 242.000 106.400 ;
        RECT 243.000 104.200 243.600 106.400 ;
        RECT 246.200 106.200 246.800 107.600 ;
        RECT 247.800 106.200 248.400 107.600 ;
        RECT 251.600 107.200 252.400 107.600 ;
        RECT 254.800 107.200 255.600 107.600 ;
        RECT 249.400 106.200 253.000 106.600 ;
        RECT 254.200 106.200 257.800 106.600 ;
        RECT 258.800 106.200 259.400 107.600 ;
        RECT 263.600 106.200 264.200 109.800 ;
        RECT 265.200 109.600 266.000 109.800 ;
        RECT 274.600 106.800 275.400 111.200 ;
        RECT 276.200 110.600 276.800 112.400 ;
        RECT 300.200 111.800 301.200 112.000 ;
        RECT 303.600 111.800 304.400 112.400 ;
        RECT 277.400 111.200 304.400 111.800 ;
        RECT 277.400 111.000 278.200 111.200 ;
        RECT 276.000 110.000 276.800 110.600 ;
        RECT 276.000 108.000 276.600 110.000 ;
        RECT 277.200 108.600 281.000 109.400 ;
        RECT 276.000 107.400 277.200 108.000 ;
        RECT 265.200 106.300 266.000 106.400 ;
        RECT 266.800 106.300 267.600 106.400 ;
        RECT 242.800 102.200 243.600 104.200 ;
        RECT 246.000 102.200 246.800 106.200 ;
        RECT 247.600 102.200 248.400 106.200 ;
        RECT 249.200 106.000 253.200 106.200 ;
        RECT 249.200 102.200 250.000 106.000 ;
        RECT 252.400 102.200 253.200 106.000 ;
        RECT 254.000 106.000 258.000 106.200 ;
        RECT 254.000 102.200 254.800 106.000 ;
        RECT 257.200 102.200 258.000 106.000 ;
        RECT 258.800 102.200 259.600 106.200 ;
        RECT 263.600 102.200 264.400 106.200 ;
        RECT 265.200 105.700 267.600 106.300 ;
        RECT 274.600 106.000 275.600 106.800 ;
        RECT 265.200 105.600 266.000 105.700 ;
        RECT 266.800 105.600 267.600 105.700 ;
        RECT 265.000 104.800 265.800 105.600 ;
        RECT 274.800 102.200 275.600 106.000 ;
        RECT 276.400 102.200 277.200 107.400 ;
        RECT 280.200 107.400 281.000 108.600 ;
        RECT 280.200 106.800 282.000 107.400 ;
        RECT 281.200 106.200 282.000 106.800 ;
        RECT 286.000 106.400 286.800 109.200 ;
        RECT 289.200 108.600 292.400 109.400 ;
        RECT 296.200 108.600 298.200 109.400 ;
        RECT 306.800 109.000 307.600 114.600 ;
        RECT 311.000 112.400 311.800 119.800 ;
        RECT 312.400 113.600 313.200 114.400 ;
        RECT 312.600 112.400 313.200 113.600 ;
        RECT 315.600 113.600 316.400 114.400 ;
        RECT 315.600 112.400 316.200 113.600 ;
        RECT 317.000 112.400 317.800 119.800 ;
        RECT 311.000 111.800 312.000 112.400 ;
        RECT 312.600 111.800 314.000 112.400 ;
        RECT 288.800 107.800 289.600 108.000 ;
        RECT 288.800 107.200 293.200 107.800 ;
        RECT 292.400 107.000 293.200 107.200 ;
        RECT 294.000 106.800 294.800 108.400 ;
        RECT 281.200 105.400 283.600 106.200 ;
        RECT 286.000 105.600 287.000 106.400 ;
        RECT 290.000 105.600 291.600 106.400 ;
        RECT 292.400 106.200 293.200 106.400 ;
        RECT 296.200 106.200 297.000 108.600 ;
        RECT 298.800 108.200 307.600 109.000 ;
        RECT 311.400 110.300 312.000 111.800 ;
        RECT 313.200 111.600 314.000 111.800 ;
        RECT 314.800 111.800 316.200 112.400 ;
        RECT 316.800 111.800 317.800 112.400 ;
        RECT 314.800 111.600 315.600 111.800 ;
        RECT 314.900 110.300 315.500 111.600 ;
        RECT 311.400 109.700 315.500 110.300 ;
        RECT 311.400 108.400 312.000 109.700 ;
        RECT 316.800 108.400 317.400 111.800 ;
        RECT 318.000 108.800 318.800 110.400 ;
        RECT 302.200 106.800 305.200 107.600 ;
        RECT 302.200 106.200 303.000 106.800 ;
        RECT 292.400 105.600 297.000 106.200 ;
        RECT 282.800 102.200 283.600 105.400 ;
        RECT 300.400 105.400 303.000 106.200 ;
        RECT 284.400 102.200 285.200 105.000 ;
        RECT 286.000 102.200 286.800 105.000 ;
        RECT 287.600 102.200 288.400 105.000 ;
        RECT 289.200 102.200 290.000 105.000 ;
        RECT 292.400 102.200 293.200 105.000 ;
        RECT 295.600 102.200 296.400 105.000 ;
        RECT 297.200 102.200 298.000 105.000 ;
        RECT 298.800 102.200 299.600 105.000 ;
        RECT 300.400 102.200 301.200 105.400 ;
        RECT 306.800 102.200 307.600 108.200 ;
        RECT 308.400 108.200 309.200 108.400 ;
        RECT 308.400 107.600 310.000 108.200 ;
        RECT 311.400 107.600 314.000 108.400 ;
        RECT 314.800 107.600 317.400 108.400 ;
        RECT 319.600 108.300 320.400 108.400 ;
        RECT 322.800 108.300 323.600 119.800 ;
        RECT 326.000 111.200 326.800 119.800 ;
        RECT 329.200 111.200 330.000 119.800 ;
        RECT 332.400 111.200 333.200 119.800 ;
        RECT 335.600 111.200 336.400 119.800 ;
        RECT 340.400 116.400 341.200 119.800 ;
        RECT 340.200 115.800 341.200 116.400 ;
        RECT 340.200 115.200 340.800 115.800 ;
        RECT 343.600 115.200 344.400 119.800 ;
        RECT 346.800 117.000 347.600 119.800 ;
        RECT 348.400 117.000 349.200 119.800 ;
        RECT 319.600 108.200 323.600 108.300 ;
        RECT 318.800 107.700 323.600 108.200 ;
        RECT 318.800 107.600 320.400 107.700 ;
        RECT 309.200 107.200 310.000 107.600 ;
        RECT 308.600 106.200 312.200 106.600 ;
        RECT 313.200 106.200 313.800 107.600 ;
        RECT 315.000 106.200 315.600 107.600 ;
        RECT 318.800 107.200 319.600 107.600 ;
        RECT 316.600 106.200 320.200 106.600 ;
        RECT 308.400 106.000 312.400 106.200 ;
        RECT 308.400 102.200 309.200 106.000 ;
        RECT 311.600 102.200 312.400 106.000 ;
        RECT 313.200 102.200 314.000 106.200 ;
        RECT 314.800 102.200 315.600 106.200 ;
        RECT 316.400 106.000 320.400 106.200 ;
        RECT 316.400 102.200 317.200 106.000 ;
        RECT 319.600 102.200 320.400 106.000 ;
        RECT 321.200 104.800 322.000 106.400 ;
        RECT 322.800 102.200 323.600 107.700 ;
        RECT 324.400 110.400 326.800 111.200 ;
        RECT 327.800 110.400 330.000 111.200 ;
        RECT 331.000 110.400 333.200 111.200 ;
        RECT 334.600 110.400 336.400 111.200 ;
        RECT 338.800 114.600 340.800 115.200 ;
        RECT 324.400 107.600 325.200 110.400 ;
        RECT 327.800 109.000 328.600 110.400 ;
        RECT 331.000 109.000 331.800 110.400 ;
        RECT 334.600 109.000 335.400 110.400 ;
        RECT 326.000 108.200 328.600 109.000 ;
        RECT 329.400 108.200 331.800 109.000 ;
        RECT 332.800 108.200 335.400 109.000 ;
        RECT 327.800 107.600 328.600 108.200 ;
        RECT 331.000 107.600 331.800 108.200 ;
        RECT 334.600 107.600 335.400 108.200 ;
        RECT 338.800 109.000 339.600 114.600 ;
        RECT 341.400 114.400 345.600 115.200 ;
        RECT 350.000 115.000 350.800 119.800 ;
        RECT 353.200 115.000 354.000 119.800 ;
        RECT 341.400 114.000 342.000 114.400 ;
        RECT 340.400 113.200 342.000 114.000 ;
        RECT 345.000 113.800 350.800 114.400 ;
        RECT 343.000 113.200 344.400 113.800 ;
        RECT 343.000 113.000 349.200 113.200 ;
        RECT 343.800 112.600 349.200 113.000 ;
        RECT 348.400 112.400 349.200 112.600 ;
        RECT 350.200 113.000 350.800 113.800 ;
        RECT 351.400 113.600 354.000 114.400 ;
        RECT 356.400 113.600 357.200 119.800 ;
        RECT 358.000 117.000 358.800 119.800 ;
        RECT 359.600 117.000 360.400 119.800 ;
        RECT 361.200 117.000 362.000 119.800 ;
        RECT 359.600 114.400 363.800 115.200 ;
        RECT 364.400 114.400 365.200 119.800 ;
        RECT 367.600 115.200 368.400 119.800 ;
        RECT 367.600 114.600 370.200 115.200 ;
        RECT 364.400 113.600 367.000 114.400 ;
        RECT 358.000 113.000 358.800 113.200 ;
        RECT 350.200 112.400 358.800 113.000 ;
        RECT 361.200 113.000 362.000 113.200 ;
        RECT 369.600 113.000 370.200 114.600 ;
        RECT 361.200 112.400 370.200 113.000 ;
        RECT 369.600 110.600 370.200 112.400 ;
        RECT 370.800 112.000 371.600 119.800 ;
        RECT 370.800 111.200 371.800 112.000 ;
        RECT 376.600 111.800 378.600 119.800 ;
        RECT 340.200 110.000 363.600 110.600 ;
        RECT 369.600 110.000 370.400 110.600 ;
        RECT 340.200 109.800 341.000 110.000 ;
        RECT 342.000 109.600 342.800 110.000 ;
        RECT 345.200 109.600 346.000 110.000 ;
        RECT 362.800 109.400 363.600 110.000 ;
        RECT 338.800 108.200 347.600 109.000 ;
        RECT 348.200 108.600 350.200 109.400 ;
        RECT 354.000 108.600 357.200 109.400 ;
        RECT 324.400 106.800 326.800 107.600 ;
        RECT 327.800 106.800 330.000 107.600 ;
        RECT 331.000 106.800 333.200 107.600 ;
        RECT 334.600 106.800 336.400 107.600 ;
        RECT 326.000 102.200 326.800 106.800 ;
        RECT 329.200 102.200 330.000 106.800 ;
        RECT 332.400 102.200 333.200 106.800 ;
        RECT 335.600 102.200 336.400 106.800 ;
        RECT 338.800 102.200 339.600 108.200 ;
        RECT 341.200 106.800 344.200 107.600 ;
        RECT 343.400 106.200 344.200 106.800 ;
        RECT 349.400 106.200 350.200 108.600 ;
        RECT 351.600 106.800 352.400 108.400 ;
        RECT 356.800 107.800 357.600 108.000 ;
        RECT 353.200 107.200 357.600 107.800 ;
        RECT 353.200 107.000 354.000 107.200 ;
        RECT 359.600 106.400 360.400 109.200 ;
        RECT 365.400 108.600 369.200 109.400 ;
        RECT 365.400 107.400 366.200 108.600 ;
        RECT 369.800 108.000 370.400 110.000 ;
        RECT 353.200 106.200 354.000 106.400 ;
        RECT 343.400 105.400 346.000 106.200 ;
        RECT 349.400 105.600 354.000 106.200 ;
        RECT 354.800 105.600 356.400 106.400 ;
        RECT 359.400 105.600 360.400 106.400 ;
        RECT 364.400 106.800 366.200 107.400 ;
        RECT 369.200 107.400 370.400 108.000 ;
        RECT 364.400 106.200 365.200 106.800 ;
        RECT 345.200 102.200 346.000 105.400 ;
        RECT 362.800 105.400 365.200 106.200 ;
        RECT 346.800 102.200 347.600 105.000 ;
        RECT 348.400 102.200 349.200 105.000 ;
        RECT 350.000 102.200 350.800 105.000 ;
        RECT 353.200 102.200 354.000 105.000 ;
        RECT 356.400 102.200 357.200 105.000 ;
        RECT 358.000 102.200 358.800 105.000 ;
        RECT 359.600 102.200 360.400 105.000 ;
        RECT 361.200 102.200 362.000 105.000 ;
        RECT 362.800 102.200 363.600 105.400 ;
        RECT 369.200 102.200 370.000 107.400 ;
        RECT 371.000 106.800 371.800 111.200 ;
        RECT 374.000 107.600 374.800 109.200 ;
        RECT 375.600 108.800 376.400 110.400 ;
        RECT 377.400 108.400 378.000 111.800 ;
        RECT 378.800 108.800 379.600 110.400 ;
        RECT 377.200 108.200 378.000 108.400 ;
        RECT 380.400 108.300 381.200 108.400 ;
        RECT 382.000 108.300 382.800 119.800 ;
        RECT 385.200 112.400 386.000 119.800 ;
        RECT 388.400 119.200 392.400 119.800 ;
        RECT 388.400 112.400 389.200 119.200 ;
        RECT 385.200 111.800 389.200 112.400 ;
        RECT 390.000 111.800 390.800 118.600 ;
        RECT 391.600 111.800 392.400 119.200 ;
        RECT 393.800 112.600 394.600 119.800 ;
        RECT 393.800 111.800 395.600 112.600 ;
        RECT 390.000 111.200 390.600 111.800 ;
        RECT 386.000 110.400 386.800 110.800 ;
        RECT 388.600 110.600 390.600 111.200 ;
        RECT 388.600 110.400 389.200 110.600 ;
        RECT 385.200 109.800 386.800 110.400 ;
        RECT 385.200 109.600 386.000 109.800 ;
        RECT 388.400 109.600 389.200 110.400 ;
        RECT 391.600 109.600 392.400 111.200 ;
        RECT 393.200 109.600 394.000 111.200 ;
        RECT 380.400 108.200 382.800 108.300 ;
        RECT 375.600 107.600 378.000 108.200 ;
        RECT 379.600 107.700 382.800 108.200 ;
        RECT 379.600 107.600 381.200 107.700 ;
        RECT 370.800 106.000 371.800 106.800 ;
        RECT 375.600 106.200 376.200 107.600 ;
        RECT 379.600 107.200 380.400 107.600 ;
        RECT 377.400 106.200 381.000 106.600 ;
        RECT 370.800 102.200 371.600 106.000 ;
        RECT 374.000 102.800 374.800 106.200 ;
        RECT 375.600 103.400 376.400 106.200 ;
        RECT 377.200 106.000 381.200 106.200 ;
        RECT 377.200 102.800 378.000 106.000 ;
        RECT 374.000 102.200 378.000 102.800 ;
        RECT 380.400 102.200 381.200 106.000 ;
        RECT 382.000 102.200 382.800 107.700 ;
        RECT 383.600 108.300 384.400 108.400 ;
        RECT 386.800 108.300 387.600 109.200 ;
        RECT 383.600 107.700 387.600 108.300 ;
        RECT 383.600 107.600 384.400 107.700 ;
        RECT 386.800 107.600 387.600 107.700 ;
        RECT 383.600 104.800 384.400 106.400 ;
        RECT 388.600 106.200 389.200 109.600 ;
        RECT 389.800 108.800 390.600 109.600 ;
        RECT 390.000 108.400 390.600 108.800 ;
        RECT 394.800 108.400 395.400 111.800 ;
        RECT 399.600 110.300 400.400 119.800 ;
        RECT 401.800 112.600 402.600 119.800 ;
        RECT 401.800 111.800 403.600 112.600 ;
        RECT 408.600 111.800 410.600 119.800 ;
        RECT 414.800 113.600 415.600 114.400 ;
        RECT 414.800 112.400 415.400 113.600 ;
        RECT 416.200 112.400 417.000 119.800 ;
        RECT 421.000 112.600 421.800 119.800 ;
        RECT 414.000 111.800 415.400 112.400 ;
        RECT 401.200 110.300 402.000 111.200 ;
        RECT 399.600 109.700 402.000 110.300 ;
        RECT 390.000 107.600 390.800 108.400 ;
        RECT 394.800 107.600 395.600 108.400 ;
        RECT 393.200 106.300 394.000 106.400 ;
        RECT 394.800 106.300 395.400 107.600 ;
        RECT 388.200 102.200 389.800 106.200 ;
        RECT 393.200 105.700 395.500 106.300 ;
        RECT 393.200 105.600 394.000 105.700 ;
        RECT 394.800 104.200 395.400 105.700 ;
        RECT 396.400 104.800 397.200 106.400 ;
        RECT 394.800 102.200 395.600 104.200 ;
        RECT 399.600 102.200 400.400 109.700 ;
        RECT 401.200 109.600 402.000 109.700 ;
        RECT 402.800 108.400 403.400 111.800 ;
        RECT 402.800 107.600 403.600 108.400 ;
        RECT 406.000 107.600 406.800 109.200 ;
        RECT 407.600 108.800 408.400 110.400 ;
        RECT 409.400 108.400 410.000 111.800 ;
        RECT 414.000 111.600 414.800 111.800 ;
        RECT 416.000 111.600 418.000 112.400 ;
        RECT 421.000 111.800 422.800 112.600 ;
        RECT 434.200 111.800 436.200 119.800 ;
        RECT 441.200 115.800 442.000 119.800 ;
        RECT 441.400 115.600 442.000 115.800 ;
        RECT 444.400 115.800 445.200 119.800 ;
        RECT 444.400 115.600 445.000 115.800 ;
        RECT 441.400 115.000 445.000 115.600 ;
        RECT 442.800 112.800 443.600 114.400 ;
        RECT 444.400 112.400 445.000 115.000 ;
        RECT 446.000 112.400 446.800 119.800 ;
        RECT 449.200 112.400 450.000 119.800 ;
        RECT 410.800 110.300 411.600 110.400 ;
        RECT 412.400 110.300 413.200 110.400 ;
        RECT 410.800 109.700 413.200 110.300 ;
        RECT 410.800 108.800 411.600 109.700 ;
        RECT 412.400 109.600 413.200 109.700 ;
        RECT 416.000 108.400 416.600 111.600 ;
        RECT 417.200 108.800 418.000 110.400 ;
        RECT 418.800 110.300 419.600 110.400 ;
        RECT 420.400 110.300 421.200 111.200 ;
        RECT 418.800 109.700 421.200 110.300 ;
        RECT 418.800 109.600 419.600 109.700 ;
        RECT 420.400 109.600 421.200 109.700 ;
        RECT 422.000 108.400 422.600 111.800 ;
        RECT 409.200 108.200 410.000 108.400 ;
        RECT 412.400 108.200 413.200 108.400 ;
        RECT 407.600 107.600 410.000 108.200 ;
        RECT 411.600 107.600 413.200 108.200 ;
        RECT 414.000 107.600 416.600 108.400 ;
        RECT 418.800 108.200 419.600 108.400 ;
        RECT 418.000 107.600 419.600 108.200 ;
        RECT 422.000 107.600 422.800 108.400 ;
        RECT 431.600 107.600 432.400 109.200 ;
        RECT 433.200 108.800 434.000 110.400 ;
        RECT 435.000 108.400 435.600 111.800 ;
        RECT 439.600 110.800 440.400 112.400 ;
        RECT 444.400 111.600 445.200 112.400 ;
        RECT 446.000 111.800 450.000 112.400 ;
        RECT 450.800 111.800 451.600 119.800 ;
        RECT 436.400 110.300 437.200 110.400 ;
        RECT 438.000 110.300 438.800 110.400 ;
        RECT 436.400 109.700 438.800 110.300 ;
        RECT 436.400 108.800 437.200 109.700 ;
        RECT 438.000 109.600 438.800 109.700 ;
        RECT 441.200 109.600 442.800 110.400 ;
        RECT 444.400 108.400 445.000 111.600 ;
        RECT 446.800 110.400 447.600 110.800 ;
        RECT 450.800 110.400 451.400 111.800 ;
        RECT 452.400 111.600 453.200 113.200 ;
        RECT 446.000 109.800 447.600 110.400 ;
        RECT 449.200 109.800 451.600 110.400 ;
        RECT 446.000 109.600 446.800 109.800 ;
        RECT 434.800 108.200 435.600 108.400 ;
        RECT 438.000 108.200 438.800 108.400 ;
        RECT 443.400 108.200 445.000 108.400 ;
        RECT 433.200 107.600 435.600 108.200 ;
        RECT 437.200 107.600 438.800 108.200 ;
        RECT 443.200 107.800 445.000 108.200 ;
        RECT 402.800 104.400 403.400 107.600 ;
        RECT 404.400 104.800 405.200 106.400 ;
        RECT 407.600 106.200 408.200 107.600 ;
        RECT 411.600 107.200 412.400 107.600 ;
        RECT 409.400 106.200 413.000 106.600 ;
        RECT 414.200 106.200 414.800 107.600 ;
        RECT 418.000 107.200 418.800 107.600 ;
        RECT 415.800 106.200 419.400 106.600 ;
        RECT 402.800 102.200 403.600 104.400 ;
        RECT 406.000 102.800 406.800 106.200 ;
        RECT 407.600 103.400 408.400 106.200 ;
        RECT 409.200 106.000 413.200 106.200 ;
        RECT 409.200 102.800 410.000 106.000 ;
        RECT 406.000 102.200 410.000 102.800 ;
        RECT 412.400 102.200 413.200 106.000 ;
        RECT 414.000 102.200 414.800 106.200 ;
        RECT 415.600 106.000 419.600 106.200 ;
        RECT 415.600 102.200 416.400 106.000 ;
        RECT 418.800 102.200 419.600 106.000 ;
        RECT 422.000 104.400 422.600 107.600 ;
        RECT 433.200 106.400 433.800 107.600 ;
        RECT 437.200 107.200 438.000 107.600 ;
        RECT 423.600 104.800 424.400 106.400 ;
        RECT 422.000 102.200 422.800 104.400 ;
        RECT 431.600 102.800 432.400 106.200 ;
        RECT 433.200 103.400 434.000 106.400 ;
        RECT 435.000 106.200 438.600 106.600 ;
        RECT 434.800 106.000 438.800 106.200 ;
        RECT 434.800 102.800 435.600 106.000 ;
        RECT 431.600 102.200 435.600 102.800 ;
        RECT 438.000 102.200 438.800 106.000 ;
        RECT 443.200 102.200 444.000 107.800 ;
        RECT 447.600 107.600 448.400 109.200 ;
        RECT 449.200 108.400 449.800 109.800 ;
        RECT 450.800 109.600 451.600 109.800 ;
        RECT 449.200 107.600 450.000 108.400 ;
        RECT 449.200 106.200 449.800 107.600 ;
        RECT 450.800 106.300 451.600 106.400 ;
        RECT 454.000 106.300 454.800 119.800 ;
        RECT 459.800 112.400 460.600 119.800 ;
        RECT 461.200 113.600 462.000 114.400 ;
        RECT 461.400 112.400 462.000 113.600 ;
        RECT 466.200 112.600 467.000 119.800 ;
        RECT 459.800 111.800 460.800 112.400 ;
        RECT 461.400 111.800 462.800 112.400 ;
        RECT 465.200 111.800 467.000 112.600 ;
        RECT 455.600 110.300 456.400 110.400 ;
        RECT 458.800 110.300 459.600 110.400 ;
        RECT 455.600 109.700 459.600 110.300 ;
        RECT 455.600 109.600 456.400 109.700 ;
        RECT 458.800 108.800 459.600 109.700 ;
        RECT 460.200 110.300 460.800 111.800 ;
        RECT 462.000 111.600 462.800 111.800 ;
        RECT 463.600 110.300 464.400 110.400 ;
        RECT 460.200 109.700 464.400 110.300 ;
        RECT 460.200 108.400 460.800 109.700 ;
        RECT 463.600 109.600 464.400 109.700 ;
        RECT 465.400 108.400 466.000 111.800 ;
        RECT 466.800 109.600 467.600 111.200 ;
        RECT 455.600 106.800 456.400 108.400 ;
        RECT 457.200 108.200 458.000 108.400 ;
        RECT 457.200 107.600 458.800 108.200 ;
        RECT 460.200 107.600 462.800 108.400 ;
        RECT 465.200 107.600 466.000 108.400 ;
        RECT 458.000 107.200 458.800 107.600 ;
        RECT 449.200 102.200 450.000 106.200 ;
        RECT 450.800 105.700 454.800 106.300 ;
        RECT 457.400 106.200 461.000 106.600 ;
        RECT 462.000 106.200 462.600 107.600 ;
        RECT 450.800 105.600 451.600 105.700 ;
        RECT 453.000 105.600 454.800 105.700 ;
        RECT 457.200 106.000 461.200 106.200 ;
        RECT 450.600 104.800 451.400 105.600 ;
        RECT 453.000 102.200 453.800 105.600 ;
        RECT 457.200 102.200 458.000 106.000 ;
        RECT 460.400 102.200 461.200 106.000 ;
        RECT 462.000 102.200 462.800 106.200 ;
        RECT 463.600 104.800 464.400 106.400 ;
        RECT 465.400 104.400 466.000 107.600 ;
        RECT 470.000 106.200 470.800 119.800 ;
        RECT 471.600 111.600 472.400 113.200 ;
        RECT 471.600 110.300 472.400 110.400 ;
        RECT 474.800 110.300 475.600 119.800 ;
        RECT 476.400 112.400 477.200 119.800 ;
        RECT 479.600 119.200 483.600 119.800 ;
        RECT 479.600 112.400 480.400 119.200 ;
        RECT 476.400 111.800 480.400 112.400 ;
        RECT 481.200 111.800 482.000 118.600 ;
        RECT 482.800 111.800 483.600 119.200 ;
        RECT 484.400 115.000 485.200 119.000 ;
        RECT 481.200 111.200 481.800 111.800 ;
        RECT 484.400 111.600 485.000 115.000 ;
        RECT 488.600 112.800 489.400 119.800 ;
        RECT 488.600 112.200 490.200 112.800 ;
        RECT 477.200 110.400 478.000 110.800 ;
        RECT 479.800 110.600 481.800 111.200 ;
        RECT 479.800 110.400 480.400 110.600 ;
        RECT 471.600 109.700 475.600 110.300 ;
        RECT 471.600 109.600 472.400 109.700 ;
        RECT 473.200 106.800 474.000 108.400 ;
        RECT 470.000 105.600 471.800 106.200 ;
        RECT 471.000 104.400 471.800 105.600 ;
        RECT 465.200 102.200 466.000 104.400 ;
        RECT 470.000 103.600 471.800 104.400 ;
        RECT 471.000 102.200 471.800 103.600 ;
        RECT 474.800 102.200 475.600 109.700 ;
        RECT 476.400 109.800 478.000 110.400 ;
        RECT 476.400 109.600 477.200 109.800 ;
        RECT 479.600 109.600 480.400 110.400 ;
        RECT 482.800 109.600 483.600 111.200 ;
        RECT 484.400 111.000 488.200 111.600 ;
        RECT 478.000 107.600 478.800 109.200 ;
        RECT 479.800 106.200 480.400 109.600 ;
        RECT 481.000 108.800 481.800 109.600 ;
        RECT 484.400 108.800 485.200 110.400 ;
        RECT 486.000 108.800 486.800 110.400 ;
        RECT 487.600 109.000 488.200 111.000 ;
        RECT 481.200 108.400 481.800 108.800 ;
        RECT 481.200 107.600 482.000 108.400 ;
        RECT 487.600 108.200 489.000 109.000 ;
        RECT 489.600 108.400 490.200 112.200 ;
        RECT 490.800 109.600 491.600 111.200 ;
        RECT 487.600 107.800 488.600 108.200 ;
        RECT 484.400 107.200 488.600 107.800 ;
        RECT 489.600 107.600 491.600 108.400 ;
        RECT 492.400 108.300 493.200 108.400 ;
        RECT 494.000 108.300 494.800 108.400 ;
        RECT 492.400 107.700 494.800 108.300 ;
        RECT 492.400 107.600 493.200 107.700 ;
        RECT 479.400 102.200 481.000 106.200 ;
        RECT 484.400 105.000 485.000 107.200 ;
        RECT 489.600 107.000 490.200 107.600 ;
        RECT 489.400 106.600 490.200 107.000 ;
        RECT 494.000 106.800 494.800 107.700 ;
        RECT 488.600 106.000 490.200 106.600 ;
        RECT 495.600 106.200 496.400 119.800 ;
        RECT 497.200 111.600 498.000 113.200 ;
        RECT 501.400 112.400 502.200 119.800 ;
        RECT 502.800 113.600 503.600 114.400 ;
        RECT 503.000 112.400 503.600 113.600 ;
        RECT 501.400 111.800 502.400 112.400 ;
        RECT 503.000 111.800 504.400 112.400 ;
        RECT 500.400 108.800 501.200 110.400 ;
        RECT 501.800 108.400 502.400 111.800 ;
        RECT 503.600 111.600 504.400 111.800 ;
        RECT 505.200 111.600 506.000 113.200 ;
        RECT 503.700 110.300 504.300 111.600 ;
        RECT 506.800 110.300 507.600 119.800 ;
        RECT 510.800 113.600 511.600 114.400 ;
        RECT 510.800 112.400 511.400 113.600 ;
        RECT 512.200 112.400 513.000 119.800 ;
        RECT 510.000 111.800 511.400 112.400 ;
        RECT 512.000 111.800 513.000 112.400 ;
        RECT 518.000 112.000 518.800 119.800 ;
        RECT 521.200 115.200 522.000 119.800 ;
        RECT 510.000 111.600 510.800 111.800 ;
        RECT 503.700 109.700 507.600 110.300 ;
        RECT 498.800 108.200 499.600 108.400 ;
        RECT 498.800 107.600 500.400 108.200 ;
        RECT 501.800 107.600 504.400 108.400 ;
        RECT 499.600 107.200 500.400 107.600 ;
        RECT 499.000 106.200 502.600 106.600 ;
        RECT 503.600 106.200 504.200 107.600 ;
        RECT 506.800 106.200 507.600 109.700 ;
        RECT 512.000 108.400 512.600 111.800 ;
        RECT 517.800 111.200 518.800 112.000 ;
        RECT 519.400 114.600 522.000 115.200 ;
        RECT 519.400 113.000 520.000 114.600 ;
        RECT 524.400 114.400 525.200 119.800 ;
        RECT 527.600 117.000 528.400 119.800 ;
        RECT 529.200 117.000 530.000 119.800 ;
        RECT 530.800 117.000 531.600 119.800 ;
        RECT 525.800 114.400 530.000 115.200 ;
        RECT 522.600 113.600 525.200 114.400 ;
        RECT 532.400 113.600 533.200 119.800 ;
        RECT 535.600 115.000 536.400 119.800 ;
        RECT 538.800 115.000 539.600 119.800 ;
        RECT 540.400 117.000 541.200 119.800 ;
        RECT 542.000 117.000 542.800 119.800 ;
        RECT 545.200 115.200 546.000 119.800 ;
        RECT 548.400 116.400 549.200 119.800 ;
        RECT 548.400 115.800 549.400 116.400 ;
        RECT 548.800 115.200 549.400 115.800 ;
        RECT 544.000 114.400 548.200 115.200 ;
        RECT 548.800 114.600 550.800 115.200 ;
        RECT 535.600 113.600 538.200 114.400 ;
        RECT 538.800 113.800 544.600 114.400 ;
        RECT 547.600 114.000 548.200 114.400 ;
        RECT 527.600 113.000 528.400 113.200 ;
        RECT 519.400 112.400 528.400 113.000 ;
        RECT 530.800 113.000 531.600 113.200 ;
        RECT 538.800 113.000 539.400 113.800 ;
        RECT 545.200 113.200 546.600 113.800 ;
        RECT 547.600 113.200 549.200 114.000 ;
        RECT 530.800 112.400 539.400 113.000 ;
        RECT 540.400 113.000 546.600 113.200 ;
        RECT 540.400 112.600 545.800 113.000 ;
        RECT 540.400 112.400 541.200 112.600 ;
        RECT 513.200 108.800 514.000 110.400 ;
        RECT 508.400 106.800 509.200 108.400 ;
        RECT 510.000 107.600 512.600 108.400 ;
        RECT 514.800 108.200 515.600 108.400 ;
        RECT 514.000 107.600 515.600 108.200 ;
        RECT 510.200 106.200 510.800 107.600 ;
        RECT 514.000 107.200 514.800 107.600 ;
        RECT 517.800 106.800 518.600 111.200 ;
        RECT 519.400 110.600 520.000 112.400 ;
        RECT 519.200 110.000 520.000 110.600 ;
        RECT 526.000 110.000 549.400 110.600 ;
        RECT 519.200 108.000 519.800 110.000 ;
        RECT 526.000 109.400 526.800 110.000 ;
        RECT 543.600 109.600 544.400 110.000 ;
        RECT 545.200 109.600 546.000 110.000 ;
        RECT 548.600 109.800 549.400 110.000 ;
        RECT 520.400 108.600 524.200 109.400 ;
        RECT 519.200 107.400 520.400 108.000 ;
        RECT 511.800 106.200 515.400 106.600 ;
        RECT 484.400 103.000 485.200 105.000 ;
        RECT 488.600 103.000 489.400 106.000 ;
        RECT 495.600 105.600 497.400 106.200 ;
        RECT 496.600 104.400 497.400 105.600 ;
        RECT 498.800 106.000 502.800 106.200 ;
        RECT 496.600 103.600 498.000 104.400 ;
        RECT 496.600 102.200 497.400 103.600 ;
        RECT 498.800 102.200 499.600 106.000 ;
        RECT 502.000 102.200 502.800 106.000 ;
        RECT 503.600 102.200 504.400 106.200 ;
        RECT 505.800 105.600 507.600 106.200 ;
        RECT 505.800 102.200 506.600 105.600 ;
        RECT 510.000 102.200 510.800 106.200 ;
        RECT 511.600 106.000 515.600 106.200 ;
        RECT 517.800 106.000 518.800 106.800 ;
        RECT 511.600 102.200 512.400 106.000 ;
        RECT 514.800 102.200 515.600 106.000 ;
        RECT 518.000 102.200 518.800 106.000 ;
        RECT 519.600 102.200 520.400 107.400 ;
        RECT 523.400 107.400 524.200 108.600 ;
        RECT 523.400 106.800 525.200 107.400 ;
        RECT 524.400 106.200 525.200 106.800 ;
        RECT 529.200 106.400 530.000 109.200 ;
        RECT 532.400 108.600 535.600 109.400 ;
        RECT 539.400 108.600 541.400 109.400 ;
        RECT 550.000 109.000 550.800 114.600 ;
        RECT 532.000 107.800 532.800 108.000 ;
        RECT 532.000 107.200 536.400 107.800 ;
        RECT 535.600 107.000 536.400 107.200 ;
        RECT 537.200 106.800 538.000 108.400 ;
        RECT 524.400 105.400 526.800 106.200 ;
        RECT 529.200 105.600 530.200 106.400 ;
        RECT 533.200 105.600 534.800 106.400 ;
        RECT 535.600 106.200 536.400 106.400 ;
        RECT 539.400 106.200 540.200 108.600 ;
        RECT 542.000 108.200 550.800 109.000 ;
        RECT 545.400 106.800 548.400 107.600 ;
        RECT 545.400 106.200 546.200 106.800 ;
        RECT 535.600 105.600 540.200 106.200 ;
        RECT 526.000 102.200 526.800 105.400 ;
        RECT 543.600 105.400 546.200 106.200 ;
        RECT 527.600 102.200 528.400 105.000 ;
        RECT 529.200 102.200 530.000 105.000 ;
        RECT 530.800 102.200 531.600 105.000 ;
        RECT 532.400 102.200 533.200 105.000 ;
        RECT 535.600 102.200 536.400 105.000 ;
        RECT 538.800 102.200 539.600 105.000 ;
        RECT 540.400 102.200 541.200 105.000 ;
        RECT 542.000 102.200 542.800 105.000 ;
        RECT 543.600 102.200 544.400 105.400 ;
        RECT 550.000 102.200 550.800 108.200 ;
        RECT 3.800 96.400 4.600 99.800 ;
        RECT 2.800 95.800 4.600 96.400 ;
        RECT 7.600 97.800 8.400 99.800 ;
        RECT 12.000 98.300 12.800 99.800 ;
        RECT 14.000 98.300 14.800 98.400 ;
        RECT 1.200 93.600 2.000 95.200 ;
        RECT 2.800 92.300 3.600 95.800 ;
        RECT 7.600 94.400 8.200 97.800 ;
        RECT 12.000 97.700 14.800 98.300 ;
        RECT 9.200 95.600 10.000 97.200 ;
        RECT 7.600 93.600 8.400 94.400 ;
        RECT 12.000 94.200 12.800 97.700 ;
        RECT 14.000 97.600 14.800 97.700 ;
        RECT 18.400 94.200 19.200 99.800 ;
        RECT 23.600 96.000 24.400 99.800 ;
        RECT 26.800 96.000 27.600 99.800 ;
        RECT 23.600 95.800 27.600 96.000 ;
        RECT 28.400 95.800 29.200 99.800 ;
        RECT 32.600 96.400 33.400 99.800 ;
        RECT 37.400 98.400 38.200 99.800 ;
        RECT 37.400 97.600 38.800 98.400 ;
        RECT 37.400 96.400 38.200 97.600 ;
        RECT 31.600 95.800 33.400 96.400 ;
        RECT 36.400 95.800 38.200 96.400 ;
        RECT 39.600 96.000 40.400 99.800 ;
        RECT 42.800 96.000 43.600 99.800 ;
        RECT 39.600 95.800 43.600 96.000 ;
        RECT 44.400 95.800 45.200 99.800 ;
        RECT 23.800 95.400 27.400 95.800 ;
        RECT 24.400 94.400 25.200 94.800 ;
        RECT 28.400 94.400 29.000 95.800 ;
        RECT 11.000 93.800 12.800 94.200 ;
        RECT 17.400 93.800 19.200 94.200 ;
        RECT 23.600 93.800 25.200 94.400 ;
        RECT 11.000 93.600 12.600 93.800 ;
        RECT 17.400 93.600 19.000 93.800 ;
        RECT 23.600 93.600 24.400 93.800 ;
        RECT 26.600 93.600 29.200 94.400 ;
        RECT 30.000 93.600 30.800 95.200 ;
        RECT 31.600 94.300 32.400 95.800 ;
        RECT 34.800 94.300 35.600 95.200 ;
        RECT 31.600 93.700 35.600 94.300 ;
        RECT 6.000 92.300 6.800 92.400 ;
        RECT 2.800 91.700 6.800 92.300 ;
        RECT 2.800 82.200 3.600 91.700 ;
        RECT 6.000 90.800 6.800 91.700 ;
        RECT 4.400 88.800 5.200 90.400 ;
        RECT 7.600 90.200 8.200 93.600 ;
        RECT 11.000 90.400 11.600 93.600 ;
        RECT 13.200 91.600 14.800 92.400 ;
        RECT 6.600 89.400 8.400 90.200 ;
        RECT 10.800 89.600 11.600 90.400 ;
        RECT 15.600 89.600 16.400 91.200 ;
        RECT 17.400 90.400 18.000 93.600 ;
        RECT 19.600 91.600 21.200 92.400 ;
        RECT 23.600 92.300 24.400 92.400 ;
        RECT 25.200 92.300 26.000 93.200 ;
        RECT 23.600 91.700 26.000 92.300 ;
        RECT 23.600 91.600 24.400 91.700 ;
        RECT 25.200 91.600 26.000 91.700 ;
        RECT 26.600 92.300 27.200 93.600 ;
        RECT 30.000 92.300 30.800 92.400 ;
        RECT 26.600 91.700 30.800 92.300 ;
        RECT 17.200 89.600 18.000 90.400 ;
        RECT 22.000 89.600 22.800 91.200 ;
        RECT 26.600 90.200 27.200 91.700 ;
        RECT 30.000 91.600 30.800 91.700 ;
        RECT 28.400 90.200 29.200 90.400 ;
        RECT 26.200 89.600 27.200 90.200 ;
        RECT 27.800 89.600 29.200 90.200 ;
        RECT 6.600 84.400 7.400 89.400 ;
        RECT 11.000 87.000 11.600 89.600 ;
        RECT 12.400 87.600 13.200 89.200 ;
        RECT 17.400 87.000 18.000 89.600 ;
        RECT 18.800 87.600 19.600 89.200 ;
        RECT 11.000 86.400 14.600 87.000 ;
        RECT 11.000 86.200 11.600 86.400 ;
        RECT 6.600 83.600 8.400 84.400 ;
        RECT 6.600 82.200 7.400 83.600 ;
        RECT 10.800 82.200 11.600 86.200 ;
        RECT 14.000 86.200 14.600 86.400 ;
        RECT 17.400 86.400 21.000 87.000 ;
        RECT 17.400 86.200 18.000 86.400 ;
        RECT 14.000 82.200 14.800 86.200 ;
        RECT 17.200 82.200 18.000 86.200 ;
        RECT 20.400 86.200 21.000 86.400 ;
        RECT 20.400 82.200 21.200 86.200 ;
        RECT 26.200 82.200 27.000 89.600 ;
        RECT 27.800 88.400 28.400 89.600 ;
        RECT 27.600 87.600 28.400 88.400 ;
        RECT 31.600 82.200 32.400 93.700 ;
        RECT 34.800 93.600 35.600 93.700 ;
        RECT 33.200 88.800 34.000 90.400 ;
        RECT 36.400 82.200 37.200 95.800 ;
        RECT 39.800 95.400 43.400 95.800 ;
        RECT 40.400 94.400 41.200 94.800 ;
        RECT 44.400 94.400 45.000 95.800 ;
        RECT 39.600 93.800 41.200 94.400 ;
        RECT 39.600 93.600 40.400 93.800 ;
        RECT 42.600 93.600 45.200 94.400 ;
        RECT 46.000 93.800 46.800 99.800 ;
        RECT 52.400 96.600 53.200 99.800 ;
        RECT 54.000 97.000 54.800 99.800 ;
        RECT 55.600 97.000 56.400 99.800 ;
        RECT 57.200 97.000 58.000 99.800 ;
        RECT 60.400 97.000 61.200 99.800 ;
        RECT 63.600 97.000 64.400 99.800 ;
        RECT 65.200 97.000 66.000 99.800 ;
        RECT 66.800 97.000 67.600 99.800 ;
        RECT 68.400 97.000 69.200 99.800 ;
        RECT 50.600 95.800 53.200 96.600 ;
        RECT 70.000 96.600 70.800 99.800 ;
        RECT 56.600 95.800 61.200 96.400 ;
        RECT 50.600 95.200 51.400 95.800 ;
        RECT 48.400 94.400 51.400 95.200 ;
        RECT 41.200 91.600 42.000 93.200 ;
        RECT 38.000 88.800 38.800 90.400 ;
        RECT 42.600 90.200 43.200 93.600 ;
        RECT 46.000 93.000 54.800 93.800 ;
        RECT 56.600 93.400 57.400 95.800 ;
        RECT 60.400 95.600 61.200 95.800 ;
        RECT 62.000 95.600 63.600 96.400 ;
        RECT 66.600 95.600 67.600 96.400 ;
        RECT 70.000 95.800 72.400 96.600 ;
        RECT 58.800 93.600 59.600 95.200 ;
        RECT 60.400 94.800 61.200 95.000 ;
        RECT 60.400 94.200 64.800 94.800 ;
        RECT 64.000 94.000 64.800 94.200 ;
        RECT 44.400 90.200 45.200 90.400 ;
        RECT 42.200 89.600 43.200 90.200 ;
        RECT 43.800 89.600 45.200 90.200 ;
        RECT 42.200 82.200 43.000 89.600 ;
        RECT 43.800 88.400 44.400 89.600 ;
        RECT 43.600 87.600 44.400 88.400 ;
        RECT 46.000 87.400 46.800 93.000 ;
        RECT 55.400 92.600 57.400 93.400 ;
        RECT 61.200 92.600 64.400 93.400 ;
        RECT 66.800 92.800 67.600 95.600 ;
        RECT 71.600 95.200 72.400 95.800 ;
        RECT 71.600 94.600 73.400 95.200 ;
        RECT 72.600 93.400 73.400 94.600 ;
        RECT 76.400 94.600 77.200 99.800 ;
        RECT 78.000 96.000 78.800 99.800 ;
        RECT 78.000 95.200 79.000 96.000 ;
        RECT 81.200 95.800 82.000 99.800 ;
        RECT 82.800 96.000 83.600 99.800 ;
        RECT 86.000 96.000 86.800 99.800 ;
        RECT 89.200 97.800 90.000 99.800 ;
        RECT 82.800 95.800 86.800 96.000 ;
        RECT 76.400 94.000 77.600 94.600 ;
        RECT 72.600 92.600 76.400 93.400 ;
        RECT 77.000 92.000 77.600 94.000 ;
        RECT 76.800 91.400 77.600 92.000 ;
        RECT 75.400 90.800 76.200 91.000 ;
        RECT 47.600 90.300 48.400 90.400 ;
        RECT 49.200 90.300 76.200 90.800 ;
        RECT 47.600 90.200 76.200 90.300 ;
        RECT 47.600 89.700 50.000 90.200 ;
        RECT 52.600 90.000 53.400 90.200 ;
        RECT 47.600 89.600 48.400 89.700 ;
        RECT 49.200 89.600 50.000 89.700 ;
        RECT 76.800 89.600 77.400 91.400 ;
        RECT 78.200 90.800 79.000 95.200 ;
        RECT 81.400 94.400 82.000 95.800 ;
        RECT 83.000 95.400 86.600 95.800 ;
        RECT 87.600 95.600 88.400 97.200 ;
        RECT 89.400 96.300 90.000 97.800 ;
        RECT 92.600 96.400 93.400 97.200 ;
        RECT 92.400 96.300 93.200 96.400 ;
        RECT 89.300 95.700 93.200 96.300 ;
        RECT 94.000 95.800 94.800 99.800 ;
        RECT 85.200 94.400 86.000 94.800 ;
        RECT 89.400 94.400 90.000 95.700 ;
        RECT 92.400 95.600 93.200 95.700 ;
        RECT 81.200 93.600 83.800 94.400 ;
        RECT 85.200 94.300 86.800 94.400 ;
        RECT 87.600 94.300 88.400 94.400 ;
        RECT 85.200 93.800 88.400 94.300 ;
        RECT 86.000 93.700 88.400 93.800 ;
        RECT 86.000 93.600 86.800 93.700 ;
        RECT 87.600 93.600 88.400 93.700 ;
        RECT 89.200 93.600 90.000 94.400 ;
        RECT 90.800 94.300 91.600 94.400 ;
        RECT 94.200 94.300 94.800 95.800 ;
        RECT 90.800 93.700 94.800 94.300 ;
        RECT 90.800 93.600 91.600 93.700 ;
        RECT 55.600 89.400 56.400 89.600 ;
        RECT 51.000 89.000 56.400 89.400 ;
        RECT 50.200 88.800 56.400 89.000 ;
        RECT 57.400 89.000 66.000 89.600 ;
        RECT 47.600 88.000 49.200 88.800 ;
        RECT 50.200 88.200 51.600 88.800 ;
        RECT 57.400 88.200 58.000 89.000 ;
        RECT 65.200 88.800 66.000 89.000 ;
        RECT 68.400 89.000 77.400 89.600 ;
        RECT 68.400 88.800 69.200 89.000 ;
        RECT 48.600 87.600 49.200 88.000 ;
        RECT 52.200 87.600 58.000 88.200 ;
        RECT 58.600 87.600 61.200 88.400 ;
        RECT 46.000 86.800 48.000 87.400 ;
        RECT 48.600 86.800 52.800 87.600 ;
        RECT 47.400 86.200 48.000 86.800 ;
        RECT 47.400 85.600 48.400 86.200 ;
        RECT 47.600 82.200 48.400 85.600 ;
        RECT 50.800 82.200 51.600 86.800 ;
        RECT 54.000 82.200 54.800 85.000 ;
        RECT 55.600 82.200 56.400 85.000 ;
        RECT 57.200 82.200 58.000 87.000 ;
        RECT 60.400 82.200 61.200 87.000 ;
        RECT 63.600 82.200 64.400 88.400 ;
        RECT 71.600 87.600 74.200 88.400 ;
        RECT 66.800 86.800 71.000 87.600 ;
        RECT 65.200 82.200 66.000 85.000 ;
        RECT 66.800 82.200 67.600 85.000 ;
        RECT 68.400 82.200 69.200 85.000 ;
        RECT 71.600 82.200 72.400 87.600 ;
        RECT 76.800 87.400 77.400 89.000 ;
        RECT 74.800 86.800 77.400 87.400 ;
        RECT 78.000 90.000 79.000 90.800 ;
        RECT 81.200 90.200 82.000 90.400 ;
        RECT 83.200 90.200 83.800 93.600 ;
        RECT 84.400 91.600 85.200 93.200 ;
        RECT 89.400 90.200 90.000 93.600 ;
        RECT 90.800 90.800 91.600 92.400 ;
        RECT 92.400 92.200 93.200 92.400 ;
        RECT 94.200 92.200 94.800 93.700 ;
        RECT 95.600 92.800 96.400 94.400 ;
        RECT 98.800 93.800 99.600 99.800 ;
        RECT 105.200 96.600 106.000 99.800 ;
        RECT 106.800 97.000 107.600 99.800 ;
        RECT 108.400 97.000 109.200 99.800 ;
        RECT 110.000 97.000 110.800 99.800 ;
        RECT 113.200 97.000 114.000 99.800 ;
        RECT 116.400 97.000 117.200 99.800 ;
        RECT 118.000 97.000 118.800 99.800 ;
        RECT 119.600 97.000 120.400 99.800 ;
        RECT 121.200 97.000 122.000 99.800 ;
        RECT 103.400 95.800 106.000 96.600 ;
        RECT 122.800 96.600 123.600 99.800 ;
        RECT 109.400 95.800 114.000 96.400 ;
        RECT 103.400 95.200 104.200 95.800 ;
        RECT 101.200 94.400 104.200 95.200 ;
        RECT 98.800 93.000 107.600 93.800 ;
        RECT 109.400 93.400 110.200 95.800 ;
        RECT 113.200 95.600 114.000 95.800 ;
        RECT 114.800 95.600 116.400 96.400 ;
        RECT 119.400 95.600 120.400 96.400 ;
        RECT 122.800 95.800 125.200 96.600 ;
        RECT 111.600 93.600 112.400 95.200 ;
        RECT 113.200 94.800 114.000 95.000 ;
        RECT 113.200 94.200 117.600 94.800 ;
        RECT 116.800 94.000 117.600 94.200 ;
        RECT 97.200 92.200 98.000 92.400 ;
        RECT 92.400 91.600 94.800 92.200 ;
        RECT 96.400 91.600 98.000 92.200 ;
        RECT 92.600 90.200 93.200 91.600 ;
        RECT 96.400 91.200 97.200 91.600 ;
        RECT 78.000 88.300 78.800 90.000 ;
        RECT 81.200 89.600 82.600 90.200 ;
        RECT 83.200 89.600 84.200 90.200 ;
        RECT 82.000 88.400 82.600 89.600 ;
        RECT 79.600 88.300 80.400 88.400 ;
        RECT 78.000 87.700 80.400 88.300 ;
        RECT 74.800 82.200 75.600 86.800 ;
        RECT 78.000 82.200 78.800 87.700 ;
        RECT 79.600 87.600 80.400 87.700 ;
        RECT 82.000 87.600 82.800 88.400 ;
        RECT 83.400 82.200 84.200 89.600 ;
        RECT 89.200 89.400 91.000 90.200 ;
        RECT 90.200 82.200 91.000 89.400 ;
        RECT 92.400 82.200 93.200 90.200 ;
        RECT 94.000 89.600 98.000 90.200 ;
        RECT 94.000 82.200 94.800 89.600 ;
        RECT 97.200 82.200 98.000 89.600 ;
        RECT 98.800 87.400 99.600 93.000 ;
        RECT 108.200 92.600 110.200 93.400 ;
        RECT 114.000 92.600 117.200 93.400 ;
        RECT 119.600 92.800 120.400 95.600 ;
        RECT 124.400 95.200 125.200 95.800 ;
        RECT 124.400 94.600 126.200 95.200 ;
        RECT 125.400 93.400 126.200 94.600 ;
        RECT 129.200 94.600 130.000 99.800 ;
        RECT 130.800 96.300 131.600 99.800 ;
        RECT 137.200 96.300 138.000 96.400 ;
        RECT 130.800 95.700 138.000 96.300 ;
        RECT 130.800 95.200 131.800 95.700 ;
        RECT 137.200 95.600 138.000 95.700 ;
        RECT 129.200 94.000 130.400 94.600 ;
        RECT 125.400 92.600 129.200 93.400 ;
        RECT 100.200 92.000 101.000 92.200 ;
        RECT 103.600 92.000 104.400 92.400 ;
        RECT 105.200 92.000 106.000 92.400 ;
        RECT 122.800 92.000 123.600 92.600 ;
        RECT 129.800 92.000 130.400 94.000 ;
        RECT 100.200 91.400 123.600 92.000 ;
        RECT 129.600 91.400 130.400 92.000 ;
        RECT 129.600 89.600 130.200 91.400 ;
        RECT 131.000 90.800 131.800 95.200 ;
        RECT 108.400 89.400 109.200 89.600 ;
        RECT 103.800 89.000 109.200 89.400 ;
        RECT 103.000 88.800 109.200 89.000 ;
        RECT 110.200 89.000 118.800 89.600 ;
        RECT 100.400 88.000 102.000 88.800 ;
        RECT 103.000 88.200 104.400 88.800 ;
        RECT 110.200 88.200 110.800 89.000 ;
        RECT 118.000 88.800 118.800 89.000 ;
        RECT 121.200 89.000 130.200 89.600 ;
        RECT 121.200 88.800 122.000 89.000 ;
        RECT 101.400 87.600 102.000 88.000 ;
        RECT 105.000 87.600 110.800 88.200 ;
        RECT 111.400 87.600 114.000 88.400 ;
        RECT 98.800 86.800 100.800 87.400 ;
        RECT 101.400 86.800 105.600 87.600 ;
        RECT 100.200 86.200 100.800 86.800 ;
        RECT 100.200 85.600 101.200 86.200 ;
        RECT 100.400 82.200 101.200 85.600 ;
        RECT 103.600 82.200 104.400 86.800 ;
        RECT 106.800 82.200 107.600 85.000 ;
        RECT 108.400 82.200 109.200 85.000 ;
        RECT 110.000 82.200 110.800 87.000 ;
        RECT 113.200 82.200 114.000 87.000 ;
        RECT 116.400 82.200 117.200 88.400 ;
        RECT 124.400 87.600 127.000 88.400 ;
        RECT 119.600 86.800 123.800 87.600 ;
        RECT 118.000 82.200 118.800 85.000 ;
        RECT 119.600 82.200 120.400 85.000 ;
        RECT 121.200 82.200 122.000 85.000 ;
        RECT 124.400 82.200 125.200 87.600 ;
        RECT 129.600 87.400 130.200 89.000 ;
        RECT 127.600 86.800 130.200 87.400 ;
        RECT 130.800 90.000 131.800 90.800 ;
        RECT 127.600 82.200 128.400 86.800 ;
        RECT 130.800 82.200 131.600 90.000 ;
        RECT 140.400 82.200 141.200 99.800 ;
        RECT 145.200 97.800 146.000 99.800 ;
        RECT 142.000 95.600 142.800 97.200 ;
        RECT 143.600 95.600 144.400 97.200 ;
        RECT 145.400 95.600 146.000 97.800 ;
        RECT 148.400 95.800 149.200 99.800 ;
        RECT 150.000 95.800 150.800 99.800 ;
        RECT 151.600 96.000 152.400 99.800 ;
        RECT 154.800 96.000 155.600 99.800 ;
        RECT 151.600 95.800 155.600 96.000 ;
        RECT 145.400 95.000 147.800 95.600 ;
        RECT 145.200 93.600 146.200 94.400 ;
        RECT 145.600 92.800 146.400 93.600 ;
        RECT 147.200 92.000 147.800 95.000 ;
        RECT 148.600 92.400 149.200 95.800 ;
        RECT 150.200 94.400 150.800 95.800 ;
        RECT 151.800 95.400 155.400 95.800 ;
        RECT 156.400 95.000 157.200 99.800 ;
        RECT 160.800 98.400 161.600 99.800 ;
        RECT 159.600 97.800 161.600 98.400 ;
        RECT 165.200 97.800 166.000 99.800 ;
        RECT 169.400 98.400 170.600 99.800 ;
        RECT 169.200 97.800 170.600 98.400 ;
        RECT 159.600 97.000 160.400 97.800 ;
        RECT 165.200 97.200 165.800 97.800 ;
        RECT 161.200 96.400 162.000 97.200 ;
        RECT 163.000 96.600 165.800 97.200 ;
        RECT 169.200 97.000 170.000 97.800 ;
        RECT 163.000 96.400 163.800 96.600 ;
        RECT 154.000 94.400 154.800 94.800 ;
        RECT 150.000 93.600 152.600 94.400 ;
        RECT 154.000 93.800 155.600 94.400 ;
        RECT 154.800 93.600 155.600 93.800 ;
        RECT 157.200 94.200 158.800 94.400 ;
        RECT 161.400 94.200 162.000 96.400 ;
        RECT 171.000 95.400 171.800 95.600 ;
        RECT 174.000 95.400 174.800 99.800 ;
        RECT 171.000 94.800 174.800 95.400 ;
        RECT 164.400 94.200 165.200 94.400 ;
        RECT 167.000 94.200 167.800 94.400 ;
        RECT 157.200 93.600 168.200 94.200 ;
        RECT 147.000 91.400 147.800 92.000 ;
        RECT 148.400 92.300 149.200 92.400 ;
        RECT 150.000 92.300 150.800 92.400 ;
        RECT 148.400 91.700 150.800 92.300 ;
        RECT 148.400 91.600 149.200 91.700 ;
        RECT 150.000 91.600 150.800 91.700 ;
        RECT 143.600 91.200 147.800 91.400 ;
        RECT 143.600 90.800 147.600 91.200 ;
        RECT 143.600 82.200 144.400 90.800 ;
        RECT 148.600 90.200 149.200 91.600 ;
        RECT 152.000 90.400 152.600 93.600 ;
        RECT 160.200 93.400 161.000 93.600 ;
        RECT 153.200 91.600 154.000 93.200 ;
        RECT 158.600 92.400 159.400 92.600 ;
        RECT 161.200 92.400 162.000 92.600 ;
        RECT 158.600 91.800 163.600 92.400 ;
        RECT 162.800 91.600 163.600 91.800 ;
        RECT 156.400 91.000 162.000 91.200 ;
        RECT 156.400 90.800 162.200 91.000 ;
        RECT 156.400 90.600 166.200 90.800 ;
        RECT 147.800 89.600 149.200 90.200 ;
        RECT 150.000 90.200 150.800 90.400 ;
        RECT 150.000 89.600 151.400 90.200 ;
        RECT 152.000 89.600 154.000 90.400 ;
        RECT 147.800 82.200 148.600 89.600 ;
        RECT 150.800 88.400 151.400 89.600 ;
        RECT 150.800 87.600 151.600 88.400 ;
        RECT 152.200 82.200 153.000 89.600 ;
        RECT 156.400 82.200 157.200 90.600 ;
        RECT 161.400 90.200 166.200 90.600 ;
        RECT 159.600 89.000 165.000 89.600 ;
        RECT 159.600 88.800 160.400 89.000 ;
        RECT 164.200 88.800 165.000 89.000 ;
        RECT 165.600 89.000 166.200 90.200 ;
        RECT 167.600 90.400 168.200 93.600 ;
        RECT 169.200 92.800 170.000 93.000 ;
        RECT 169.200 92.200 173.000 92.800 ;
        RECT 172.200 92.000 173.000 92.200 ;
        RECT 170.600 91.400 171.400 91.600 ;
        RECT 174.000 91.400 174.800 94.800 ;
        RECT 175.600 95.200 176.400 99.800 ;
        RECT 175.600 94.600 177.800 95.200 ;
        RECT 170.600 90.800 174.800 91.400 ;
        RECT 167.600 89.800 170.000 90.400 ;
        RECT 167.000 89.000 167.800 89.200 ;
        RECT 165.600 88.400 167.800 89.000 ;
        RECT 169.400 88.800 170.000 89.800 ;
        RECT 169.400 88.000 170.800 88.800 ;
        RECT 163.000 87.400 163.800 87.600 ;
        RECT 165.800 87.400 166.600 87.600 ;
        RECT 159.600 86.200 160.400 87.000 ;
        RECT 163.000 86.800 166.600 87.400 ;
        RECT 165.200 86.200 165.800 86.800 ;
        RECT 169.200 86.200 170.000 87.000 ;
        RECT 159.600 85.600 161.600 86.200 ;
        RECT 160.800 82.200 161.600 85.600 ;
        RECT 165.200 82.200 166.000 86.200 ;
        RECT 169.400 82.200 170.600 86.200 ;
        RECT 174.000 82.200 174.800 90.800 ;
        RECT 177.200 91.600 177.800 94.600 ;
        RECT 178.800 92.400 179.600 99.800 ;
        RECT 180.400 95.200 181.200 99.800 ;
        RECT 180.400 94.600 182.600 95.200 ;
        RECT 177.200 90.800 178.400 91.600 ;
        RECT 177.200 90.200 177.800 90.800 ;
        RECT 179.000 90.200 179.600 92.400 ;
        RECT 182.000 91.600 182.600 94.600 ;
        RECT 183.600 92.400 184.400 99.800 ;
        RECT 185.200 95.600 186.000 97.200 ;
        RECT 182.000 90.800 183.200 91.600 ;
        RECT 182.000 90.200 182.600 90.800 ;
        RECT 183.800 90.200 184.400 92.400 ;
        RECT 175.600 89.600 177.800 90.200 ;
        RECT 175.600 82.200 176.400 89.600 ;
        RECT 178.800 82.200 179.600 90.200 ;
        RECT 180.400 89.600 182.600 90.200 ;
        RECT 180.400 82.200 181.200 89.600 ;
        RECT 183.600 82.200 184.400 90.200 ;
        RECT 186.800 94.300 187.600 99.800 ;
        RECT 191.600 95.800 192.400 99.800 ;
        RECT 193.000 96.400 193.800 97.200 ;
        RECT 197.400 96.400 198.200 99.800 ;
        RECT 190.000 94.300 190.800 94.400 ;
        RECT 186.800 93.700 190.800 94.300 ;
        RECT 186.800 82.200 187.600 93.700 ;
        RECT 190.000 92.800 190.800 93.700 ;
        RECT 188.400 92.200 189.200 92.400 ;
        RECT 191.600 92.200 192.200 95.800 ;
        RECT 193.200 95.600 194.000 96.400 ;
        RECT 196.400 95.800 198.200 96.400 ;
        RECT 200.200 96.400 201.000 99.800 ;
        RECT 200.200 95.800 202.000 96.400 ;
        RECT 204.400 95.800 205.200 99.800 ;
        RECT 206.000 96.000 206.800 99.800 ;
        RECT 209.200 96.000 210.000 99.800 ;
        RECT 206.000 95.800 210.000 96.000 ;
        RECT 193.200 94.300 194.000 94.400 ;
        RECT 194.800 94.300 195.600 95.200 ;
        RECT 193.200 93.700 195.600 94.300 ;
        RECT 193.200 93.600 194.000 93.700 ;
        RECT 194.800 93.600 195.600 93.700 ;
        RECT 193.200 92.200 194.000 92.400 ;
        RECT 188.400 91.600 190.000 92.200 ;
        RECT 191.600 91.600 194.000 92.200 ;
        RECT 189.200 91.200 190.000 91.600 ;
        RECT 193.200 90.200 193.800 91.600 ;
        RECT 188.400 89.600 192.400 90.200 ;
        RECT 188.400 82.200 189.200 89.600 ;
        RECT 191.600 82.200 192.400 89.600 ;
        RECT 193.200 82.200 194.000 90.200 ;
        RECT 196.400 82.200 197.200 95.800 ;
        RECT 201.200 92.300 202.000 95.800 ;
        RECT 202.800 94.300 203.600 95.200 ;
        RECT 204.600 94.400 205.200 95.800 ;
        RECT 206.200 95.400 209.800 95.800 ;
        RECT 208.400 94.400 209.200 94.800 ;
        RECT 204.400 94.300 207.000 94.400 ;
        RECT 202.800 93.700 207.000 94.300 ;
        RECT 208.400 93.800 210.000 94.400 ;
        RECT 202.800 93.600 203.600 93.700 ;
        RECT 204.400 93.600 207.000 93.700 ;
        RECT 209.200 93.600 210.000 93.800 ;
        RECT 210.800 94.300 211.600 99.800 ;
        RECT 212.400 95.600 213.200 97.200 ;
        RECT 216.600 96.400 217.400 99.800 ;
        RECT 220.400 97.800 221.200 99.800 ;
        RECT 215.600 95.800 217.400 96.400 ;
        RECT 214.000 94.300 214.800 95.200 ;
        RECT 210.800 93.700 214.800 94.300 ;
        RECT 198.100 91.700 202.000 92.300 ;
        RECT 198.100 90.400 198.700 91.700 ;
        RECT 198.000 88.800 198.800 90.400 ;
        RECT 199.600 88.800 200.400 90.400 ;
        RECT 201.200 82.200 202.000 91.700 ;
        RECT 204.400 90.200 205.200 90.400 ;
        RECT 206.400 90.200 207.000 93.600 ;
        RECT 207.600 91.600 208.400 93.200 ;
        RECT 204.400 89.600 205.800 90.200 ;
        RECT 206.400 89.600 207.400 90.200 ;
        RECT 205.200 88.400 205.800 89.600 ;
        RECT 205.200 87.600 206.000 88.400 ;
        RECT 206.600 82.200 207.400 89.600 ;
        RECT 210.800 82.200 211.600 93.700 ;
        RECT 214.000 93.600 214.800 93.700 ;
        RECT 212.400 90.300 213.200 90.400 ;
        RECT 215.600 90.300 216.400 95.800 ;
        RECT 218.800 95.600 219.600 97.200 ;
        RECT 220.600 94.400 221.200 97.800 ;
        RECT 226.200 96.400 227.000 99.800 ;
        RECT 225.200 95.600 227.600 96.400 ;
        RECT 228.400 95.600 229.200 97.200 ;
        RECT 220.400 93.600 221.200 94.400 ;
        RECT 223.600 93.600 224.400 95.200 ;
        RECT 220.600 92.300 221.200 93.600 ;
        RECT 217.300 91.700 221.200 92.300 ;
        RECT 217.300 90.400 217.900 91.700 ;
        RECT 212.400 89.700 216.400 90.300 ;
        RECT 212.400 89.600 213.200 89.700 ;
        RECT 215.600 82.200 216.400 89.700 ;
        RECT 217.200 88.800 218.000 90.400 ;
        RECT 220.600 90.200 221.200 91.700 ;
        RECT 222.000 90.800 222.800 92.400 ;
        RECT 220.400 89.400 222.200 90.200 ;
        RECT 221.400 88.300 222.200 89.400 ;
        RECT 223.600 88.300 224.400 88.400 ;
        RECT 221.400 87.700 224.400 88.300 ;
        RECT 221.400 82.200 222.200 87.700 ;
        RECT 223.600 87.600 224.400 87.700 ;
        RECT 225.200 82.200 226.000 95.600 ;
        RECT 230.000 94.300 230.800 99.800 ;
        RECT 231.800 96.400 232.600 97.200 ;
        RECT 231.600 95.600 232.400 96.400 ;
        RECT 233.200 95.800 234.000 99.800 ;
        RECT 238.000 96.000 238.800 99.800 ;
        RECT 241.200 96.000 242.000 99.800 ;
        RECT 238.000 95.800 242.000 96.000 ;
        RECT 242.800 95.800 243.600 99.800 ;
        RECT 247.600 98.400 248.400 99.800 ;
        RECT 247.600 97.800 248.600 98.400 ;
        RECT 248.000 97.600 248.600 97.800 ;
        RECT 250.800 97.800 251.600 99.800 ;
        RECT 250.800 97.600 252.000 97.800 ;
        RECT 248.000 97.000 252.000 97.600 ;
        RECT 246.000 96.300 247.800 96.400 ;
        RECT 249.200 96.300 250.000 96.400 ;
        RECT 231.600 94.300 232.400 94.400 ;
        RECT 230.000 93.700 232.400 94.300 ;
        RECT 226.800 88.800 227.600 90.400 ;
        RECT 230.000 82.200 230.800 93.700 ;
        RECT 231.600 93.600 232.400 93.700 ;
        RECT 231.600 92.200 232.400 92.400 ;
        RECT 233.400 92.200 234.000 95.800 ;
        RECT 238.200 95.400 241.800 95.800 ;
        RECT 238.800 94.400 239.600 94.800 ;
        RECT 242.800 94.400 243.400 95.800 ;
        RECT 246.000 95.700 250.000 96.300 ;
        RECT 246.000 95.600 247.800 95.700 ;
        RECT 249.200 95.600 250.000 95.700 ;
        RECT 234.800 92.800 235.600 94.400 ;
        RECT 238.000 93.800 239.600 94.400 ;
        RECT 238.000 93.600 238.800 93.800 ;
        RECT 241.000 93.600 243.600 94.400 ;
        RECT 244.400 94.300 245.200 94.400 ;
        RECT 247.600 94.300 249.200 94.400 ;
        RECT 244.400 93.700 249.200 94.300 ;
        RECT 244.400 93.600 245.200 93.700 ;
        RECT 247.600 93.600 249.200 93.700 ;
        RECT 236.400 92.300 237.200 92.400 ;
        RECT 239.600 92.300 240.400 93.200 ;
        RECT 236.400 92.200 240.400 92.300 ;
        RECT 231.600 91.600 234.000 92.200 ;
        RECT 235.600 91.700 240.400 92.200 ;
        RECT 235.600 91.600 237.200 91.700 ;
        RECT 239.600 91.600 240.400 91.700 ;
        RECT 241.000 92.300 241.600 93.600 ;
        RECT 246.000 92.300 246.800 92.400 ;
        RECT 241.000 91.700 246.800 92.300 ;
        RECT 231.800 90.200 232.400 91.600 ;
        RECT 235.600 91.200 236.400 91.600 ;
        RECT 241.000 90.200 241.600 91.700 ;
        RECT 246.000 91.600 246.800 91.700 ;
        RECT 247.600 92.300 248.400 92.400 ;
        RECT 249.200 92.300 250.800 92.400 ;
        RECT 247.600 91.700 250.800 92.300 ;
        RECT 247.600 91.600 248.400 91.700 ;
        RECT 249.200 91.600 250.800 91.700 ;
        RECT 251.400 90.400 252.000 97.000 ;
        RECT 258.800 97.600 259.600 99.800 ;
        RECT 258.800 94.400 259.400 97.600 ;
        RECT 260.400 96.300 261.200 97.200 ;
        RECT 270.000 96.300 270.800 99.800 ;
        RECT 260.400 95.700 270.800 96.300 ;
        RECT 260.400 95.600 261.200 95.700 ;
        RECT 269.800 95.200 270.800 95.700 ;
        RECT 258.800 93.600 259.600 94.400 ;
        RECT 257.200 90.800 258.000 92.400 ;
        RECT 242.800 90.200 243.600 90.400 ;
        RECT 231.600 82.200 232.400 90.200 ;
        RECT 233.200 89.600 237.200 90.200 ;
        RECT 233.200 82.200 234.000 89.600 ;
        RECT 236.400 82.200 237.200 89.600 ;
        RECT 240.600 89.600 241.600 90.200 ;
        RECT 242.200 89.600 243.600 90.200 ;
        RECT 251.400 89.800 254.800 90.400 ;
        RECT 258.800 90.200 259.400 93.600 ;
        RECT 269.800 90.800 270.600 95.200 ;
        RECT 271.600 94.600 272.400 99.800 ;
        RECT 278.000 96.600 278.800 99.800 ;
        RECT 279.600 97.000 280.400 99.800 ;
        RECT 281.200 97.000 282.000 99.800 ;
        RECT 282.800 97.000 283.600 99.800 ;
        RECT 284.400 97.000 285.200 99.800 ;
        RECT 287.600 97.000 288.400 99.800 ;
        RECT 290.800 97.000 291.600 99.800 ;
        RECT 292.400 97.000 293.200 99.800 ;
        RECT 294.000 97.000 294.800 99.800 ;
        RECT 276.400 95.800 278.800 96.600 ;
        RECT 295.600 96.600 296.400 99.800 ;
        RECT 276.400 95.200 277.200 95.800 ;
        RECT 271.200 94.000 272.400 94.600 ;
        RECT 275.400 94.600 277.200 95.200 ;
        RECT 281.200 95.600 282.200 96.400 ;
        RECT 285.200 95.600 286.800 96.400 ;
        RECT 287.600 95.800 292.200 96.400 ;
        RECT 295.600 95.800 298.200 96.600 ;
        RECT 287.600 95.600 288.400 95.800 ;
        RECT 271.200 92.000 271.800 94.000 ;
        RECT 275.400 93.400 276.200 94.600 ;
        RECT 272.400 92.600 276.200 93.400 ;
        RECT 281.200 92.800 282.000 95.600 ;
        RECT 287.600 94.800 288.400 95.000 ;
        RECT 284.000 94.200 288.400 94.800 ;
        RECT 284.000 94.000 284.800 94.200 ;
        RECT 289.200 93.600 290.000 95.200 ;
        RECT 291.400 93.400 292.200 95.800 ;
        RECT 297.400 95.200 298.200 95.800 ;
        RECT 297.400 94.400 300.400 95.200 ;
        RECT 302.000 93.800 302.800 99.800 ;
        RECT 303.600 95.600 304.400 97.200 ;
        RECT 284.400 92.600 287.600 93.400 ;
        RECT 291.400 92.600 293.400 93.400 ;
        RECT 294.000 93.000 302.800 93.800 ;
        RECT 278.000 92.000 278.800 92.600 ;
        RECT 295.600 92.000 296.400 92.400 ;
        RECT 300.400 92.200 301.200 92.400 ;
        RECT 300.400 92.000 301.400 92.200 ;
        RECT 271.200 91.400 272.000 92.000 ;
        RECT 278.000 91.400 301.400 92.000 ;
        RECT 254.000 89.600 254.800 89.800 ;
        RECT 240.600 82.200 241.400 89.600 ;
        RECT 242.200 88.400 242.800 89.600 ;
        RECT 242.000 87.600 242.800 88.400 ;
        RECT 244.600 88.800 248.200 89.400 ;
        RECT 244.600 88.200 245.200 88.800 ;
        RECT 244.400 82.200 245.200 88.200 ;
        RECT 247.600 88.200 248.200 88.800 ;
        RECT 249.400 89.000 253.000 89.200 ;
        RECT 254.000 89.000 254.600 89.600 ;
        RECT 257.800 89.400 259.600 90.200 ;
        RECT 269.800 90.000 270.800 90.800 ;
        RECT 249.400 88.600 253.200 89.000 ;
        RECT 249.400 88.200 250.000 88.600 ;
        RECT 247.600 82.800 248.400 88.200 ;
        RECT 249.200 83.400 250.000 88.200 ;
        RECT 250.800 82.800 251.600 88.000 ;
        RECT 252.400 83.000 253.200 88.600 ;
        RECT 254.000 83.400 254.800 89.000 ;
        RECT 247.600 82.200 251.600 82.800 ;
        RECT 252.600 82.800 253.200 83.000 ;
        RECT 255.600 83.000 256.400 89.000 ;
        RECT 255.600 82.800 256.200 83.000 ;
        RECT 252.600 82.200 256.200 82.800 ;
        RECT 257.800 82.200 258.600 89.400 ;
        RECT 270.000 82.200 270.800 90.000 ;
        RECT 271.400 89.600 272.000 91.400 ;
        RECT 271.400 89.000 280.400 89.600 ;
        RECT 271.400 87.400 272.000 89.000 ;
        RECT 279.600 88.800 280.400 89.000 ;
        RECT 282.800 89.000 291.400 89.600 ;
        RECT 282.800 88.800 283.600 89.000 ;
        RECT 274.600 87.600 277.200 88.400 ;
        RECT 271.400 86.800 274.000 87.400 ;
        RECT 273.200 82.200 274.000 86.800 ;
        RECT 276.400 82.200 277.200 87.600 ;
        RECT 277.800 86.800 282.000 87.600 ;
        RECT 279.600 82.200 280.400 85.000 ;
        RECT 281.200 82.200 282.000 85.000 ;
        RECT 282.800 82.200 283.600 85.000 ;
        RECT 284.400 82.200 285.200 88.400 ;
        RECT 287.600 87.600 290.200 88.400 ;
        RECT 290.800 88.200 291.400 89.000 ;
        RECT 292.400 89.400 293.200 89.600 ;
        RECT 292.400 89.000 297.800 89.400 ;
        RECT 292.400 88.800 298.600 89.000 ;
        RECT 297.200 88.200 298.600 88.800 ;
        RECT 290.800 87.600 296.600 88.200 ;
        RECT 299.600 88.000 301.200 88.800 ;
        RECT 299.600 87.600 300.200 88.000 ;
        RECT 287.600 82.200 288.400 87.000 ;
        RECT 290.800 82.200 291.600 87.000 ;
        RECT 296.000 86.800 300.200 87.600 ;
        RECT 302.000 87.400 302.800 93.000 ;
        RECT 300.800 86.800 302.800 87.400 ;
        RECT 292.400 82.200 293.200 85.000 ;
        RECT 294.000 82.200 294.800 85.000 ;
        RECT 297.200 82.200 298.000 86.800 ;
        RECT 300.800 86.200 301.400 86.800 ;
        RECT 300.400 85.600 301.400 86.200 ;
        RECT 300.400 82.200 301.200 85.600 ;
        RECT 305.200 82.200 306.000 99.800 ;
        RECT 306.800 96.300 307.600 96.400 ;
        RECT 308.400 96.300 309.200 99.800 ;
        RECT 306.800 95.700 309.200 96.300 ;
        RECT 306.800 95.600 307.600 95.700 ;
        RECT 308.200 95.200 309.200 95.700 ;
        RECT 308.200 90.800 309.000 95.200 ;
        RECT 310.000 94.600 310.800 99.800 ;
        RECT 316.400 96.600 317.200 99.800 ;
        RECT 318.000 97.000 318.800 99.800 ;
        RECT 319.600 97.000 320.400 99.800 ;
        RECT 321.200 97.000 322.000 99.800 ;
        RECT 322.800 97.000 323.600 99.800 ;
        RECT 326.000 97.000 326.800 99.800 ;
        RECT 329.200 97.000 330.000 99.800 ;
        RECT 330.800 97.000 331.600 99.800 ;
        RECT 332.400 97.000 333.200 99.800 ;
        RECT 314.800 95.800 317.200 96.600 ;
        RECT 334.000 96.600 334.800 99.800 ;
        RECT 314.800 95.200 315.600 95.800 ;
        RECT 309.600 94.000 310.800 94.600 ;
        RECT 313.800 94.600 315.600 95.200 ;
        RECT 319.600 95.600 320.600 96.400 ;
        RECT 323.600 95.600 325.200 96.400 ;
        RECT 326.000 95.800 330.600 96.400 ;
        RECT 334.000 95.800 336.600 96.600 ;
        RECT 326.000 95.600 326.800 95.800 ;
        RECT 309.600 92.000 310.200 94.000 ;
        RECT 313.800 93.400 314.600 94.600 ;
        RECT 310.800 92.600 314.600 93.400 ;
        RECT 319.600 92.800 320.400 95.600 ;
        RECT 326.000 94.800 326.800 95.000 ;
        RECT 322.400 94.200 326.800 94.800 ;
        RECT 322.400 94.000 323.200 94.200 ;
        RECT 327.600 93.600 328.400 95.200 ;
        RECT 329.800 93.400 330.600 95.800 ;
        RECT 335.800 95.200 336.600 95.800 ;
        RECT 335.800 94.400 338.800 95.200 ;
        RECT 340.400 93.800 341.200 99.800 ;
        RECT 342.000 96.000 342.800 99.800 ;
        RECT 345.200 96.000 346.000 99.800 ;
        RECT 342.000 95.800 346.000 96.000 ;
        RECT 346.800 95.800 347.600 99.800 ;
        RECT 348.400 95.800 349.200 99.800 ;
        RECT 350.000 96.000 350.800 99.800 ;
        RECT 353.200 96.000 354.000 99.800 ;
        RECT 350.000 95.800 354.000 96.000 ;
        RECT 342.200 95.400 345.800 95.800 ;
        RECT 342.800 94.400 343.600 94.800 ;
        RECT 346.800 94.400 347.400 95.800 ;
        RECT 348.600 94.400 349.200 95.800 ;
        RECT 350.200 95.400 353.800 95.800 ;
        RECT 352.400 94.400 353.200 94.800 ;
        RECT 322.800 92.600 326.000 93.400 ;
        RECT 329.800 92.600 331.800 93.400 ;
        RECT 332.400 93.000 341.200 93.800 ;
        RECT 342.000 93.800 343.600 94.400 ;
        RECT 342.000 93.600 342.800 93.800 ;
        RECT 345.000 93.600 347.600 94.400 ;
        RECT 348.400 93.600 351.000 94.400 ;
        RECT 352.400 93.800 354.000 94.400 ;
        RECT 353.200 93.600 354.000 93.800 ;
        RECT 354.800 93.800 355.600 99.800 ;
        RECT 361.200 96.600 362.000 99.800 ;
        RECT 362.800 97.000 363.600 99.800 ;
        RECT 364.400 97.000 365.200 99.800 ;
        RECT 366.000 97.000 366.800 99.800 ;
        RECT 369.200 97.000 370.000 99.800 ;
        RECT 372.400 97.000 373.200 99.800 ;
        RECT 374.000 97.000 374.800 99.800 ;
        RECT 375.600 97.000 376.400 99.800 ;
        RECT 377.200 97.000 378.000 99.800 ;
        RECT 359.400 95.800 362.000 96.600 ;
        RECT 378.800 96.600 379.600 99.800 ;
        RECT 365.400 95.800 370.000 96.400 ;
        RECT 359.400 95.200 360.200 95.800 ;
        RECT 357.200 94.400 360.200 95.200 ;
        RECT 309.600 91.400 310.400 92.000 ;
        RECT 308.200 90.000 309.200 90.800 ;
        RECT 308.400 82.200 309.200 90.000 ;
        RECT 309.800 89.600 310.400 91.400 ;
        RECT 311.000 90.800 311.800 91.000 ;
        RECT 311.000 90.200 338.000 90.800 ;
        RECT 333.800 90.000 334.600 90.200 ;
        RECT 337.200 89.600 338.000 90.200 ;
        RECT 309.800 89.000 318.800 89.600 ;
        RECT 309.800 87.400 310.400 89.000 ;
        RECT 318.000 88.800 318.800 89.000 ;
        RECT 321.200 89.000 329.800 89.600 ;
        RECT 321.200 88.800 322.000 89.000 ;
        RECT 313.000 87.600 315.600 88.400 ;
        RECT 309.800 86.800 312.400 87.400 ;
        RECT 311.600 82.200 312.400 86.800 ;
        RECT 314.800 82.200 315.600 87.600 ;
        RECT 316.200 86.800 320.400 87.600 ;
        RECT 318.000 82.200 318.800 85.000 ;
        RECT 319.600 82.200 320.400 85.000 ;
        RECT 321.200 82.200 322.000 85.000 ;
        RECT 322.800 82.200 323.600 88.400 ;
        RECT 326.000 87.600 328.600 88.400 ;
        RECT 329.200 88.200 329.800 89.000 ;
        RECT 330.800 89.400 331.600 89.600 ;
        RECT 330.800 89.000 336.200 89.400 ;
        RECT 330.800 88.800 337.000 89.000 ;
        RECT 335.600 88.200 337.000 88.800 ;
        RECT 329.200 87.600 335.000 88.200 ;
        RECT 338.000 88.000 339.600 88.800 ;
        RECT 338.000 87.600 338.600 88.000 ;
        RECT 326.000 82.200 326.800 87.000 ;
        RECT 329.200 82.200 330.000 87.000 ;
        RECT 334.400 86.800 338.600 87.600 ;
        RECT 340.400 87.400 341.200 93.000 ;
        RECT 343.600 91.600 344.400 93.200 ;
        RECT 345.000 90.200 345.600 93.600 ;
        RECT 350.400 92.300 351.000 93.600 ;
        RECT 346.900 91.700 351.000 92.300 ;
        RECT 346.900 90.400 347.500 91.700 ;
        RECT 346.800 90.200 347.600 90.400 ;
        RECT 339.200 86.800 341.200 87.400 ;
        RECT 344.600 89.600 345.600 90.200 ;
        RECT 346.200 89.600 347.600 90.200 ;
        RECT 348.400 90.200 349.200 90.400 ;
        RECT 350.400 90.200 351.000 91.700 ;
        RECT 354.800 93.000 363.600 93.800 ;
        RECT 365.400 93.400 366.200 95.800 ;
        RECT 369.200 95.600 370.000 95.800 ;
        RECT 370.800 95.600 372.400 96.400 ;
        RECT 375.400 95.600 376.400 96.400 ;
        RECT 378.800 95.800 381.200 96.600 ;
        RECT 367.600 93.600 368.400 95.200 ;
        RECT 369.200 94.800 370.000 95.000 ;
        RECT 369.200 94.200 373.600 94.800 ;
        RECT 372.800 94.000 373.600 94.200 ;
        RECT 348.400 89.600 349.800 90.200 ;
        RECT 350.400 89.600 351.400 90.200 ;
        RECT 330.800 82.200 331.600 85.000 ;
        RECT 332.400 82.200 333.200 85.000 ;
        RECT 335.600 82.200 336.400 86.800 ;
        RECT 339.200 86.200 339.800 86.800 ;
        RECT 338.800 85.600 339.800 86.200 ;
        RECT 338.800 82.200 339.600 85.600 ;
        RECT 344.600 82.200 345.400 89.600 ;
        RECT 346.200 88.400 346.800 89.600 ;
        RECT 346.000 87.600 346.800 88.400 ;
        RECT 349.200 88.400 349.800 89.600 ;
        RECT 349.200 87.600 350.000 88.400 ;
        RECT 350.600 82.200 351.400 89.600 ;
        RECT 354.800 87.400 355.600 93.000 ;
        RECT 364.200 92.600 366.200 93.400 ;
        RECT 370.000 92.600 373.200 93.400 ;
        RECT 375.600 92.800 376.400 95.600 ;
        RECT 380.400 95.200 381.200 95.800 ;
        RECT 380.400 94.600 382.200 95.200 ;
        RECT 381.400 93.400 382.200 94.600 ;
        RECT 385.200 94.600 386.000 99.800 ;
        RECT 386.800 96.000 387.600 99.800 ;
        RECT 390.600 96.400 391.400 99.800 ;
        RECT 395.400 96.400 396.200 99.800 ;
        RECT 402.200 96.400 403.000 99.800 ;
        RECT 407.000 96.400 407.800 99.800 ;
        RECT 386.800 95.200 387.800 96.000 ;
        RECT 390.600 95.800 392.400 96.400 ;
        RECT 395.400 95.800 397.200 96.400 ;
        RECT 385.200 94.000 386.400 94.600 ;
        RECT 381.400 92.600 385.200 93.400 ;
        RECT 356.200 92.000 357.000 92.200 ;
        RECT 361.200 92.000 362.000 92.400 ;
        RECT 367.600 92.000 368.400 92.400 ;
        RECT 378.800 92.000 379.600 92.600 ;
        RECT 385.800 92.000 386.400 94.000 ;
        RECT 356.200 91.400 379.600 92.000 ;
        RECT 385.600 91.400 386.400 92.000 ;
        RECT 387.000 92.300 387.800 95.200 ;
        RECT 390.000 92.300 390.800 92.400 ;
        RECT 387.000 91.700 390.800 92.300 ;
        RECT 385.600 89.600 386.200 91.400 ;
        RECT 387.000 90.800 387.800 91.700 ;
        RECT 390.000 91.600 390.800 91.700 ;
        RECT 364.400 89.400 365.200 89.600 ;
        RECT 359.800 89.000 365.200 89.400 ;
        RECT 359.000 88.800 365.200 89.000 ;
        RECT 366.200 89.000 374.800 89.600 ;
        RECT 356.400 88.000 358.000 88.800 ;
        RECT 359.000 88.200 360.400 88.800 ;
        RECT 366.200 88.200 366.800 89.000 ;
        RECT 374.000 88.800 374.800 89.000 ;
        RECT 377.200 89.000 386.200 89.600 ;
        RECT 377.200 88.800 378.000 89.000 ;
        RECT 357.400 87.600 358.000 88.000 ;
        RECT 361.000 87.600 366.800 88.200 ;
        RECT 367.400 87.600 370.000 88.400 ;
        RECT 354.800 86.800 356.800 87.400 ;
        RECT 357.400 86.800 361.600 87.600 ;
        RECT 356.200 86.200 356.800 86.800 ;
        RECT 356.200 85.600 357.200 86.200 ;
        RECT 356.400 82.200 357.200 85.600 ;
        RECT 359.600 82.200 360.400 86.800 ;
        RECT 362.800 82.200 363.600 85.000 ;
        RECT 364.400 82.200 365.200 85.000 ;
        RECT 366.000 82.200 366.800 87.000 ;
        RECT 369.200 82.200 370.000 87.000 ;
        RECT 372.400 82.200 373.200 88.400 ;
        RECT 380.400 87.600 383.000 88.400 ;
        RECT 375.600 86.800 379.800 87.600 ;
        RECT 374.000 82.200 374.800 85.000 ;
        RECT 375.600 82.200 376.400 85.000 ;
        RECT 377.200 82.200 378.000 85.000 ;
        RECT 380.400 82.200 381.200 87.600 ;
        RECT 385.600 87.400 386.200 89.000 ;
        RECT 383.600 86.800 386.200 87.400 ;
        RECT 386.800 90.000 387.800 90.800 ;
        RECT 383.600 82.200 384.400 86.800 ;
        RECT 386.800 82.200 387.600 90.000 ;
        RECT 388.400 88.300 389.200 88.400 ;
        RECT 390.000 88.300 390.800 90.400 ;
        RECT 388.400 87.700 390.800 88.300 ;
        RECT 388.400 87.600 389.200 87.700 ;
        RECT 391.600 82.200 392.400 95.800 ;
        RECT 393.200 93.600 394.000 95.200 ;
        RECT 393.200 90.300 394.000 90.400 ;
        RECT 394.800 90.300 395.600 90.400 ;
        RECT 393.200 89.700 395.600 90.300 ;
        RECT 393.200 89.600 394.000 89.700 ;
        RECT 394.800 88.800 395.600 89.700 ;
        RECT 396.400 82.200 397.200 95.800 ;
        RECT 401.200 95.800 403.000 96.400 ;
        RECT 406.000 95.800 407.800 96.400 ;
        RECT 409.200 95.800 410.000 99.800 ;
        RECT 410.800 96.000 411.600 99.800 ;
        RECT 414.000 96.000 414.800 99.800 ;
        RECT 410.800 95.800 414.800 96.000 ;
        RECT 398.000 93.600 398.800 95.200 ;
        RECT 399.600 93.600 400.400 95.200 ;
        RECT 401.200 82.200 402.000 95.800 ;
        RECT 404.400 93.600 405.200 95.200 ;
        RECT 406.000 92.300 406.800 95.800 ;
        RECT 409.400 94.400 410.000 95.800 ;
        RECT 411.000 95.400 414.600 95.800 ;
        RECT 415.600 95.600 416.400 97.200 ;
        RECT 413.200 94.400 414.000 94.800 ;
        RECT 409.200 93.600 411.800 94.400 ;
        RECT 413.200 94.300 414.800 94.400 ;
        RECT 417.200 94.300 418.000 99.800 ;
        RECT 413.200 93.800 418.000 94.300 ;
        RECT 414.000 93.700 418.000 93.800 ;
        RECT 414.000 93.600 414.800 93.700 ;
        RECT 406.000 91.700 409.900 92.300 ;
        RECT 402.800 88.800 403.600 90.400 ;
        RECT 406.000 82.200 406.800 91.700 ;
        RECT 409.300 90.400 409.900 91.700 ;
        RECT 407.600 88.800 408.400 90.400 ;
        RECT 409.200 90.200 410.000 90.400 ;
        RECT 411.200 90.200 411.800 93.600 ;
        RECT 412.400 91.600 413.200 93.200 ;
        RECT 409.200 89.600 410.600 90.200 ;
        RECT 411.200 89.600 412.200 90.200 ;
        RECT 410.000 88.400 410.600 89.600 ;
        RECT 410.000 87.600 410.800 88.400 ;
        RECT 411.400 82.200 412.200 89.600 ;
        RECT 417.200 82.200 418.000 93.700 ;
        RECT 418.800 92.400 419.600 99.800 ;
        RECT 422.000 95.200 422.800 99.800 ;
        RECT 430.000 95.600 430.800 97.200 ;
        RECT 420.600 94.600 422.800 95.200 ;
        RECT 418.800 90.200 419.400 92.400 ;
        RECT 420.600 91.600 421.200 94.600 ;
        RECT 420.000 90.800 421.200 91.600 ;
        RECT 420.600 90.200 421.200 90.800 ;
        RECT 418.800 82.200 419.600 90.200 ;
        RECT 420.600 89.600 422.800 90.200 ;
        RECT 422.000 82.200 422.800 89.600 ;
        RECT 431.600 82.200 432.400 99.800 ;
        RECT 433.400 96.400 434.200 97.200 ;
        RECT 433.200 95.600 434.000 96.400 ;
        RECT 434.800 95.800 435.600 99.800 ;
        RECT 433.200 92.200 434.000 92.400 ;
        RECT 435.000 92.200 435.600 95.800 ;
        RECT 436.400 92.800 437.200 94.400 ;
        RECT 443.200 94.200 444.000 99.800 ;
        RECT 448.600 96.400 449.400 99.800 ;
        RECT 447.600 95.800 449.400 96.400 ;
        RECT 443.200 93.800 445.000 94.200 ;
        RECT 443.400 93.600 445.000 93.800 ;
        RECT 446.000 93.600 446.800 95.200 ;
        RECT 438.000 92.200 438.800 92.400 ;
        RECT 433.200 91.600 435.600 92.200 ;
        RECT 437.200 91.600 438.800 92.200 ;
        RECT 441.200 91.600 442.800 92.400 ;
        RECT 433.400 90.200 434.000 91.600 ;
        RECT 437.200 91.200 438.000 91.600 ;
        RECT 433.200 82.200 434.000 90.200 ;
        RECT 434.800 89.600 438.800 90.200 ;
        RECT 439.600 89.600 440.400 91.200 ;
        RECT 444.400 90.400 445.000 93.600 ;
        RECT 444.400 89.600 445.200 90.400 ;
        RECT 434.800 82.200 435.600 89.600 ;
        RECT 438.000 82.200 438.800 89.600 ;
        RECT 441.200 88.300 442.000 88.400 ;
        RECT 442.800 88.300 443.600 89.200 ;
        RECT 441.200 87.700 443.600 88.300 ;
        RECT 441.200 87.600 442.000 87.700 ;
        RECT 442.800 87.600 443.600 87.700 ;
        RECT 444.400 87.000 445.000 89.600 ;
        RECT 441.400 86.400 445.000 87.000 ;
        RECT 441.400 86.200 442.000 86.400 ;
        RECT 441.200 82.200 442.000 86.200 ;
        RECT 444.400 86.200 445.000 86.400 ;
        RECT 444.400 82.200 445.200 86.200 ;
        RECT 447.600 82.200 448.400 95.800 ;
        RECT 450.800 95.200 451.600 99.800 ;
        RECT 450.800 94.600 453.000 95.200 ;
        RECT 452.400 91.600 453.000 94.600 ;
        RECT 454.000 92.400 454.800 99.800 ;
        RECT 459.400 96.000 460.200 99.000 ;
        RECT 463.600 97.000 464.400 99.000 ;
        RECT 458.600 95.400 460.200 96.000 ;
        RECT 458.600 95.000 459.400 95.400 ;
        RECT 458.600 94.400 459.200 95.000 ;
        RECT 463.800 94.800 464.400 97.000 ;
        RECT 468.200 95.800 469.800 99.800 ;
        RECT 475.800 98.400 477.400 99.800 ;
        RECT 474.800 97.600 477.400 98.400 ;
        RECT 475.800 95.800 477.400 97.600 ;
        RECT 482.800 96.000 483.600 99.800 ;
        RECT 457.200 93.600 459.200 94.400 ;
        RECT 460.200 94.200 464.400 94.800 ;
        RECT 460.200 93.800 461.200 94.200 ;
        RECT 452.400 90.800 453.600 91.600 ;
        RECT 449.200 88.800 450.000 90.400 ;
        RECT 452.400 90.200 453.000 90.800 ;
        RECT 454.200 90.200 454.800 92.400 ;
        RECT 455.600 92.300 456.400 92.400 ;
        RECT 457.200 92.300 458.000 92.400 ;
        RECT 455.600 91.700 458.000 92.300 ;
        RECT 455.600 91.600 456.400 91.700 ;
        RECT 457.200 90.800 458.000 91.700 ;
        RECT 450.800 89.600 453.000 90.200 ;
        RECT 450.800 82.200 451.600 89.600 ;
        RECT 454.000 82.200 454.800 90.200 ;
        RECT 458.600 89.800 459.200 93.600 ;
        RECT 459.800 93.000 461.200 93.800 ;
        RECT 460.600 91.000 461.200 93.000 ;
        RECT 462.000 91.600 462.800 93.200 ;
        RECT 463.600 91.600 464.400 93.200 ;
        RECT 466.800 92.800 467.600 94.400 ;
        RECT 468.600 92.400 469.200 95.800 ;
        RECT 470.000 94.300 470.800 94.400 ;
        RECT 471.600 94.300 472.400 94.400 ;
        RECT 474.800 94.300 475.600 94.400 ;
        RECT 470.000 93.700 475.600 94.300 ;
        RECT 470.000 93.600 470.800 93.700 ;
        RECT 471.600 93.600 472.400 93.700 ;
        RECT 474.800 93.600 475.600 93.700 ;
        RECT 470.000 93.200 470.600 93.600 ;
        RECT 469.800 92.400 470.600 93.200 ;
        RECT 475.000 93.200 475.600 93.600 ;
        RECT 475.000 92.400 475.800 93.200 ;
        RECT 476.400 92.400 477.000 95.800 ;
        RECT 482.600 95.200 483.600 96.000 ;
        RECT 478.000 94.300 478.800 94.400 ;
        RECT 482.600 94.300 483.400 95.200 ;
        RECT 484.400 94.600 485.200 99.800 ;
        RECT 490.800 96.600 491.600 99.800 ;
        RECT 492.400 97.000 493.200 99.800 ;
        RECT 494.000 97.000 494.800 99.800 ;
        RECT 495.600 97.000 496.400 99.800 ;
        RECT 497.200 97.000 498.000 99.800 ;
        RECT 500.400 97.000 501.200 99.800 ;
        RECT 503.600 97.000 504.400 99.800 ;
        RECT 505.200 97.000 506.000 99.800 ;
        RECT 506.800 97.000 507.600 99.800 ;
        RECT 489.200 95.800 491.600 96.600 ;
        RECT 508.400 96.600 509.200 99.800 ;
        RECT 489.200 95.200 490.000 95.800 ;
        RECT 478.000 93.700 483.400 94.300 ;
        RECT 478.000 92.800 478.800 93.700 ;
        RECT 465.200 92.200 466.000 92.400 ;
        RECT 465.200 91.600 466.800 92.200 ;
        RECT 468.400 91.600 469.200 92.400 ;
        RECT 466.000 91.200 466.800 91.600 ;
        RECT 468.600 91.400 469.200 91.600 ;
        RECT 460.600 90.400 464.400 91.000 ;
        RECT 468.600 90.800 470.600 91.400 ;
        RECT 471.600 90.800 472.400 92.400 ;
        RECT 473.200 90.800 474.000 92.400 ;
        RECT 476.400 91.600 477.200 92.400 ;
        RECT 479.600 92.200 480.400 92.400 ;
        RECT 478.800 91.600 480.400 92.200 ;
        RECT 476.400 91.400 477.000 91.600 ;
        RECT 475.000 90.800 477.000 91.400 ;
        RECT 478.800 91.200 479.600 91.600 ;
        RECT 482.600 90.800 483.400 93.700 ;
        RECT 484.000 94.000 485.200 94.600 ;
        RECT 488.200 94.600 490.000 95.200 ;
        RECT 494.000 95.600 495.000 96.400 ;
        RECT 498.000 95.600 499.600 96.400 ;
        RECT 500.400 95.800 505.000 96.400 ;
        RECT 508.400 95.800 511.000 96.600 ;
        RECT 500.400 95.600 501.200 95.800 ;
        RECT 484.000 92.000 484.600 94.000 ;
        RECT 488.200 93.400 489.000 94.600 ;
        RECT 485.200 92.600 489.000 93.400 ;
        RECT 494.000 92.800 494.800 95.600 ;
        RECT 500.400 94.800 501.200 95.000 ;
        RECT 496.800 94.200 501.200 94.800 ;
        RECT 496.800 94.000 497.600 94.200 ;
        RECT 502.000 93.600 502.800 95.200 ;
        RECT 504.200 93.400 505.000 95.800 ;
        RECT 510.200 95.200 511.000 95.800 ;
        RECT 510.200 94.400 513.200 95.200 ;
        RECT 514.800 93.800 515.600 99.800 ;
        RECT 518.000 96.000 518.800 99.800 ;
        RECT 497.200 92.600 500.400 93.400 ;
        RECT 504.200 92.600 506.200 93.400 ;
        RECT 506.800 93.000 515.600 93.800 ;
        RECT 490.800 92.000 491.600 92.600 ;
        RECT 508.400 92.000 509.200 92.400 ;
        RECT 511.600 92.000 512.400 92.400 ;
        RECT 513.400 92.000 514.200 92.200 ;
        RECT 484.000 91.400 484.800 92.000 ;
        RECT 490.800 91.400 514.200 92.000 ;
        RECT 458.600 89.200 460.200 89.800 ;
        RECT 459.400 84.400 460.200 89.200 ;
        RECT 463.800 87.000 464.400 90.400 ;
        RECT 470.000 90.200 470.600 90.800 ;
        RECT 475.000 90.200 475.600 90.800 ;
        RECT 459.400 83.600 461.200 84.400 ;
        RECT 459.400 82.200 460.200 83.600 ;
        RECT 463.600 83.000 464.400 87.000 ;
        RECT 465.200 89.600 469.200 90.200 ;
        RECT 465.200 82.200 466.000 89.600 ;
        RECT 468.400 82.800 469.200 89.600 ;
        RECT 470.000 83.400 470.800 90.200 ;
        RECT 471.600 82.800 472.400 90.200 ;
        RECT 468.400 82.200 472.400 82.800 ;
        RECT 473.200 82.800 474.000 90.200 ;
        RECT 474.800 83.400 475.600 90.200 ;
        RECT 476.400 89.600 480.400 90.200 ;
        RECT 482.600 90.000 483.600 90.800 ;
        RECT 476.400 82.800 477.200 89.600 ;
        RECT 473.200 82.200 477.200 82.800 ;
        RECT 479.600 82.200 480.400 89.600 ;
        RECT 482.800 82.200 483.600 90.000 ;
        RECT 484.200 89.600 484.800 91.400 ;
        RECT 484.200 89.000 493.200 89.600 ;
        RECT 484.200 87.400 484.800 89.000 ;
        RECT 492.400 88.800 493.200 89.000 ;
        RECT 495.600 89.000 504.200 89.600 ;
        RECT 495.600 88.800 496.400 89.000 ;
        RECT 487.400 87.600 490.000 88.400 ;
        RECT 484.200 86.800 486.800 87.400 ;
        RECT 486.000 82.200 486.800 86.800 ;
        RECT 489.200 82.200 490.000 87.600 ;
        RECT 490.600 86.800 494.800 87.600 ;
        RECT 492.400 82.200 493.200 85.000 ;
        RECT 494.000 82.200 494.800 85.000 ;
        RECT 495.600 82.200 496.400 85.000 ;
        RECT 497.200 82.200 498.000 88.400 ;
        RECT 500.400 87.600 503.000 88.400 ;
        RECT 503.600 88.200 504.200 89.000 ;
        RECT 505.200 89.400 506.000 89.600 ;
        RECT 505.200 89.000 510.600 89.400 ;
        RECT 505.200 88.800 511.400 89.000 ;
        RECT 510.000 88.200 511.400 88.800 ;
        RECT 503.600 87.600 509.400 88.200 ;
        RECT 512.400 88.000 514.000 88.800 ;
        RECT 512.400 87.600 513.000 88.000 ;
        RECT 500.400 82.200 501.200 87.000 ;
        RECT 503.600 82.200 504.400 87.000 ;
        RECT 508.800 86.800 513.000 87.600 ;
        RECT 514.800 87.400 515.600 93.000 ;
        RECT 517.800 95.200 518.800 96.000 ;
        RECT 517.800 90.800 518.600 95.200 ;
        RECT 519.600 94.600 520.400 99.800 ;
        RECT 526.000 96.600 526.800 99.800 ;
        RECT 527.600 97.000 528.400 99.800 ;
        RECT 529.200 97.000 530.000 99.800 ;
        RECT 530.800 97.000 531.600 99.800 ;
        RECT 532.400 97.000 533.200 99.800 ;
        RECT 535.600 97.000 536.400 99.800 ;
        RECT 538.800 97.000 539.600 99.800 ;
        RECT 540.400 97.000 541.200 99.800 ;
        RECT 542.000 97.000 542.800 99.800 ;
        RECT 524.400 95.800 526.800 96.600 ;
        RECT 543.600 96.600 544.400 99.800 ;
        RECT 524.400 95.200 525.200 95.800 ;
        RECT 519.200 94.000 520.400 94.600 ;
        RECT 523.400 94.600 525.200 95.200 ;
        RECT 529.200 95.600 530.200 96.400 ;
        RECT 533.200 95.600 534.800 96.400 ;
        RECT 535.600 95.800 540.200 96.400 ;
        RECT 543.600 95.800 546.200 96.600 ;
        RECT 535.600 95.600 536.400 95.800 ;
        RECT 519.200 92.000 519.800 94.000 ;
        RECT 523.400 93.400 524.200 94.600 ;
        RECT 520.400 92.600 524.200 93.400 ;
        RECT 529.200 92.800 530.000 95.600 ;
        RECT 535.600 94.800 536.400 95.000 ;
        RECT 532.000 94.200 536.400 94.800 ;
        RECT 532.000 94.000 532.800 94.200 ;
        RECT 537.200 93.600 538.000 95.200 ;
        RECT 539.400 93.400 540.200 95.800 ;
        RECT 545.400 95.200 546.200 95.800 ;
        RECT 545.400 94.400 548.400 95.200 ;
        RECT 550.000 93.800 550.800 99.800 ;
        RECT 532.400 92.600 535.600 93.400 ;
        RECT 539.400 92.600 541.400 93.400 ;
        RECT 542.000 93.000 550.800 93.800 ;
        RECT 526.000 92.000 526.800 92.600 ;
        RECT 543.600 92.000 544.400 92.400 ;
        RECT 545.200 92.000 546.000 92.400 ;
        RECT 548.600 92.000 549.400 92.200 ;
        RECT 519.200 91.400 520.000 92.000 ;
        RECT 526.000 91.400 549.400 92.000 ;
        RECT 517.800 90.000 518.800 90.800 ;
        RECT 513.600 86.800 515.600 87.400 ;
        RECT 505.200 82.200 506.000 85.000 ;
        RECT 506.800 82.200 507.600 85.000 ;
        RECT 510.000 82.200 510.800 86.800 ;
        RECT 513.600 86.200 514.200 86.800 ;
        RECT 513.200 85.600 514.200 86.200 ;
        RECT 513.200 82.200 514.000 85.600 ;
        RECT 518.000 82.200 518.800 90.000 ;
        RECT 519.400 89.600 520.000 91.400 ;
        RECT 519.400 89.000 528.400 89.600 ;
        RECT 519.400 87.400 520.000 89.000 ;
        RECT 527.600 88.800 528.400 89.000 ;
        RECT 530.800 89.000 539.400 89.600 ;
        RECT 530.800 88.800 531.600 89.000 ;
        RECT 522.600 87.600 525.200 88.400 ;
        RECT 519.400 86.800 522.000 87.400 ;
        RECT 521.200 82.200 522.000 86.800 ;
        RECT 524.400 82.200 525.200 87.600 ;
        RECT 525.800 86.800 530.000 87.600 ;
        RECT 527.600 82.200 528.400 85.000 ;
        RECT 529.200 82.200 530.000 85.000 ;
        RECT 530.800 82.200 531.600 85.000 ;
        RECT 532.400 82.200 533.200 88.400 ;
        RECT 535.600 87.600 538.200 88.400 ;
        RECT 538.800 88.200 539.400 89.000 ;
        RECT 540.400 89.400 541.200 89.600 ;
        RECT 540.400 89.000 545.800 89.400 ;
        RECT 540.400 88.800 546.600 89.000 ;
        RECT 545.200 88.200 546.600 88.800 ;
        RECT 538.800 87.600 544.600 88.200 ;
        RECT 547.600 88.000 549.200 88.800 ;
        RECT 547.600 87.600 548.200 88.000 ;
        RECT 535.600 82.200 536.400 87.000 ;
        RECT 538.800 82.200 539.600 87.000 ;
        RECT 544.000 86.800 548.200 87.600 ;
        RECT 550.000 87.400 550.800 93.000 ;
        RECT 548.800 86.800 550.800 87.400 ;
        RECT 540.400 82.200 541.200 85.000 ;
        RECT 542.000 82.200 542.800 85.000 ;
        RECT 545.200 82.200 546.000 86.800 ;
        RECT 548.800 86.200 549.400 86.800 ;
        RECT 548.400 85.600 549.400 86.200 ;
        RECT 548.400 82.200 549.200 85.600 ;
        RECT 3.800 78.400 4.600 79.800 ;
        RECT 2.800 77.600 4.600 78.400 ;
        RECT 3.800 72.600 4.600 77.600 ;
        RECT 2.800 71.800 4.600 72.600 ;
        RECT 3.000 68.400 3.600 71.800 ;
        RECT 4.400 69.600 5.200 71.200 ;
        RECT 7.600 70.300 8.400 79.800 ;
        RECT 11.800 72.600 12.600 79.800 ;
        RECT 10.800 71.800 12.600 72.600 ;
        RECT 14.600 78.400 15.400 79.800 ;
        RECT 14.600 77.600 16.400 78.400 ;
        RECT 14.600 72.600 15.400 77.600 ;
        RECT 14.600 71.800 16.400 72.600 ;
        RECT 9.200 70.300 10.000 70.400 ;
        RECT 7.600 69.700 10.000 70.300 ;
        RECT 2.800 67.600 3.600 68.400 ;
        RECT 3.000 66.400 3.600 67.600 ;
        RECT 1.200 64.800 2.000 66.400 ;
        RECT 2.800 65.600 3.600 66.400 ;
        RECT 3.000 64.200 3.600 65.600 ;
        RECT 6.000 64.800 6.800 66.400 ;
        RECT 2.800 62.200 3.600 64.200 ;
        RECT 7.600 62.200 8.400 69.700 ;
        RECT 9.200 69.600 10.000 69.700 ;
        RECT 11.000 68.400 11.600 71.800 ;
        RECT 12.400 70.300 13.200 71.200 ;
        RECT 14.000 70.300 14.800 71.200 ;
        RECT 12.400 69.700 14.800 70.300 ;
        RECT 12.400 69.600 13.200 69.700 ;
        RECT 14.000 69.600 14.800 69.700 ;
        RECT 15.600 68.400 16.200 71.800 ;
        RECT 20.400 70.300 21.200 79.800 ;
        RECT 22.600 78.400 23.400 79.800 ;
        RECT 27.400 78.400 28.200 79.800 ;
        RECT 22.600 77.600 24.400 78.400 ;
        RECT 26.800 77.600 28.200 78.400 ;
        RECT 22.600 72.600 23.400 77.600 ;
        RECT 27.400 72.600 28.200 77.600 ;
        RECT 32.200 72.600 33.000 79.800 ;
        RECT 22.600 71.800 24.400 72.600 ;
        RECT 27.400 71.800 29.200 72.600 ;
        RECT 32.200 71.800 34.000 72.600 ;
        RECT 22.000 70.300 22.800 71.200 ;
        RECT 20.400 69.700 22.800 70.300 ;
        RECT 10.800 68.300 11.600 68.400 ;
        RECT 14.000 68.300 14.800 68.400 ;
        RECT 10.800 67.700 14.800 68.300 ;
        RECT 10.800 67.600 11.600 67.700 ;
        RECT 14.000 67.600 14.800 67.700 ;
        RECT 15.600 67.600 16.400 68.400 ;
        RECT 9.200 64.800 10.000 66.400 ;
        RECT 11.000 64.200 11.600 67.600 ;
        RECT 10.800 62.200 11.600 64.200 ;
        RECT 15.600 64.200 16.200 67.600 ;
        RECT 17.200 64.800 18.000 66.400 ;
        RECT 18.800 64.800 19.600 66.400 ;
        RECT 15.600 62.200 16.400 64.200 ;
        RECT 20.400 62.200 21.200 69.700 ;
        RECT 22.000 69.600 22.800 69.700 ;
        RECT 23.600 68.400 24.200 71.800 ;
        RECT 26.800 69.600 27.600 71.200 ;
        RECT 28.400 68.400 29.000 71.800 ;
        RECT 31.600 69.600 32.400 71.200 ;
        RECT 33.200 68.400 33.800 71.800 ;
        RECT 36.400 71.600 37.200 73.200 ;
        RECT 23.600 67.600 24.400 68.400 ;
        RECT 28.400 67.600 29.200 68.400 ;
        RECT 30.000 68.300 30.800 68.400 ;
        RECT 33.200 68.300 34.000 68.400 ;
        RECT 30.000 67.700 34.000 68.300 ;
        RECT 30.000 67.600 30.800 67.700 ;
        RECT 33.200 67.600 34.000 67.700 ;
        RECT 23.600 64.200 24.200 67.600 ;
        RECT 25.200 64.800 26.000 66.400 ;
        RECT 28.400 64.200 29.000 67.600 ;
        RECT 30.000 64.800 30.800 66.400 ;
        RECT 33.200 64.200 33.800 67.600 ;
        RECT 34.800 64.800 35.600 66.400 ;
        RECT 38.000 66.200 38.800 79.800 ;
        RECT 39.600 72.300 40.400 72.400 ;
        RECT 41.200 72.300 42.000 79.800 ;
        RECT 39.600 71.700 42.000 72.300 ;
        RECT 47.000 71.800 49.000 79.800 ;
        RECT 55.000 72.400 55.800 79.800 ;
        RECT 56.400 73.600 57.200 74.400 ;
        RECT 56.600 72.400 57.200 73.600 ;
        RECT 55.000 71.800 56.000 72.400 ;
        RECT 56.600 71.800 58.000 72.400 ;
        RECT 39.600 71.600 40.400 71.700 ;
        RECT 39.600 66.800 40.400 68.400 ;
        RECT 37.000 65.600 38.800 66.200 ;
        RECT 37.000 64.400 37.800 65.600 ;
        RECT 23.600 62.200 24.400 64.200 ;
        RECT 28.400 62.200 29.200 64.200 ;
        RECT 33.200 62.200 34.000 64.200 ;
        RECT 36.400 63.600 37.800 64.400 ;
        RECT 37.000 62.200 37.800 63.600 ;
        RECT 41.200 62.200 42.000 71.700 ;
        RECT 46.000 68.800 46.800 70.400 ;
        RECT 47.600 68.400 48.200 71.800 ;
        RECT 49.200 68.800 50.000 70.400 ;
        RECT 44.400 68.200 45.200 68.400 ;
        RECT 47.600 68.200 48.400 68.400 ;
        RECT 44.400 67.600 46.000 68.200 ;
        RECT 47.600 67.600 50.000 68.200 ;
        RECT 50.800 67.600 51.600 69.200 ;
        RECT 54.000 68.800 54.800 70.400 ;
        RECT 55.400 68.400 56.000 71.800 ;
        RECT 57.200 71.600 58.000 71.800 ;
        RECT 58.800 71.600 59.600 73.200 ;
        RECT 57.300 70.300 57.900 71.600 ;
        RECT 60.400 70.300 61.200 79.800 ;
        RECT 65.200 71.200 66.000 79.800 ;
        RECT 68.400 71.200 69.200 79.800 ;
        RECT 71.600 71.200 72.400 79.800 ;
        RECT 74.800 71.200 75.600 79.800 ;
        RECT 79.600 75.800 80.400 79.800 ;
        RECT 79.800 75.600 80.400 75.800 ;
        RECT 82.800 75.800 83.600 79.800 ;
        RECT 84.400 75.800 85.200 79.800 ;
        RECT 82.800 75.600 83.400 75.800 ;
        RECT 79.800 75.000 83.400 75.600 ;
        RECT 81.200 72.800 82.000 74.400 ;
        RECT 82.800 72.400 83.400 75.000 ;
        RECT 84.600 75.600 85.200 75.800 ;
        RECT 87.600 75.800 88.400 79.800 ;
        RECT 87.600 75.600 88.200 75.800 ;
        RECT 84.600 75.000 88.200 75.600 ;
        RECT 84.600 72.400 85.200 75.000 ;
        RECT 86.000 72.800 86.800 74.400 ;
        RECT 57.300 69.700 61.200 70.300 ;
        RECT 52.400 68.200 53.200 68.400 ;
        RECT 52.400 67.600 54.000 68.200 ;
        RECT 55.400 67.600 58.000 68.400 ;
        RECT 45.200 67.200 46.000 67.600 ;
        RECT 42.800 64.800 43.600 66.400 ;
        RECT 44.600 66.200 48.200 66.600 ;
        RECT 49.400 66.200 50.000 67.600 ;
        RECT 53.200 67.200 54.000 67.600 ;
        RECT 52.600 66.200 56.200 66.600 ;
        RECT 57.200 66.200 57.800 67.600 ;
        RECT 60.400 66.200 61.200 69.700 ;
        RECT 63.600 70.400 66.000 71.200 ;
        RECT 67.000 70.400 69.200 71.200 ;
        RECT 70.200 70.400 72.400 71.200 ;
        RECT 73.800 70.400 75.600 71.200 ;
        RECT 62.000 66.800 62.800 68.400 ;
        RECT 63.600 67.600 64.400 70.400 ;
        RECT 67.000 69.000 67.800 70.400 ;
        RECT 70.200 69.000 71.000 70.400 ;
        RECT 73.800 69.000 74.600 70.400 ;
        RECT 76.400 70.300 77.200 70.400 ;
        RECT 78.000 70.300 78.800 72.400 ;
        RECT 82.800 71.600 83.600 72.400 ;
        RECT 84.400 71.600 85.200 72.400 ;
        RECT 76.400 69.700 78.800 70.300 ;
        RECT 76.400 69.600 77.200 69.700 ;
        RECT 79.600 69.600 81.200 70.400 ;
        RECT 65.200 68.200 67.800 69.000 ;
        RECT 68.600 68.200 71.000 69.000 ;
        RECT 72.000 68.200 74.600 69.000 ;
        RECT 82.800 68.400 83.400 71.600 ;
        RECT 81.800 68.200 83.400 68.400 ;
        RECT 67.000 67.600 67.800 68.200 ;
        RECT 70.200 67.600 71.000 68.200 ;
        RECT 73.800 67.600 74.600 68.200 ;
        RECT 81.600 67.800 83.400 68.200 ;
        RECT 84.600 68.400 85.200 71.600 ;
        RECT 86.800 69.600 88.400 70.400 ;
        RECT 89.200 70.300 90.000 72.400 ;
        RECT 92.400 72.000 93.200 79.800 ;
        RECT 95.600 75.200 96.400 79.800 ;
        RECT 92.200 71.200 93.200 72.000 ;
        RECT 93.800 74.600 96.400 75.200 ;
        RECT 93.800 73.000 94.400 74.600 ;
        RECT 98.800 74.400 99.600 79.800 ;
        RECT 102.000 77.000 102.800 79.800 ;
        RECT 103.600 77.000 104.400 79.800 ;
        RECT 105.200 77.000 106.000 79.800 ;
        RECT 100.200 74.400 104.400 75.200 ;
        RECT 97.000 73.600 99.600 74.400 ;
        RECT 106.800 73.600 107.600 79.800 ;
        RECT 110.000 75.000 110.800 79.800 ;
        RECT 113.200 75.000 114.000 79.800 ;
        RECT 114.800 77.000 115.600 79.800 ;
        RECT 116.400 77.000 117.200 79.800 ;
        RECT 119.600 75.200 120.400 79.800 ;
        RECT 122.800 76.400 123.600 79.800 ;
        RECT 122.800 75.800 123.800 76.400 ;
        RECT 123.200 75.200 123.800 75.800 ;
        RECT 118.400 74.400 122.600 75.200 ;
        RECT 123.200 74.600 125.200 75.200 ;
        RECT 110.000 73.600 112.600 74.400 ;
        RECT 113.200 73.800 119.000 74.400 ;
        RECT 122.000 74.000 122.600 74.400 ;
        RECT 102.000 73.000 102.800 73.200 ;
        RECT 93.800 72.400 102.800 73.000 ;
        RECT 105.200 73.000 106.000 73.200 ;
        RECT 113.200 73.000 113.800 73.800 ;
        RECT 119.600 73.200 121.000 73.800 ;
        RECT 122.000 73.200 123.600 74.000 ;
        RECT 105.200 72.400 113.800 73.000 ;
        RECT 114.800 73.000 121.000 73.200 ;
        RECT 114.800 72.600 120.200 73.000 ;
        RECT 114.800 72.400 115.600 72.600 ;
        RECT 92.200 70.300 93.000 71.200 ;
        RECT 93.800 70.600 94.400 72.400 ;
        RECT 89.200 69.700 93.000 70.300 ;
        RECT 84.600 68.200 86.200 68.400 ;
        RECT 84.600 67.800 86.400 68.200 ;
        RECT 63.600 66.800 66.000 67.600 ;
        RECT 67.000 66.800 69.200 67.600 ;
        RECT 70.200 66.800 72.400 67.600 ;
        RECT 73.800 66.800 75.600 67.600 ;
        RECT 44.400 66.000 48.400 66.200 ;
        RECT 44.400 62.200 45.200 66.000 ;
        RECT 47.600 62.800 48.400 66.000 ;
        RECT 49.200 63.400 50.000 66.200 ;
        RECT 50.800 62.800 51.600 66.200 ;
        RECT 47.600 62.200 51.600 62.800 ;
        RECT 52.400 66.000 56.400 66.200 ;
        RECT 52.400 62.200 53.200 66.000 ;
        RECT 55.600 62.200 56.400 66.000 ;
        RECT 57.200 62.200 58.000 66.200 ;
        RECT 59.400 65.600 61.200 66.200 ;
        RECT 59.400 62.200 60.200 65.600 ;
        RECT 65.200 62.200 66.000 66.800 ;
        RECT 68.400 62.200 69.200 66.800 ;
        RECT 71.600 62.200 72.400 66.800 ;
        RECT 74.800 62.200 75.600 66.800 ;
        RECT 81.600 62.200 82.400 67.800 ;
        RECT 85.600 62.200 86.400 67.800 ;
        RECT 92.200 66.800 93.000 69.700 ;
        RECT 93.600 70.000 94.400 70.600 ;
        RECT 100.400 70.000 123.800 70.600 ;
        RECT 93.600 68.000 94.200 70.000 ;
        RECT 100.400 69.400 101.200 70.000 ;
        RECT 118.000 69.600 118.800 70.000 ;
        RECT 119.600 69.600 120.400 70.000 ;
        RECT 123.000 69.800 123.800 70.000 ;
        RECT 94.800 68.600 98.600 69.400 ;
        RECT 93.600 67.400 94.800 68.000 ;
        RECT 92.200 66.000 93.200 66.800 ;
        RECT 92.400 62.200 93.200 66.000 ;
        RECT 94.000 62.200 94.800 67.400 ;
        RECT 97.800 67.400 98.600 68.600 ;
        RECT 97.800 66.800 99.600 67.400 ;
        RECT 98.800 66.200 99.600 66.800 ;
        RECT 103.600 66.400 104.400 69.200 ;
        RECT 106.800 68.600 110.000 69.400 ;
        RECT 113.800 68.600 115.800 69.400 ;
        RECT 124.400 69.000 125.200 74.600 ;
        RECT 134.000 72.000 134.800 79.800 ;
        RECT 137.200 75.200 138.000 79.800 ;
        RECT 106.400 67.800 107.200 68.000 ;
        RECT 106.400 67.200 110.800 67.800 ;
        RECT 110.000 67.000 110.800 67.200 ;
        RECT 111.600 66.800 112.400 68.400 ;
        RECT 98.800 65.400 101.200 66.200 ;
        RECT 103.600 65.600 104.600 66.400 ;
        RECT 107.600 65.600 109.200 66.400 ;
        RECT 110.000 66.200 110.800 66.400 ;
        RECT 113.800 66.200 114.600 68.600 ;
        RECT 116.400 68.200 125.200 69.000 ;
        RECT 119.800 66.800 122.800 67.600 ;
        RECT 119.800 66.200 120.600 66.800 ;
        RECT 110.000 65.600 114.600 66.200 ;
        RECT 100.400 62.200 101.200 65.400 ;
        RECT 118.000 65.400 120.600 66.200 ;
        RECT 102.000 62.200 102.800 65.000 ;
        RECT 103.600 62.200 104.400 65.000 ;
        RECT 105.200 62.200 106.000 65.000 ;
        RECT 106.800 62.200 107.600 65.000 ;
        RECT 110.000 62.200 110.800 65.000 ;
        RECT 113.200 62.200 114.000 65.000 ;
        RECT 114.800 62.200 115.600 65.000 ;
        RECT 116.400 62.200 117.200 65.000 ;
        RECT 118.000 62.200 118.800 65.400 ;
        RECT 124.400 62.200 125.200 68.200 ;
        RECT 133.800 71.200 134.800 72.000 ;
        RECT 135.400 74.600 138.000 75.200 ;
        RECT 135.400 73.000 136.000 74.600 ;
        RECT 140.400 74.400 141.200 79.800 ;
        RECT 143.600 77.000 144.400 79.800 ;
        RECT 145.200 77.000 146.000 79.800 ;
        RECT 146.800 77.000 147.600 79.800 ;
        RECT 141.800 74.400 146.000 75.200 ;
        RECT 138.600 73.600 141.200 74.400 ;
        RECT 148.400 73.600 149.200 79.800 ;
        RECT 151.600 75.000 152.400 79.800 ;
        RECT 154.800 75.000 155.600 79.800 ;
        RECT 156.400 77.000 157.200 79.800 ;
        RECT 158.000 77.000 158.800 79.800 ;
        RECT 161.200 75.200 162.000 79.800 ;
        RECT 164.400 76.400 165.200 79.800 ;
        RECT 164.400 75.800 165.400 76.400 ;
        RECT 164.800 75.200 165.400 75.800 ;
        RECT 160.000 74.400 164.200 75.200 ;
        RECT 164.800 74.600 166.800 75.200 ;
        RECT 151.600 73.600 154.200 74.400 ;
        RECT 154.800 73.800 160.600 74.400 ;
        RECT 163.600 74.000 164.200 74.400 ;
        RECT 143.600 73.000 144.400 73.200 ;
        RECT 135.400 72.400 144.400 73.000 ;
        RECT 146.800 73.000 147.600 73.200 ;
        RECT 154.800 73.000 155.400 73.800 ;
        RECT 161.200 73.200 162.600 73.800 ;
        RECT 163.600 73.200 165.200 74.000 ;
        RECT 146.800 72.400 155.400 73.000 ;
        RECT 156.400 73.000 162.600 73.200 ;
        RECT 156.400 72.600 161.800 73.000 ;
        RECT 156.400 72.400 157.200 72.600 ;
        RECT 133.800 66.800 134.600 71.200 ;
        RECT 135.400 70.600 136.000 72.400 ;
        RECT 159.400 71.800 160.200 72.000 ;
        RECT 162.800 71.800 163.600 72.400 ;
        RECT 136.600 71.200 163.600 71.800 ;
        RECT 136.600 71.000 137.400 71.200 ;
        RECT 135.200 70.000 136.000 70.600 ;
        RECT 135.200 68.000 135.800 70.000 ;
        RECT 136.400 68.600 140.200 69.400 ;
        RECT 135.200 67.400 136.400 68.000 ;
        RECT 133.800 66.000 134.800 66.800 ;
        RECT 134.000 62.200 134.800 66.000 ;
        RECT 135.600 62.200 136.400 67.400 ;
        RECT 139.400 67.400 140.200 68.600 ;
        RECT 139.400 66.800 141.200 67.400 ;
        RECT 140.400 66.200 141.200 66.800 ;
        RECT 145.200 66.400 146.000 69.200 ;
        RECT 148.400 68.600 151.600 69.400 ;
        RECT 155.400 68.600 157.400 69.400 ;
        RECT 166.000 69.000 166.800 74.600 ;
        RECT 148.000 67.800 148.800 68.000 ;
        RECT 148.000 67.200 152.400 67.800 ;
        RECT 151.600 67.000 152.400 67.200 ;
        RECT 153.200 66.800 154.000 68.400 ;
        RECT 140.400 65.400 142.800 66.200 ;
        RECT 145.200 65.600 146.200 66.400 ;
        RECT 149.200 65.600 150.800 66.400 ;
        RECT 151.600 66.200 152.400 66.400 ;
        RECT 155.400 66.200 156.200 68.600 ;
        RECT 158.000 68.200 166.800 69.000 ;
        RECT 161.400 66.800 164.400 67.600 ;
        RECT 161.400 66.200 162.200 66.800 ;
        RECT 151.600 65.600 156.200 66.200 ;
        RECT 142.000 62.200 142.800 65.400 ;
        RECT 159.600 65.400 162.200 66.200 ;
        RECT 143.600 62.200 144.400 65.000 ;
        RECT 145.200 62.200 146.000 65.000 ;
        RECT 146.800 62.200 147.600 65.000 ;
        RECT 148.400 62.200 149.200 65.000 ;
        RECT 151.600 62.200 152.400 65.000 ;
        RECT 154.800 62.200 155.600 65.000 ;
        RECT 156.400 62.200 157.200 65.000 ;
        RECT 158.000 62.200 158.800 65.000 ;
        RECT 159.600 62.200 160.400 65.400 ;
        RECT 166.000 62.200 166.800 68.200 ;
        RECT 167.600 71.800 168.400 79.800 ;
        RECT 170.800 72.400 171.600 79.800 ;
        RECT 174.000 76.400 174.800 79.800 ;
        RECT 173.800 75.800 174.800 76.400 ;
        RECT 173.800 75.200 174.400 75.800 ;
        RECT 177.200 75.200 178.000 79.800 ;
        RECT 180.400 77.000 181.200 79.800 ;
        RECT 182.000 77.000 182.800 79.800 ;
        RECT 169.400 71.800 171.600 72.400 ;
        RECT 172.400 74.600 174.400 75.200 ;
        RECT 167.600 69.600 168.200 71.800 ;
        RECT 169.400 71.200 170.000 71.800 ;
        RECT 168.800 70.400 170.000 71.200 ;
        RECT 167.600 62.200 168.400 69.600 ;
        RECT 169.400 67.400 170.000 70.400 ;
        RECT 172.400 69.000 173.200 74.600 ;
        RECT 175.000 74.400 179.200 75.200 ;
        RECT 183.600 75.000 184.400 79.800 ;
        RECT 186.800 75.000 187.600 79.800 ;
        RECT 175.000 74.000 175.600 74.400 ;
        RECT 174.000 73.200 175.600 74.000 ;
        RECT 178.600 73.800 184.400 74.400 ;
        RECT 176.600 73.200 178.000 73.800 ;
        RECT 176.600 73.000 182.800 73.200 ;
        RECT 177.400 72.600 182.800 73.000 ;
        RECT 182.000 72.400 182.800 72.600 ;
        RECT 183.800 73.000 184.400 73.800 ;
        RECT 185.000 73.600 187.600 74.400 ;
        RECT 190.000 73.600 190.800 79.800 ;
        RECT 191.600 77.000 192.400 79.800 ;
        RECT 193.200 77.000 194.000 79.800 ;
        RECT 194.800 77.000 195.600 79.800 ;
        RECT 193.200 74.400 197.400 75.200 ;
        RECT 198.000 74.400 198.800 79.800 ;
        RECT 201.200 75.200 202.000 79.800 ;
        RECT 201.200 74.600 203.800 75.200 ;
        RECT 198.000 73.600 200.600 74.400 ;
        RECT 191.600 73.000 192.400 73.200 ;
        RECT 183.800 72.400 192.400 73.000 ;
        RECT 194.800 73.000 195.600 73.200 ;
        RECT 203.200 73.000 203.800 74.600 ;
        RECT 194.800 72.400 203.800 73.000 ;
        RECT 203.200 70.600 203.800 72.400 ;
        RECT 204.400 72.000 205.200 79.800 ;
        RECT 209.200 72.000 210.000 79.800 ;
        RECT 212.400 75.200 213.200 79.800 ;
        RECT 204.400 71.200 205.400 72.000 ;
        RECT 173.800 70.000 197.200 70.600 ;
        RECT 203.200 70.000 204.000 70.600 ;
        RECT 173.800 69.800 174.600 70.000 ;
        RECT 177.200 69.600 178.000 70.000 ;
        RECT 178.800 69.600 179.600 70.000 ;
        RECT 196.400 69.400 197.200 70.000 ;
        RECT 172.400 68.200 181.200 69.000 ;
        RECT 181.800 68.600 183.800 69.400 ;
        RECT 187.600 68.600 190.800 69.400 ;
        RECT 169.400 66.800 171.600 67.400 ;
        RECT 170.800 62.200 171.600 66.800 ;
        RECT 172.400 62.200 173.200 68.200 ;
        RECT 174.800 66.800 177.800 67.600 ;
        RECT 177.000 66.200 177.800 66.800 ;
        RECT 183.000 66.200 183.800 68.600 ;
        RECT 185.200 66.800 186.000 68.400 ;
        RECT 190.400 67.800 191.200 68.000 ;
        RECT 186.800 67.200 191.200 67.800 ;
        RECT 186.800 67.000 187.600 67.200 ;
        RECT 193.200 66.400 194.000 69.200 ;
        RECT 199.000 68.600 202.800 69.400 ;
        RECT 199.000 67.400 199.800 68.600 ;
        RECT 203.400 68.000 204.000 70.000 ;
        RECT 186.800 66.200 187.600 66.400 ;
        RECT 177.000 65.400 179.600 66.200 ;
        RECT 183.000 65.600 187.600 66.200 ;
        RECT 188.400 65.600 190.000 66.400 ;
        RECT 193.000 65.600 194.000 66.400 ;
        RECT 198.000 66.800 199.800 67.400 ;
        RECT 202.800 67.400 204.000 68.000 ;
        RECT 198.000 66.200 198.800 66.800 ;
        RECT 178.800 62.200 179.600 65.400 ;
        RECT 196.400 65.400 198.800 66.200 ;
        RECT 180.400 62.200 181.200 65.000 ;
        RECT 182.000 62.200 182.800 65.000 ;
        RECT 183.600 62.200 184.400 65.000 ;
        RECT 186.800 62.200 187.600 65.000 ;
        RECT 190.000 62.200 190.800 65.000 ;
        RECT 191.600 62.200 192.400 65.000 ;
        RECT 193.200 62.200 194.000 65.000 ;
        RECT 194.800 62.200 195.600 65.000 ;
        RECT 196.400 62.200 197.200 65.400 ;
        RECT 202.800 62.200 203.600 67.400 ;
        RECT 204.600 66.800 205.400 71.200 ;
        RECT 204.400 66.000 205.400 66.800 ;
        RECT 209.000 71.200 210.000 72.000 ;
        RECT 210.600 74.600 213.200 75.200 ;
        RECT 210.600 73.000 211.200 74.600 ;
        RECT 215.600 74.400 216.400 79.800 ;
        RECT 218.800 77.000 219.600 79.800 ;
        RECT 220.400 77.000 221.200 79.800 ;
        RECT 222.000 77.000 222.800 79.800 ;
        RECT 217.000 74.400 221.200 75.200 ;
        RECT 213.800 73.600 216.400 74.400 ;
        RECT 223.600 73.600 224.400 79.800 ;
        RECT 226.800 75.000 227.600 79.800 ;
        RECT 230.000 75.000 230.800 79.800 ;
        RECT 231.600 77.000 232.400 79.800 ;
        RECT 233.200 77.000 234.000 79.800 ;
        RECT 236.400 75.200 237.200 79.800 ;
        RECT 239.600 76.400 240.400 79.800 ;
        RECT 239.600 75.800 240.600 76.400 ;
        RECT 240.000 75.200 240.600 75.800 ;
        RECT 235.200 74.400 239.400 75.200 ;
        RECT 240.000 74.600 242.000 75.200 ;
        RECT 226.800 73.600 229.400 74.400 ;
        RECT 230.000 73.800 235.800 74.400 ;
        RECT 238.800 74.000 239.400 74.400 ;
        RECT 218.800 73.000 219.600 73.200 ;
        RECT 210.600 72.400 219.600 73.000 ;
        RECT 222.000 73.000 222.800 73.200 ;
        RECT 230.000 73.000 230.600 73.800 ;
        RECT 236.400 73.200 237.800 73.800 ;
        RECT 238.800 73.200 240.400 74.000 ;
        RECT 222.000 72.400 230.600 73.000 ;
        RECT 231.600 73.000 237.800 73.200 ;
        RECT 231.600 72.600 237.000 73.000 ;
        RECT 231.600 72.400 232.400 72.600 ;
        RECT 209.000 66.800 209.800 71.200 ;
        RECT 210.600 70.600 211.200 72.400 ;
        RECT 210.400 70.000 211.200 70.600 ;
        RECT 217.200 70.000 240.600 70.600 ;
        RECT 210.400 68.000 211.000 70.000 ;
        RECT 217.200 69.400 218.000 70.000 ;
        RECT 234.800 69.600 235.600 70.000 ;
        RECT 239.600 69.800 240.600 70.000 ;
        RECT 239.600 69.600 240.400 69.800 ;
        RECT 211.600 68.600 215.400 69.400 ;
        RECT 210.400 67.400 211.600 68.000 ;
        RECT 209.000 66.000 210.000 66.800 ;
        RECT 204.400 62.200 205.200 66.000 ;
        RECT 209.200 62.200 210.000 66.000 ;
        RECT 210.800 62.200 211.600 67.400 ;
        RECT 214.600 67.400 215.400 68.600 ;
        RECT 214.600 66.800 216.400 67.400 ;
        RECT 215.600 66.200 216.400 66.800 ;
        RECT 220.400 66.400 221.200 69.200 ;
        RECT 223.600 68.600 226.800 69.400 ;
        RECT 230.600 68.600 232.600 69.400 ;
        RECT 241.200 69.000 242.000 74.600 ;
        RECT 223.200 67.800 224.000 68.000 ;
        RECT 223.200 67.200 227.600 67.800 ;
        RECT 226.800 67.000 227.600 67.200 ;
        RECT 228.400 66.800 229.200 68.400 ;
        RECT 215.600 65.400 218.000 66.200 ;
        RECT 220.400 65.600 221.400 66.400 ;
        RECT 224.400 65.600 226.000 66.400 ;
        RECT 226.800 66.200 227.600 66.400 ;
        RECT 230.600 66.200 231.400 68.600 ;
        RECT 233.200 68.200 242.000 69.000 ;
        RECT 236.600 66.800 239.600 67.600 ;
        RECT 236.600 66.200 237.400 66.800 ;
        RECT 226.800 65.600 231.400 66.200 ;
        RECT 217.200 62.200 218.000 65.400 ;
        RECT 234.800 65.400 237.400 66.200 ;
        RECT 218.800 62.200 219.600 65.000 ;
        RECT 220.400 62.200 221.200 65.000 ;
        RECT 222.000 62.200 222.800 65.000 ;
        RECT 223.600 62.200 224.400 65.000 ;
        RECT 226.800 62.200 227.600 65.000 ;
        RECT 230.000 62.200 230.800 65.000 ;
        RECT 231.600 62.200 232.400 65.000 ;
        RECT 233.200 62.200 234.000 65.000 ;
        RECT 234.800 62.200 235.600 65.400 ;
        RECT 241.200 62.200 242.000 68.200 ;
        RECT 242.800 71.800 243.600 79.800 ;
        RECT 246.000 72.400 246.800 79.800 ;
        RECT 244.600 71.800 246.800 72.400 ;
        RECT 242.800 69.600 243.400 71.800 ;
        RECT 244.600 71.200 245.200 71.800 ;
        RECT 244.000 70.400 245.200 71.200 ;
        RECT 242.800 62.200 243.600 69.600 ;
        RECT 244.600 67.400 245.200 70.400 ;
        RECT 249.200 68.300 250.000 79.800 ;
        RECT 253.400 72.400 254.200 79.800 ;
        RECT 254.800 73.600 255.600 74.400 ;
        RECT 255.000 72.400 255.600 73.600 ;
        RECT 258.000 73.600 258.800 74.400 ;
        RECT 258.000 72.400 258.600 73.600 ;
        RECT 259.400 72.400 260.200 79.800 ;
        RECT 253.400 71.800 254.400 72.400 ;
        RECT 255.000 71.800 256.400 72.400 ;
        RECT 252.400 68.800 253.200 70.400 ;
        RECT 253.800 68.400 254.400 71.800 ;
        RECT 255.600 71.600 256.400 71.800 ;
        RECT 257.200 71.800 258.600 72.400 ;
        RECT 259.200 71.800 260.200 72.400 ;
        RECT 257.200 71.600 258.000 71.800 ;
        RECT 255.700 70.300 256.300 71.600 ;
        RECT 259.200 70.300 259.800 71.800 ;
        RECT 255.700 69.700 259.800 70.300 ;
        RECT 259.200 68.400 259.800 69.700 ;
        RECT 265.200 70.300 266.000 79.800 ;
        RECT 274.800 72.000 275.600 79.800 ;
        RECT 278.000 75.200 278.800 79.800 ;
        RECT 274.600 71.200 275.600 72.000 ;
        RECT 276.200 74.600 278.800 75.200 ;
        RECT 276.200 73.000 276.800 74.600 ;
        RECT 281.200 74.400 282.000 79.800 ;
        RECT 284.400 77.000 285.200 79.800 ;
        RECT 286.000 77.000 286.800 79.800 ;
        RECT 287.600 77.000 288.400 79.800 ;
        RECT 282.600 74.400 286.800 75.200 ;
        RECT 279.400 73.600 282.000 74.400 ;
        RECT 289.200 73.600 290.000 79.800 ;
        RECT 292.400 75.000 293.200 79.800 ;
        RECT 295.600 75.000 296.400 79.800 ;
        RECT 297.200 77.000 298.000 79.800 ;
        RECT 298.800 77.000 299.600 79.800 ;
        RECT 302.000 75.200 302.800 79.800 ;
        RECT 305.200 76.400 306.000 79.800 ;
        RECT 305.200 75.800 306.200 76.400 ;
        RECT 305.600 75.200 306.200 75.800 ;
        RECT 300.800 74.400 305.000 75.200 ;
        RECT 305.600 74.600 307.600 75.200 ;
        RECT 292.400 73.600 295.000 74.400 ;
        RECT 295.600 73.800 301.400 74.400 ;
        RECT 304.400 74.000 305.000 74.400 ;
        RECT 284.400 73.000 285.200 73.200 ;
        RECT 276.200 72.400 285.200 73.000 ;
        RECT 287.600 73.000 288.400 73.200 ;
        RECT 295.600 73.000 296.200 73.800 ;
        RECT 302.000 73.200 303.400 73.800 ;
        RECT 304.400 73.200 306.000 74.000 ;
        RECT 287.600 72.400 296.200 73.000 ;
        RECT 297.200 73.000 303.400 73.200 ;
        RECT 297.200 72.600 302.600 73.000 ;
        RECT 297.200 72.400 298.000 72.600 ;
        RECT 273.200 70.300 274.000 70.400 ;
        RECT 265.200 69.700 274.000 70.300 ;
        RECT 250.800 68.300 251.600 68.400 ;
        RECT 249.200 68.200 251.600 68.300 ;
        RECT 249.200 67.700 252.400 68.200 ;
        RECT 244.600 66.800 246.800 67.400 ;
        RECT 246.000 62.200 246.800 66.800 ;
        RECT 247.600 64.800 248.400 66.400 ;
        RECT 249.200 62.200 250.000 67.700 ;
        RECT 250.800 67.600 252.400 67.700 ;
        RECT 253.800 67.600 256.400 68.400 ;
        RECT 257.200 67.600 259.800 68.400 ;
        RECT 262.000 68.200 262.800 68.400 ;
        RECT 261.200 67.600 262.800 68.200 ;
        RECT 251.600 67.200 252.400 67.600 ;
        RECT 251.000 66.200 254.600 66.600 ;
        RECT 255.600 66.200 256.200 67.600 ;
        RECT 257.400 66.200 258.000 67.600 ;
        RECT 261.200 67.200 262.000 67.600 ;
        RECT 259.000 66.200 262.600 66.600 ;
        RECT 250.800 66.000 254.800 66.200 ;
        RECT 250.800 62.200 251.600 66.000 ;
        RECT 254.000 62.200 254.800 66.000 ;
        RECT 255.600 62.200 256.400 66.200 ;
        RECT 257.200 62.200 258.000 66.200 ;
        RECT 258.800 66.000 262.800 66.200 ;
        RECT 258.800 62.200 259.600 66.000 ;
        RECT 262.000 62.200 262.800 66.000 ;
        RECT 263.600 64.800 264.400 66.400 ;
        RECT 265.200 62.200 266.000 69.700 ;
        RECT 273.200 69.600 274.000 69.700 ;
        RECT 274.600 66.800 275.400 71.200 ;
        RECT 276.200 70.600 276.800 72.400 ;
        RECT 300.200 71.800 301.000 72.000 ;
        RECT 303.600 71.800 304.400 72.400 ;
        RECT 277.400 71.200 304.400 71.800 ;
        RECT 277.400 71.000 278.200 71.200 ;
        RECT 276.000 70.000 276.800 70.600 ;
        RECT 276.000 68.000 276.600 70.000 ;
        RECT 277.200 68.600 281.000 69.400 ;
        RECT 276.000 67.400 277.200 68.000 ;
        RECT 266.800 66.300 267.600 66.400 ;
        RECT 274.600 66.300 275.600 66.800 ;
        RECT 266.800 65.700 275.600 66.300 ;
        RECT 266.800 65.600 267.600 65.700 ;
        RECT 274.800 62.200 275.600 65.700 ;
        RECT 276.400 62.200 277.200 67.400 ;
        RECT 280.200 67.400 281.000 68.600 ;
        RECT 280.200 66.800 282.000 67.400 ;
        RECT 281.200 66.200 282.000 66.800 ;
        RECT 286.000 66.400 286.800 69.200 ;
        RECT 289.200 68.600 292.400 69.400 ;
        RECT 296.200 68.600 298.200 69.400 ;
        RECT 306.800 69.000 307.600 74.600 ;
        RECT 311.000 72.400 311.800 79.800 ;
        RECT 312.400 73.600 313.200 74.400 ;
        RECT 312.600 72.400 313.200 73.600 ;
        RECT 315.600 73.600 316.400 74.400 ;
        RECT 315.600 72.400 316.200 73.600 ;
        RECT 317.000 72.400 317.800 79.800 ;
        RECT 311.000 71.800 312.000 72.400 ;
        RECT 312.600 71.800 314.000 72.400 ;
        RECT 288.800 67.800 289.600 68.000 ;
        RECT 288.800 67.200 293.200 67.800 ;
        RECT 292.400 67.000 293.200 67.200 ;
        RECT 294.000 66.800 294.800 68.400 ;
        RECT 281.200 65.400 283.600 66.200 ;
        RECT 286.000 65.600 287.000 66.400 ;
        RECT 290.000 65.600 291.600 66.400 ;
        RECT 292.400 66.200 293.200 66.400 ;
        RECT 296.200 66.200 297.000 68.600 ;
        RECT 298.800 68.200 307.600 69.000 ;
        RECT 310.000 68.800 310.800 70.400 ;
        RECT 311.400 68.400 312.000 71.800 ;
        RECT 313.200 71.600 314.000 71.800 ;
        RECT 314.800 71.800 316.200 72.400 ;
        RECT 316.800 71.800 317.800 72.400 ;
        RECT 321.200 72.400 322.000 79.800 ;
        RECT 321.200 71.800 323.400 72.400 ;
        RECT 324.400 71.800 325.200 79.800 ;
        RECT 328.600 71.800 330.600 79.800 ;
        RECT 314.800 71.600 315.600 71.800 ;
        RECT 313.300 70.300 313.900 71.600 ;
        RECT 316.800 70.300 317.400 71.800 ;
        RECT 313.300 69.700 317.400 70.300 ;
        RECT 316.800 68.400 317.400 69.700 ;
        RECT 322.800 71.200 323.400 71.800 ;
        RECT 322.800 70.400 324.000 71.200 ;
        RECT 302.200 66.800 305.200 67.600 ;
        RECT 302.200 66.200 303.000 66.800 ;
        RECT 292.400 65.600 297.000 66.200 ;
        RECT 282.800 62.200 283.600 65.400 ;
        RECT 300.400 65.400 303.000 66.200 ;
        RECT 284.400 62.200 285.200 65.000 ;
        RECT 286.000 62.200 286.800 65.000 ;
        RECT 287.600 62.200 288.400 65.000 ;
        RECT 289.200 62.200 290.000 65.000 ;
        RECT 292.400 62.200 293.200 65.000 ;
        RECT 295.600 62.200 296.400 65.000 ;
        RECT 297.200 62.200 298.000 65.000 ;
        RECT 298.800 62.200 299.600 65.000 ;
        RECT 300.400 62.200 301.200 65.400 ;
        RECT 306.800 62.200 307.600 68.200 ;
        RECT 308.400 68.200 309.200 68.400 ;
        RECT 308.400 67.600 310.000 68.200 ;
        RECT 311.400 67.600 314.000 68.400 ;
        RECT 314.800 67.600 317.400 68.400 ;
        RECT 319.600 68.200 320.400 68.400 ;
        RECT 318.800 67.600 320.400 68.200 ;
        RECT 309.200 67.200 310.000 67.600 ;
        RECT 308.600 66.200 312.200 66.600 ;
        RECT 313.200 66.200 313.800 67.600 ;
        RECT 315.000 66.200 315.600 67.600 ;
        RECT 318.800 67.200 319.600 67.600 ;
        RECT 322.800 67.400 323.400 70.400 ;
        RECT 324.600 69.600 325.200 71.800 ;
        RECT 321.200 66.800 323.400 67.400 ;
        RECT 316.600 66.200 320.200 66.600 ;
        RECT 308.400 66.000 312.400 66.200 ;
        RECT 308.400 62.200 309.200 66.000 ;
        RECT 311.600 62.200 312.400 66.000 ;
        RECT 313.200 62.200 314.000 66.200 ;
        RECT 314.800 62.200 315.600 66.200 ;
        RECT 316.400 66.000 320.400 66.200 ;
        RECT 316.400 62.200 317.200 66.000 ;
        RECT 319.600 62.200 320.400 66.000 ;
        RECT 321.200 62.200 322.000 66.800 ;
        RECT 324.400 62.200 325.200 69.600 ;
        RECT 326.000 67.600 326.800 69.200 ;
        RECT 327.600 68.800 328.400 70.400 ;
        RECT 329.400 68.400 330.000 71.800 ;
        RECT 330.800 68.800 331.600 70.400 ;
        RECT 329.200 68.200 330.000 68.400 ;
        RECT 332.400 68.300 333.200 68.400 ;
        RECT 334.000 68.300 334.800 79.800 ;
        RECT 338.800 72.000 339.600 79.800 ;
        RECT 342.000 75.200 342.800 79.800 ;
        RECT 332.400 68.200 334.800 68.300 ;
        RECT 327.600 67.600 330.000 68.200 ;
        RECT 331.600 67.700 334.800 68.200 ;
        RECT 331.600 67.600 333.200 67.700 ;
        RECT 327.600 66.200 328.200 67.600 ;
        RECT 331.600 67.200 332.400 67.600 ;
        RECT 329.400 66.200 333.000 66.600 ;
        RECT 326.000 62.800 326.800 66.200 ;
        RECT 327.600 63.400 328.400 66.200 ;
        RECT 329.200 66.000 333.200 66.200 ;
        RECT 329.200 62.800 330.000 66.000 ;
        RECT 326.000 62.200 330.000 62.800 ;
        RECT 332.400 62.200 333.200 66.000 ;
        RECT 334.000 62.200 334.800 67.700 ;
        RECT 338.600 71.200 339.600 72.000 ;
        RECT 340.200 74.600 342.800 75.200 ;
        RECT 340.200 73.000 340.800 74.600 ;
        RECT 345.200 74.400 346.000 79.800 ;
        RECT 348.400 77.000 349.200 79.800 ;
        RECT 350.000 77.000 350.800 79.800 ;
        RECT 351.600 77.000 352.400 79.800 ;
        RECT 346.600 74.400 350.800 75.200 ;
        RECT 343.400 73.600 346.000 74.400 ;
        RECT 353.200 73.600 354.000 79.800 ;
        RECT 356.400 75.000 357.200 79.800 ;
        RECT 359.600 75.000 360.400 79.800 ;
        RECT 361.200 77.000 362.000 79.800 ;
        RECT 362.800 77.000 363.600 79.800 ;
        RECT 366.000 75.200 366.800 79.800 ;
        RECT 369.200 76.400 370.000 79.800 ;
        RECT 369.200 75.800 370.200 76.400 ;
        RECT 369.600 75.200 370.200 75.800 ;
        RECT 364.800 74.400 369.000 75.200 ;
        RECT 369.600 74.600 371.600 75.200 ;
        RECT 356.400 73.600 359.000 74.400 ;
        RECT 359.600 73.800 365.400 74.400 ;
        RECT 368.400 74.000 369.000 74.400 ;
        RECT 348.400 73.000 349.200 73.200 ;
        RECT 340.200 72.400 349.200 73.000 ;
        RECT 351.600 73.000 352.400 73.200 ;
        RECT 359.600 73.000 360.200 73.800 ;
        RECT 366.000 73.200 367.400 73.800 ;
        RECT 368.400 73.200 370.000 74.000 ;
        RECT 351.600 72.400 360.200 73.000 ;
        RECT 361.200 73.000 367.400 73.200 ;
        RECT 361.200 72.600 366.600 73.000 ;
        RECT 361.200 72.400 362.000 72.600 ;
        RECT 338.600 66.800 339.400 71.200 ;
        RECT 340.200 70.600 340.800 72.400 ;
        RECT 340.000 70.000 340.800 70.600 ;
        RECT 346.800 70.000 370.200 70.600 ;
        RECT 340.000 68.000 340.600 70.000 ;
        RECT 346.800 69.400 347.600 70.000 ;
        RECT 364.400 69.600 365.200 70.000 ;
        RECT 367.600 69.600 368.400 70.000 ;
        RECT 369.400 69.800 370.200 70.000 ;
        RECT 341.200 68.600 345.000 69.400 ;
        RECT 340.000 67.400 341.200 68.000 ;
        RECT 335.600 66.300 336.400 66.400 ;
        RECT 338.600 66.300 339.600 66.800 ;
        RECT 335.600 65.700 339.600 66.300 ;
        RECT 335.600 64.800 336.400 65.700 ;
        RECT 338.800 62.200 339.600 65.700 ;
        RECT 340.400 62.200 341.200 67.400 ;
        RECT 344.200 67.400 345.000 68.600 ;
        RECT 344.200 66.800 346.000 67.400 ;
        RECT 345.200 66.200 346.000 66.800 ;
        RECT 350.000 66.400 350.800 69.200 ;
        RECT 353.200 68.600 356.400 69.400 ;
        RECT 360.200 68.600 362.200 69.400 ;
        RECT 370.800 69.000 371.600 74.600 ;
        RECT 375.000 72.400 375.800 79.800 ;
        RECT 376.400 73.600 377.200 74.400 ;
        RECT 376.600 72.400 377.200 73.600 ;
        RECT 375.000 71.800 376.000 72.400 ;
        RECT 376.600 71.800 378.000 72.400 ;
        RECT 381.400 71.800 383.400 79.800 ;
        RECT 389.400 72.400 390.200 79.800 ;
        RECT 390.800 73.600 391.600 74.400 ;
        RECT 391.000 72.400 391.600 73.600 ;
        RECT 389.400 71.800 390.400 72.400 ;
        RECT 391.000 71.800 392.400 72.400 ;
        RECT 375.400 70.400 376.000 71.800 ;
        RECT 377.200 71.600 378.000 71.800 ;
        RECT 352.800 67.800 353.600 68.000 ;
        RECT 352.800 67.200 357.200 67.800 ;
        RECT 356.400 67.000 357.200 67.200 ;
        RECT 358.000 66.800 358.800 68.400 ;
        RECT 345.200 65.400 347.600 66.200 ;
        RECT 350.000 65.600 351.000 66.400 ;
        RECT 354.000 65.600 355.600 66.400 ;
        RECT 356.400 66.200 357.200 66.400 ;
        RECT 360.200 66.200 361.000 68.600 ;
        RECT 362.800 68.200 371.600 69.000 ;
        RECT 374.000 68.800 374.800 70.400 ;
        RECT 375.400 69.600 376.400 70.400 ;
        RECT 375.400 68.400 376.000 69.600 ;
        RECT 366.200 66.800 369.200 67.600 ;
        RECT 366.200 66.200 367.000 66.800 ;
        RECT 356.400 65.600 361.000 66.200 ;
        RECT 346.800 62.200 347.600 65.400 ;
        RECT 364.400 65.400 367.000 66.200 ;
        RECT 348.400 62.200 349.200 65.000 ;
        RECT 350.000 62.200 350.800 65.000 ;
        RECT 351.600 62.200 352.400 65.000 ;
        RECT 353.200 62.200 354.000 65.000 ;
        RECT 356.400 62.200 357.200 65.000 ;
        RECT 359.600 62.200 360.400 65.000 ;
        RECT 361.200 62.200 362.000 65.000 ;
        RECT 362.800 62.200 363.600 65.000 ;
        RECT 364.400 62.200 365.200 65.400 ;
        RECT 370.800 62.200 371.600 68.200 ;
        RECT 372.400 68.200 373.200 68.400 ;
        RECT 372.400 67.600 374.000 68.200 ;
        RECT 375.400 67.600 378.000 68.400 ;
        RECT 378.800 67.600 379.600 69.200 ;
        RECT 380.400 68.800 381.200 70.400 ;
        RECT 382.200 68.400 382.800 71.800 ;
        RECT 383.600 70.300 384.400 70.400 ;
        RECT 385.200 70.300 386.000 70.400 ;
        RECT 383.600 69.700 386.000 70.300 ;
        RECT 383.600 68.800 384.400 69.700 ;
        RECT 385.200 69.600 386.000 69.700 ;
        RECT 388.400 68.800 389.200 70.400 ;
        RECT 389.800 68.400 390.400 71.800 ;
        RECT 391.600 71.600 392.400 71.800 ;
        RECT 382.000 68.200 382.800 68.400 ;
        RECT 385.200 68.300 386.000 68.400 ;
        RECT 386.800 68.300 387.600 68.400 ;
        RECT 385.200 68.200 387.600 68.300 ;
        RECT 380.400 67.600 382.800 68.200 ;
        RECT 384.400 67.700 388.400 68.200 ;
        RECT 384.400 67.600 386.000 67.700 ;
        RECT 386.800 67.600 388.400 67.700 ;
        RECT 389.800 67.600 392.400 68.400 ;
        RECT 373.200 67.200 374.000 67.600 ;
        RECT 372.600 66.200 376.200 66.600 ;
        RECT 377.200 66.200 377.800 67.600 ;
        RECT 380.400 66.200 381.000 67.600 ;
        RECT 384.400 67.200 385.200 67.600 ;
        RECT 387.600 67.200 388.400 67.600 ;
        RECT 382.200 66.200 385.800 66.600 ;
        RECT 387.000 66.200 390.600 66.600 ;
        RECT 391.600 66.200 392.200 67.600 ;
        RECT 372.400 66.000 376.400 66.200 ;
        RECT 372.400 62.200 373.200 66.000 ;
        RECT 375.600 62.200 376.400 66.000 ;
        RECT 377.200 62.200 378.000 66.200 ;
        RECT 378.800 62.800 379.600 66.200 ;
        RECT 380.400 63.400 381.200 66.200 ;
        RECT 382.000 66.000 386.000 66.200 ;
        RECT 382.000 62.800 382.800 66.000 ;
        RECT 378.800 62.200 382.800 62.800 ;
        RECT 385.200 62.200 386.000 66.000 ;
        RECT 386.800 66.000 390.800 66.200 ;
        RECT 386.800 62.200 387.600 66.000 ;
        RECT 390.000 62.200 390.800 66.000 ;
        RECT 391.600 62.200 392.400 66.200 ;
        RECT 393.200 62.200 394.000 79.800 ;
        RECT 394.800 72.300 395.600 72.400 ;
        RECT 396.400 72.300 397.200 73.200 ;
        RECT 394.800 71.700 397.200 72.300 ;
        RECT 394.800 71.600 395.600 71.700 ;
        RECT 396.400 71.600 397.200 71.700 ;
        RECT 394.800 64.800 395.600 66.400 ;
        RECT 398.000 66.200 398.800 79.800 ;
        RECT 401.800 72.600 402.600 79.800 ;
        RECT 407.600 78.300 408.400 79.800 ;
        RECT 410.800 78.300 411.600 78.400 ;
        RECT 407.600 77.700 411.600 78.300 ;
        RECT 401.800 71.800 403.600 72.600 ;
        RECT 401.200 69.600 402.000 71.200 ;
        RECT 402.800 68.400 403.400 71.800 ;
        RECT 399.600 66.800 400.400 68.400 ;
        RECT 402.800 67.600 403.600 68.400 ;
        RECT 397.000 65.600 398.800 66.200 ;
        RECT 397.000 62.200 397.800 65.600 ;
        RECT 402.800 64.400 403.400 67.600 ;
        RECT 404.400 64.800 405.200 66.400 ;
        RECT 406.000 64.800 406.800 66.400 ;
        RECT 402.800 62.200 403.600 64.400 ;
        RECT 407.600 62.200 408.400 77.700 ;
        RECT 410.800 77.600 411.600 77.700 ;
        RECT 417.200 72.000 418.000 79.800 ;
        RECT 420.400 75.200 421.200 79.800 ;
        RECT 417.000 71.200 418.000 72.000 ;
        RECT 418.600 74.600 421.200 75.200 ;
        RECT 418.600 73.000 419.200 74.600 ;
        RECT 423.600 74.400 424.400 79.800 ;
        RECT 426.800 77.000 427.600 79.800 ;
        RECT 428.400 77.000 429.200 79.800 ;
        RECT 430.000 77.000 430.800 79.800 ;
        RECT 425.000 74.400 429.200 75.200 ;
        RECT 421.800 73.600 424.400 74.400 ;
        RECT 431.600 73.600 432.400 79.800 ;
        RECT 434.800 75.000 435.600 79.800 ;
        RECT 438.000 75.000 438.800 79.800 ;
        RECT 439.600 77.000 440.400 79.800 ;
        RECT 441.200 77.000 442.000 79.800 ;
        RECT 444.400 75.200 445.200 79.800 ;
        RECT 447.600 76.400 448.400 79.800 ;
        RECT 447.600 75.800 448.600 76.400 ;
        RECT 448.000 75.200 448.600 75.800 ;
        RECT 443.200 74.400 447.400 75.200 ;
        RECT 448.000 74.600 450.000 75.200 ;
        RECT 434.800 73.600 437.400 74.400 ;
        RECT 438.000 73.800 443.800 74.400 ;
        RECT 446.800 74.000 447.400 74.400 ;
        RECT 426.800 73.000 427.600 73.200 ;
        RECT 418.600 72.400 427.600 73.000 ;
        RECT 430.000 73.000 430.800 73.200 ;
        RECT 438.000 73.000 438.600 73.800 ;
        RECT 444.400 73.200 445.800 73.800 ;
        RECT 446.800 73.200 448.400 74.000 ;
        RECT 430.000 72.400 438.600 73.000 ;
        RECT 439.600 73.000 445.800 73.200 ;
        RECT 439.600 72.600 445.000 73.000 ;
        RECT 439.600 72.400 440.400 72.600 ;
        RECT 417.000 66.800 417.800 71.200 ;
        RECT 418.600 70.600 419.200 72.400 ;
        RECT 418.400 70.000 419.200 70.600 ;
        RECT 425.200 70.000 448.600 70.600 ;
        RECT 418.400 68.000 419.000 70.000 ;
        RECT 425.200 69.400 426.000 70.000 ;
        RECT 442.800 69.600 443.600 70.000 ;
        RECT 446.000 69.600 446.800 70.000 ;
        RECT 447.800 69.800 448.600 70.000 ;
        RECT 419.600 68.600 423.400 69.400 ;
        RECT 418.400 67.400 419.600 68.000 ;
        RECT 417.000 66.000 418.000 66.800 ;
        RECT 417.200 62.200 418.000 66.000 ;
        RECT 418.800 62.200 419.600 67.400 ;
        RECT 422.600 67.400 423.400 68.600 ;
        RECT 422.600 66.800 424.400 67.400 ;
        RECT 423.600 66.200 424.400 66.800 ;
        RECT 428.400 66.400 429.200 69.200 ;
        RECT 431.600 68.600 434.800 69.400 ;
        RECT 438.600 68.600 440.600 69.400 ;
        RECT 449.200 69.000 450.000 74.600 ;
        RECT 451.600 73.600 452.400 74.400 ;
        RECT 451.600 72.400 452.200 73.600 ;
        RECT 453.000 72.400 453.800 79.800 ;
        RECT 450.800 71.800 452.200 72.400 ;
        RECT 452.800 71.800 453.800 72.400 ;
        RECT 450.800 71.600 451.600 71.800 ;
        RECT 431.200 67.800 432.000 68.000 ;
        RECT 431.200 67.200 435.600 67.800 ;
        RECT 434.800 67.000 435.600 67.200 ;
        RECT 436.400 66.800 437.200 68.400 ;
        RECT 423.600 65.400 426.000 66.200 ;
        RECT 428.400 65.600 429.400 66.400 ;
        RECT 432.400 65.600 434.000 66.400 ;
        RECT 434.800 66.200 435.600 66.400 ;
        RECT 438.600 66.200 439.400 68.600 ;
        RECT 441.200 68.200 450.000 69.000 ;
        RECT 452.800 68.400 453.400 71.800 ;
        RECT 454.000 70.300 454.800 70.400 ;
        RECT 455.600 70.300 456.400 70.400 ;
        RECT 454.000 69.700 456.400 70.300 ;
        RECT 454.000 68.800 454.800 69.700 ;
        RECT 455.600 69.600 456.400 69.700 ;
        RECT 444.600 66.800 447.600 67.600 ;
        RECT 444.600 66.200 445.400 66.800 ;
        RECT 434.800 65.600 439.400 66.200 ;
        RECT 425.200 62.200 426.000 65.400 ;
        RECT 442.800 65.400 445.400 66.200 ;
        RECT 426.800 62.200 427.600 65.000 ;
        RECT 428.400 62.200 429.200 65.000 ;
        RECT 430.000 62.200 430.800 65.000 ;
        RECT 431.600 62.200 432.400 65.000 ;
        RECT 434.800 62.200 435.600 65.000 ;
        RECT 438.000 62.200 438.800 65.000 ;
        RECT 439.600 62.200 440.400 65.000 ;
        RECT 441.200 62.200 442.000 65.000 ;
        RECT 442.800 62.200 443.600 65.400 ;
        RECT 449.200 62.200 450.000 68.200 ;
        RECT 450.800 67.600 453.400 68.400 ;
        RECT 455.600 68.300 456.400 68.400 ;
        RECT 457.200 68.300 458.000 79.800 ;
        RECT 460.400 71.800 461.200 79.800 ;
        RECT 462.000 72.400 462.800 79.800 ;
        RECT 465.200 72.400 466.000 79.800 ;
        RECT 462.000 71.800 466.000 72.400 ;
        RECT 460.600 70.400 461.200 71.800 ;
        RECT 466.800 71.600 467.600 73.200 ;
        RECT 464.400 70.400 465.200 70.800 ;
        RECT 460.400 69.800 462.800 70.400 ;
        RECT 464.400 70.300 466.000 70.400 ;
        RECT 466.800 70.300 467.600 70.400 ;
        RECT 464.400 69.800 467.600 70.300 ;
        RECT 460.400 69.600 461.200 69.800 ;
        RECT 455.600 68.200 458.000 68.300 ;
        RECT 454.800 67.700 458.000 68.200 ;
        RECT 454.800 67.600 456.400 67.700 ;
        RECT 451.000 66.200 451.600 67.600 ;
        RECT 454.800 67.200 455.600 67.600 ;
        RECT 452.600 66.200 456.200 66.600 ;
        RECT 450.800 62.200 451.600 66.200 ;
        RECT 452.400 66.000 456.400 66.200 ;
        RECT 452.400 62.200 453.200 66.000 ;
        RECT 455.600 62.200 456.400 66.000 ;
        RECT 457.200 62.200 458.000 67.700 ;
        RECT 458.800 68.300 459.600 68.400 ;
        RECT 462.200 68.300 462.800 69.800 ;
        RECT 465.200 69.700 467.600 69.800 ;
        RECT 465.200 69.600 466.000 69.700 ;
        RECT 466.800 69.600 467.600 69.700 ;
        RECT 458.800 67.700 462.800 68.300 ;
        RECT 458.800 67.600 459.600 67.700 ;
        RECT 458.800 64.800 459.600 66.400 ;
        RECT 460.400 65.600 461.200 66.400 ;
        RECT 462.200 66.200 462.800 67.700 ;
        RECT 463.600 68.300 464.400 69.200 ;
        RECT 465.200 68.300 466.000 68.400 ;
        RECT 463.600 67.700 466.000 68.300 ;
        RECT 463.600 67.600 464.400 67.700 ;
        RECT 465.200 67.600 466.000 67.700 ;
        RECT 468.400 66.200 469.200 79.800 ;
        RECT 471.600 71.800 472.400 79.800 ;
        RECT 473.200 72.400 474.000 79.800 ;
        RECT 476.400 72.400 477.200 79.800 ;
        RECT 481.800 72.800 482.600 79.800 ;
        RECT 486.000 75.000 486.800 79.000 ;
        RECT 473.200 71.800 477.200 72.400 ;
        RECT 481.000 72.200 482.600 72.800 ;
        RECT 471.800 70.400 472.400 71.800 ;
        RECT 475.600 70.400 476.400 70.800 ;
        RECT 471.600 69.800 474.000 70.400 ;
        RECT 475.600 69.800 477.200 70.400 ;
        RECT 471.600 69.600 472.400 69.800 ;
        RECT 470.000 68.300 470.800 68.400 ;
        RECT 473.400 68.300 474.000 69.800 ;
        RECT 476.400 69.600 477.200 69.800 ;
        RECT 478.000 70.300 478.800 70.400 ;
        RECT 479.600 70.300 480.400 71.200 ;
        RECT 478.000 69.700 480.400 70.300 ;
        RECT 478.000 69.600 478.800 69.700 ;
        RECT 479.600 69.600 480.400 69.700 ;
        RECT 470.000 67.700 474.000 68.300 ;
        RECT 470.000 66.800 470.800 67.700 ;
        RECT 460.600 64.800 461.400 65.600 ;
        RECT 462.000 62.200 462.800 66.200 ;
        RECT 467.400 65.600 469.200 66.200 ;
        RECT 471.600 65.600 472.400 66.400 ;
        RECT 473.400 66.200 474.000 67.700 ;
        RECT 474.800 67.600 475.600 69.200 ;
        RECT 481.000 68.400 481.600 72.200 ;
        RECT 486.200 71.600 486.800 75.000 ;
        RECT 483.000 71.000 486.800 71.600 ;
        RECT 483.000 69.000 483.600 71.000 ;
        RECT 479.600 67.600 481.600 68.400 ;
        RECT 482.200 68.200 483.600 69.000 ;
        RECT 484.400 68.800 485.200 70.400 ;
        RECT 486.000 70.300 486.800 70.400 ;
        RECT 487.600 70.300 488.400 70.400 ;
        RECT 486.000 69.700 488.400 70.300 ;
        RECT 486.000 68.800 486.800 69.700 ;
        RECT 487.600 69.600 488.400 69.700 ;
        RECT 489.200 70.300 490.000 79.800 ;
        RECT 490.800 71.600 491.600 73.200 ;
        RECT 495.000 72.400 495.800 79.800 ;
        RECT 501.000 78.400 501.800 79.800 ;
        RECT 501.000 77.600 502.800 78.400 ;
        RECT 496.400 73.600 497.200 74.400 ;
        RECT 496.600 72.400 497.200 73.600 ;
        RECT 499.600 73.600 500.400 74.400 ;
        RECT 499.600 72.400 500.200 73.600 ;
        RECT 501.000 72.400 501.800 77.600 ;
        RECT 495.000 71.800 496.000 72.400 ;
        RECT 496.600 71.800 498.000 72.400 ;
        RECT 492.400 70.300 493.200 70.400 ;
        RECT 489.200 69.700 493.200 70.300 ;
        RECT 467.400 62.200 468.200 65.600 ;
        RECT 471.800 64.800 472.600 65.600 ;
        RECT 473.200 62.200 474.000 66.200 ;
        RECT 481.000 67.000 481.600 67.600 ;
        RECT 482.600 67.800 483.600 68.200 ;
        RECT 482.600 67.200 486.800 67.800 ;
        RECT 481.000 66.600 481.800 67.000 ;
        RECT 481.000 66.400 482.600 66.600 ;
        RECT 481.000 66.000 483.600 66.400 ;
        RECT 481.800 65.600 483.600 66.000 ;
        RECT 481.800 63.000 482.600 65.600 ;
        RECT 486.200 65.000 486.800 67.200 ;
        RECT 487.600 66.800 488.400 68.400 ;
        RECT 489.200 66.200 490.000 69.700 ;
        RECT 492.400 69.600 493.200 69.700 ;
        RECT 494.000 68.800 494.800 70.400 ;
        RECT 495.400 68.400 496.000 71.800 ;
        RECT 497.200 71.600 498.000 71.800 ;
        RECT 498.800 71.800 500.200 72.400 ;
        RECT 500.800 71.800 501.800 72.400 ;
        RECT 498.800 71.600 499.600 71.800 ;
        RECT 500.800 68.400 501.400 71.800 ;
        RECT 505.200 71.600 506.000 73.200 ;
        RECT 502.000 68.800 502.800 70.400 ;
        RECT 490.800 68.300 491.600 68.400 ;
        RECT 492.400 68.300 493.200 68.400 ;
        RECT 490.800 68.200 493.200 68.300 ;
        RECT 490.800 67.700 494.000 68.200 ;
        RECT 490.800 67.600 491.600 67.700 ;
        RECT 492.400 67.600 494.000 67.700 ;
        RECT 495.400 67.600 498.000 68.400 ;
        RECT 498.800 67.600 501.400 68.400 ;
        RECT 503.600 68.200 504.400 68.400 ;
        RECT 502.800 67.600 504.400 68.200 ;
        RECT 493.200 67.200 494.000 67.600 ;
        RECT 492.600 66.200 496.200 66.600 ;
        RECT 497.200 66.200 497.800 67.600 ;
        RECT 499.000 66.200 499.600 67.600 ;
        RECT 502.800 67.200 503.600 67.600 ;
        RECT 500.600 66.200 504.200 66.600 ;
        RECT 506.800 66.200 507.600 79.800 ;
        RECT 508.400 72.300 509.200 72.400 ;
        RECT 510.000 72.300 510.800 73.200 ;
        RECT 508.400 71.700 510.800 72.300 ;
        RECT 508.400 71.600 509.200 71.700 ;
        RECT 510.000 71.600 510.800 71.700 ;
        RECT 508.400 68.300 509.200 68.400 ;
        RECT 510.000 68.300 510.800 68.400 ;
        RECT 508.400 67.700 510.800 68.300 ;
        RECT 508.400 66.800 509.200 67.700 ;
        RECT 510.000 67.600 510.800 67.700 ;
        RECT 511.600 66.200 512.400 79.800 ;
        RECT 516.400 72.000 517.200 79.800 ;
        RECT 519.600 75.200 520.400 79.800 ;
        RECT 516.200 71.200 517.200 72.000 ;
        RECT 517.800 74.600 520.400 75.200 ;
        RECT 517.800 73.000 518.400 74.600 ;
        RECT 522.800 74.400 523.600 79.800 ;
        RECT 526.000 77.000 526.800 79.800 ;
        RECT 527.600 77.000 528.400 79.800 ;
        RECT 529.200 77.000 530.000 79.800 ;
        RECT 524.200 74.400 528.400 75.200 ;
        RECT 521.000 73.600 523.600 74.400 ;
        RECT 530.800 73.600 531.600 79.800 ;
        RECT 534.000 75.000 534.800 79.800 ;
        RECT 537.200 75.000 538.000 79.800 ;
        RECT 538.800 77.000 539.600 79.800 ;
        RECT 540.400 77.000 541.200 79.800 ;
        RECT 543.600 75.200 544.400 79.800 ;
        RECT 546.800 76.400 547.600 79.800 ;
        RECT 546.800 75.800 547.800 76.400 ;
        RECT 547.200 75.200 547.800 75.800 ;
        RECT 542.400 74.400 546.600 75.200 ;
        RECT 547.200 74.600 549.200 75.200 ;
        RECT 534.000 73.600 536.600 74.400 ;
        RECT 537.200 73.800 543.000 74.400 ;
        RECT 546.000 74.000 546.600 74.400 ;
        RECT 526.000 73.000 526.800 73.200 ;
        RECT 517.800 72.400 526.800 73.000 ;
        RECT 529.200 73.000 530.000 73.200 ;
        RECT 537.200 73.000 537.800 73.800 ;
        RECT 543.600 73.200 545.000 73.800 ;
        RECT 546.000 73.200 547.600 74.000 ;
        RECT 529.200 72.400 537.800 73.000 ;
        RECT 538.800 73.000 545.000 73.200 ;
        RECT 538.800 72.600 544.200 73.000 ;
        RECT 538.800 72.400 539.600 72.600 ;
        RECT 513.200 68.300 514.000 68.400 ;
        RECT 514.800 68.300 515.600 68.400 ;
        RECT 513.200 67.700 515.600 68.300 ;
        RECT 513.200 66.800 514.000 67.700 ;
        RECT 514.800 67.600 515.600 67.700 ;
        RECT 516.200 66.800 517.000 71.200 ;
        RECT 517.800 70.600 518.400 72.400 ;
        RECT 517.600 70.000 518.400 70.600 ;
        RECT 524.400 70.000 547.800 70.600 ;
        RECT 517.600 68.000 518.200 70.000 ;
        RECT 524.400 69.400 525.200 70.000 ;
        RECT 542.000 69.600 542.800 70.000 ;
        RECT 547.000 69.800 547.800 70.000 ;
        RECT 518.800 68.600 522.600 69.400 ;
        RECT 517.600 67.400 518.800 68.000 ;
        RECT 489.200 65.600 491.000 66.200 ;
        RECT 486.000 63.000 486.800 65.000 ;
        RECT 490.200 62.200 491.000 65.600 ;
        RECT 492.400 66.000 496.400 66.200 ;
        RECT 492.400 62.200 493.200 66.000 ;
        RECT 495.600 62.200 496.400 66.000 ;
        RECT 497.200 62.200 498.000 66.200 ;
        RECT 498.800 62.200 499.600 66.200 ;
        RECT 500.400 66.000 504.400 66.200 ;
        RECT 500.400 62.200 501.200 66.000 ;
        RECT 503.600 62.200 504.400 66.000 ;
        RECT 505.800 65.600 507.600 66.200 ;
        RECT 510.600 65.600 512.400 66.200 ;
        RECT 516.200 66.000 517.200 66.800 ;
        RECT 505.800 64.400 506.600 65.600 ;
        RECT 505.200 63.600 506.600 64.400 ;
        RECT 505.800 62.200 506.600 63.600 ;
        RECT 510.600 64.400 511.400 65.600 ;
        RECT 510.600 63.600 512.400 64.400 ;
        RECT 510.600 62.200 511.400 63.600 ;
        RECT 516.400 62.200 517.200 66.000 ;
        RECT 518.000 62.200 518.800 67.400 ;
        RECT 521.800 67.400 522.600 68.600 ;
        RECT 521.800 66.800 523.600 67.400 ;
        RECT 522.800 66.200 523.600 66.800 ;
        RECT 527.600 66.400 528.400 69.200 ;
        RECT 530.800 68.600 534.000 69.400 ;
        RECT 537.800 68.600 539.800 69.400 ;
        RECT 548.400 69.000 549.200 74.600 ;
        RECT 530.400 67.800 531.200 68.000 ;
        RECT 530.400 67.200 534.800 67.800 ;
        RECT 534.000 67.000 534.800 67.200 ;
        RECT 535.600 66.800 536.400 68.400 ;
        RECT 522.800 65.400 525.200 66.200 ;
        RECT 527.600 65.600 528.600 66.400 ;
        RECT 531.600 65.600 533.200 66.400 ;
        RECT 534.000 66.200 534.800 66.400 ;
        RECT 537.800 66.200 538.600 68.600 ;
        RECT 540.400 68.200 549.200 69.000 ;
        RECT 543.800 66.800 546.800 67.600 ;
        RECT 543.800 66.200 544.600 66.800 ;
        RECT 534.000 65.600 538.600 66.200 ;
        RECT 524.400 62.200 525.200 65.400 ;
        RECT 542.000 65.400 544.600 66.200 ;
        RECT 526.000 62.200 526.800 65.000 ;
        RECT 527.600 62.200 528.400 65.000 ;
        RECT 529.200 62.200 530.000 65.000 ;
        RECT 530.800 62.200 531.600 65.000 ;
        RECT 534.000 62.200 534.800 65.000 ;
        RECT 537.200 62.200 538.000 65.000 ;
        RECT 538.800 62.200 539.600 65.000 ;
        RECT 540.400 62.200 541.200 65.000 ;
        RECT 542.000 62.200 542.800 65.400 ;
        RECT 548.400 62.200 549.200 68.200 ;
        RECT 1.200 55.600 2.000 57.200 ;
        RECT 2.800 50.300 3.600 59.800 ;
        RECT 7.000 58.400 7.800 59.800 ;
        RECT 7.000 57.600 8.400 58.400 ;
        RECT 7.000 56.400 7.800 57.600 ;
        RECT 6.000 55.800 7.800 56.400 ;
        RECT 4.400 53.600 5.200 55.200 ;
        RECT 4.400 50.300 5.200 50.400 ;
        RECT 2.800 49.700 5.200 50.300 ;
        RECT 2.800 42.200 3.600 49.700 ;
        RECT 4.400 49.600 5.200 49.700 ;
        RECT 6.000 42.200 6.800 55.800 ;
        RECT 9.200 55.600 10.000 57.200 ;
        RECT 7.600 50.300 8.400 50.400 ;
        RECT 10.800 50.300 11.600 59.800 ;
        RECT 15.000 58.400 15.800 59.800 ;
        RECT 15.000 57.600 16.400 58.400 ;
        RECT 15.000 56.400 15.800 57.600 ;
        RECT 14.000 55.800 15.800 56.400 ;
        RECT 17.200 56.000 18.000 59.800 ;
        RECT 20.400 59.200 24.400 59.800 ;
        RECT 20.400 56.000 21.200 59.200 ;
        RECT 17.200 55.800 21.200 56.000 ;
        RECT 22.000 55.800 22.800 58.600 ;
        RECT 23.600 55.800 24.400 59.200 ;
        RECT 25.200 56.000 26.000 59.800 ;
        RECT 28.400 59.200 32.400 59.800 ;
        RECT 28.400 56.000 29.200 59.200 ;
        RECT 25.200 55.800 29.200 56.000 ;
        RECT 30.000 55.800 30.800 58.600 ;
        RECT 31.600 55.800 32.400 59.200 ;
        RECT 35.800 58.400 36.600 59.800 ;
        RECT 34.800 57.600 36.600 58.400 ;
        RECT 35.800 56.400 36.600 57.600 ;
        RECT 34.800 55.800 36.600 56.400 ;
        RECT 12.400 53.600 13.200 55.200 ;
        RECT 7.600 49.700 11.600 50.300 ;
        RECT 7.600 48.800 8.400 49.700 ;
        RECT 10.800 42.200 11.600 49.700 ;
        RECT 14.000 42.200 14.800 55.800 ;
        RECT 17.400 55.400 21.000 55.800 ;
        RECT 18.000 54.400 18.800 54.800 ;
        RECT 22.200 54.400 22.800 55.800 ;
        RECT 25.400 55.400 29.000 55.800 ;
        RECT 26.000 54.400 26.800 54.800 ;
        RECT 30.200 54.400 30.800 55.800 ;
        RECT 17.200 53.800 18.800 54.400 ;
        RECT 20.400 53.800 22.800 54.400 ;
        RECT 17.200 53.600 18.000 53.800 ;
        RECT 20.400 53.600 21.200 53.800 ;
        RECT 18.800 51.600 19.600 53.200 ;
        RECT 15.600 48.800 16.400 50.400 ;
        RECT 20.400 50.200 21.000 53.600 ;
        RECT 22.000 51.600 22.800 53.200 ;
        RECT 23.600 52.800 24.400 54.400 ;
        RECT 25.200 53.800 26.800 54.400 ;
        RECT 28.400 53.800 30.800 54.400 ;
        RECT 25.200 53.600 26.000 53.800 ;
        RECT 28.400 53.600 29.200 53.800 ;
        RECT 26.800 51.600 27.600 53.200 ;
        RECT 28.400 50.200 29.000 53.600 ;
        RECT 30.000 51.600 30.800 53.200 ;
        RECT 31.600 52.800 32.400 54.400 ;
        RECT 33.200 53.600 34.000 55.200 ;
        RECT 19.800 42.200 21.800 50.200 ;
        RECT 27.800 44.400 29.800 50.200 ;
        RECT 26.800 43.600 29.800 44.400 ;
        RECT 27.800 42.200 29.800 43.600 ;
        RECT 34.800 42.200 35.600 55.800 ;
        RECT 36.400 50.300 37.200 50.400 ;
        RECT 38.000 50.300 38.800 59.800 ;
        RECT 39.600 55.600 40.400 57.200 ;
        RECT 36.400 49.700 38.800 50.300 ;
        RECT 36.400 48.800 37.200 49.700 ;
        RECT 38.000 42.200 38.800 49.700 ;
        RECT 41.200 53.800 42.000 59.800 ;
        RECT 47.600 56.600 48.400 59.800 ;
        RECT 49.200 57.000 50.000 59.800 ;
        RECT 50.800 57.000 51.600 59.800 ;
        RECT 52.400 57.000 53.200 59.800 ;
        RECT 55.600 57.000 56.400 59.800 ;
        RECT 58.800 57.000 59.600 59.800 ;
        RECT 60.400 57.000 61.200 59.800 ;
        RECT 62.000 57.000 62.800 59.800 ;
        RECT 63.600 57.000 64.400 59.800 ;
        RECT 45.800 55.800 48.400 56.600 ;
        RECT 65.200 56.600 66.000 59.800 ;
        RECT 51.800 55.800 56.400 56.400 ;
        RECT 45.800 55.200 46.600 55.800 ;
        RECT 43.600 54.400 46.600 55.200 ;
        RECT 41.200 53.000 50.000 53.800 ;
        RECT 51.800 53.400 52.600 55.800 ;
        RECT 55.600 55.600 56.400 55.800 ;
        RECT 57.200 55.600 58.800 56.400 ;
        RECT 61.800 55.600 62.800 56.400 ;
        RECT 65.200 55.800 67.600 56.600 ;
        RECT 54.000 53.600 54.800 55.200 ;
        RECT 55.600 54.800 56.400 55.000 ;
        RECT 55.600 54.200 60.000 54.800 ;
        RECT 59.200 54.000 60.000 54.200 ;
        RECT 41.200 47.400 42.000 53.000 ;
        RECT 50.600 52.600 52.600 53.400 ;
        RECT 56.400 52.600 59.600 53.400 ;
        RECT 62.000 52.800 62.800 55.600 ;
        RECT 66.800 55.200 67.600 55.800 ;
        RECT 66.800 54.600 68.600 55.200 ;
        RECT 67.800 53.400 68.600 54.600 ;
        RECT 71.600 54.600 72.400 59.800 ;
        RECT 73.200 56.300 74.000 59.800 ;
        RECT 74.800 56.300 75.600 56.400 ;
        RECT 73.200 55.700 75.600 56.300 ;
        RECT 73.200 55.200 74.200 55.700 ;
        RECT 74.800 55.600 75.600 55.700 ;
        RECT 71.600 54.000 72.800 54.600 ;
        RECT 67.800 52.600 71.600 53.400 ;
        RECT 42.600 52.000 43.400 52.200 ;
        RECT 46.000 52.000 46.800 52.400 ;
        RECT 47.600 52.000 48.400 52.400 ;
        RECT 65.200 52.000 66.000 52.600 ;
        RECT 72.200 52.000 72.800 54.000 ;
        RECT 42.600 51.400 66.000 52.000 ;
        RECT 72.000 51.400 72.800 52.000 ;
        RECT 72.000 49.600 72.600 51.400 ;
        RECT 73.400 50.800 74.200 55.200 ;
        RECT 78.000 55.200 78.800 59.800 ;
        RECT 81.200 55.200 82.000 59.800 ;
        RECT 84.400 55.200 85.200 59.800 ;
        RECT 87.600 55.200 88.400 59.800 ;
        RECT 78.000 54.400 79.800 55.200 ;
        RECT 81.200 54.400 83.400 55.200 ;
        RECT 84.400 54.400 86.600 55.200 ;
        RECT 87.600 54.400 90.000 55.200 ;
        RECT 79.000 53.800 79.800 54.400 ;
        RECT 82.600 53.800 83.400 54.400 ;
        RECT 85.800 53.800 86.600 54.400 ;
        RECT 79.000 53.000 81.600 53.800 ;
        RECT 82.600 53.000 85.000 53.800 ;
        RECT 85.800 53.000 88.400 53.800 ;
        RECT 79.000 51.600 79.800 53.000 ;
        RECT 82.600 51.600 83.400 53.000 ;
        RECT 85.800 51.600 86.600 53.000 ;
        RECT 89.200 51.600 90.000 54.400 ;
        RECT 50.800 49.400 51.600 49.600 ;
        RECT 46.200 49.000 51.600 49.400 ;
        RECT 45.400 48.800 51.600 49.000 ;
        RECT 52.600 49.000 61.200 49.600 ;
        RECT 42.800 48.000 44.400 48.800 ;
        RECT 45.400 48.200 46.800 48.800 ;
        RECT 52.600 48.200 53.200 49.000 ;
        RECT 60.400 48.800 61.200 49.000 ;
        RECT 63.600 49.000 72.600 49.600 ;
        RECT 63.600 48.800 64.400 49.000 ;
        RECT 43.800 47.600 44.400 48.000 ;
        RECT 47.400 47.600 53.200 48.200 ;
        RECT 53.800 47.600 56.400 48.400 ;
        RECT 41.200 46.800 43.200 47.400 ;
        RECT 43.800 46.800 48.000 47.600 ;
        RECT 42.600 46.200 43.200 46.800 ;
        RECT 42.600 45.600 43.600 46.200 ;
        RECT 42.800 42.200 43.600 45.600 ;
        RECT 46.000 42.200 46.800 46.800 ;
        RECT 49.200 42.200 50.000 45.000 ;
        RECT 50.800 42.200 51.600 45.000 ;
        RECT 52.400 42.200 53.200 47.000 ;
        RECT 55.600 42.200 56.400 47.000 ;
        RECT 58.800 42.200 59.600 48.400 ;
        RECT 66.800 47.600 69.400 48.400 ;
        RECT 62.000 46.800 66.200 47.600 ;
        RECT 60.400 42.200 61.200 45.000 ;
        RECT 62.000 42.200 62.800 45.000 ;
        RECT 63.600 42.200 64.400 45.000 ;
        RECT 66.800 42.200 67.600 47.600 ;
        RECT 72.000 47.400 72.600 49.000 ;
        RECT 70.000 46.800 72.600 47.400 ;
        RECT 73.200 50.000 74.200 50.800 ;
        RECT 78.000 50.800 79.800 51.600 ;
        RECT 81.200 50.800 83.400 51.600 ;
        RECT 84.400 50.800 86.600 51.600 ;
        RECT 87.600 50.800 90.000 51.600 ;
        RECT 90.800 53.800 91.600 59.800 ;
        RECT 97.200 56.600 98.000 59.800 ;
        RECT 98.800 57.000 99.600 59.800 ;
        RECT 100.400 57.000 101.200 59.800 ;
        RECT 102.000 57.000 102.800 59.800 ;
        RECT 105.200 57.000 106.000 59.800 ;
        RECT 108.400 57.000 109.200 59.800 ;
        RECT 110.000 57.000 110.800 59.800 ;
        RECT 111.600 57.000 112.400 59.800 ;
        RECT 113.200 57.000 114.000 59.800 ;
        RECT 95.400 55.800 98.000 56.600 ;
        RECT 114.800 56.600 115.600 59.800 ;
        RECT 101.400 55.800 106.000 56.400 ;
        RECT 95.400 55.200 96.200 55.800 ;
        RECT 93.200 54.400 96.200 55.200 ;
        RECT 90.800 53.000 99.600 53.800 ;
        RECT 101.400 53.400 102.200 55.800 ;
        RECT 105.200 55.600 106.000 55.800 ;
        RECT 106.800 55.600 108.400 56.400 ;
        RECT 111.400 55.600 112.400 56.400 ;
        RECT 114.800 55.800 117.200 56.600 ;
        RECT 103.600 53.600 104.400 55.200 ;
        RECT 105.200 54.800 106.000 55.000 ;
        RECT 105.200 54.200 109.600 54.800 ;
        RECT 108.800 54.000 109.600 54.200 ;
        RECT 70.000 42.200 70.800 46.800 ;
        RECT 73.200 42.200 74.000 50.000 ;
        RECT 78.000 42.200 78.800 50.800 ;
        RECT 81.200 42.200 82.000 50.800 ;
        RECT 84.400 42.200 85.200 50.800 ;
        RECT 87.600 42.200 88.400 50.800 ;
        RECT 90.800 47.400 91.600 53.000 ;
        RECT 100.200 52.600 102.200 53.400 ;
        RECT 106.000 52.600 109.200 53.400 ;
        RECT 111.600 52.800 112.400 55.600 ;
        RECT 116.400 55.200 117.200 55.800 ;
        RECT 116.400 54.600 118.200 55.200 ;
        RECT 117.400 53.400 118.200 54.600 ;
        RECT 121.200 54.600 122.000 59.800 ;
        RECT 122.800 56.000 123.600 59.800 ;
        RECT 134.000 57.600 134.800 59.800 ;
        RECT 122.800 55.200 123.800 56.000 ;
        RECT 132.400 55.600 133.200 57.200 ;
        RECT 121.200 54.000 122.400 54.600 ;
        RECT 117.400 52.600 121.200 53.400 ;
        RECT 121.800 52.000 122.400 54.000 ;
        RECT 121.600 51.400 122.400 52.000 ;
        RECT 120.200 50.800 121.000 51.000 ;
        RECT 94.000 50.200 121.000 50.800 ;
        RECT 94.000 49.600 94.800 50.200 ;
        RECT 97.400 50.000 98.200 50.200 ;
        RECT 121.600 49.600 122.200 51.400 ;
        RECT 123.000 50.800 123.800 55.200 ;
        RECT 134.200 54.400 134.800 57.600 ;
        RECT 135.600 56.300 136.400 56.400 ;
        RECT 137.200 56.300 138.000 59.800 ;
        RECT 142.000 57.800 142.800 59.800 ;
        RECT 135.600 55.700 138.000 56.300 ;
        RECT 135.600 55.600 136.400 55.700 ;
        RECT 134.000 53.600 134.800 54.400 ;
        RECT 100.400 49.400 101.200 49.600 ;
        RECT 95.800 49.000 101.200 49.400 ;
        RECT 95.000 48.800 101.200 49.000 ;
        RECT 102.200 49.000 110.800 49.600 ;
        RECT 92.400 48.000 94.000 48.800 ;
        RECT 95.000 48.200 96.400 48.800 ;
        RECT 102.200 48.200 102.800 49.000 ;
        RECT 110.000 48.800 110.800 49.000 ;
        RECT 113.200 49.000 122.200 49.600 ;
        RECT 113.200 48.800 114.000 49.000 ;
        RECT 93.400 47.600 94.000 48.000 ;
        RECT 97.000 47.600 102.800 48.200 ;
        RECT 103.400 47.600 106.000 48.400 ;
        RECT 90.800 46.800 92.800 47.400 ;
        RECT 93.400 46.800 97.600 47.600 ;
        RECT 92.200 46.200 92.800 46.800 ;
        RECT 92.200 45.600 93.200 46.200 ;
        RECT 92.400 42.200 93.200 45.600 ;
        RECT 95.600 42.200 96.400 46.800 ;
        RECT 98.800 42.200 99.600 45.000 ;
        RECT 100.400 42.200 101.200 45.000 ;
        RECT 102.000 42.200 102.800 47.000 ;
        RECT 105.200 42.200 106.000 47.000 ;
        RECT 108.400 42.200 109.200 48.400 ;
        RECT 116.400 47.600 119.000 48.400 ;
        RECT 111.600 46.800 115.800 47.600 ;
        RECT 110.000 42.200 110.800 45.000 ;
        RECT 111.600 42.200 112.400 45.000 ;
        RECT 113.200 42.200 114.000 45.000 ;
        RECT 116.400 42.200 117.200 47.600 ;
        RECT 121.600 47.400 122.200 49.000 ;
        RECT 119.600 46.800 122.200 47.400 ;
        RECT 122.800 50.000 123.800 50.800 ;
        RECT 134.200 50.200 134.800 53.600 ;
        RECT 135.600 50.800 136.400 52.400 ;
        RECT 137.200 52.300 138.000 55.700 ;
        RECT 138.800 55.600 139.600 57.200 ;
        RECT 142.000 54.400 142.600 57.800 ;
        RECT 143.600 56.300 144.400 57.200 ;
        RECT 145.800 56.400 146.600 59.800 ;
        RECT 152.600 56.400 153.400 59.800 ;
        RECT 156.400 57.800 157.200 59.800 ;
        RECT 160.200 58.400 161.000 59.800 ;
        RECT 145.800 56.300 147.600 56.400 ;
        RECT 143.600 55.700 147.600 56.300 ;
        RECT 143.600 55.600 144.400 55.700 ;
        RECT 142.000 53.600 142.800 54.400 ;
        RECT 140.400 52.300 141.200 52.400 ;
        RECT 137.200 51.700 141.200 52.300 ;
        RECT 119.600 42.200 120.400 46.800 ;
        RECT 122.800 42.200 123.600 50.000 ;
        RECT 134.000 49.400 135.800 50.200 ;
        RECT 135.000 42.200 135.800 49.400 ;
        RECT 137.200 42.200 138.000 51.700 ;
        RECT 140.400 50.800 141.200 51.700 ;
        RECT 142.000 50.200 142.600 53.600 ;
        RECT 141.000 49.400 142.800 50.200 ;
        RECT 141.000 44.400 141.800 49.400 ;
        RECT 145.200 48.800 146.000 50.400 ;
        RECT 141.000 43.600 142.800 44.400 ;
        RECT 141.000 42.200 141.800 43.600 ;
        RECT 146.800 42.200 147.600 55.700 ;
        RECT 151.600 55.800 153.400 56.400 ;
        RECT 148.400 54.300 149.200 55.200 ;
        RECT 150.000 54.300 150.800 55.200 ;
        RECT 148.400 53.700 150.800 54.300 ;
        RECT 148.400 53.600 149.200 53.700 ;
        RECT 150.000 53.600 150.800 53.700 ;
        RECT 148.400 52.300 149.200 52.400 ;
        RECT 151.600 52.300 152.400 55.800 ;
        RECT 154.800 55.600 155.600 57.200 ;
        RECT 156.600 54.400 157.200 57.800 ;
        RECT 159.600 57.600 161.000 58.400 ;
        RECT 160.200 56.400 161.000 57.600 ;
        RECT 160.200 55.800 162.000 56.400 ;
        RECT 156.400 53.600 157.200 54.400 ;
        RECT 156.600 52.300 157.200 53.600 ;
        RECT 148.400 51.700 152.400 52.300 ;
        RECT 148.400 51.600 149.200 51.700 ;
        RECT 151.600 42.200 152.400 51.700 ;
        RECT 153.300 51.700 157.200 52.300 ;
        RECT 153.300 50.400 153.900 51.700 ;
        RECT 153.200 48.800 154.000 50.400 ;
        RECT 156.600 50.200 157.200 51.700 ;
        RECT 158.000 50.800 158.800 52.400 ;
        RECT 156.400 49.400 158.200 50.200 ;
        RECT 157.400 42.200 158.200 49.400 ;
        RECT 159.600 48.800 160.400 50.400 ;
        RECT 161.200 42.200 162.000 55.800 ;
        RECT 162.800 53.600 163.600 55.200 ;
        RECT 162.800 52.300 163.600 52.400 ;
        RECT 164.400 52.300 165.200 59.800 ;
        RECT 169.200 57.600 170.000 59.800 ;
        RECT 166.000 55.600 166.800 57.200 ;
        RECT 169.200 54.400 169.800 57.600 ;
        RECT 170.800 55.600 171.600 57.200 ;
        RECT 169.200 53.600 170.000 54.400 ;
        RECT 170.900 54.300 171.500 55.600 ;
        RECT 172.400 54.300 173.200 55.200 ;
        RECT 170.900 53.700 173.200 54.300 ;
        RECT 172.400 53.600 173.200 53.700 ;
        RECT 162.800 51.700 165.200 52.300 ;
        RECT 162.800 51.600 163.600 51.700 ;
        RECT 164.400 42.200 165.200 51.700 ;
        RECT 166.000 52.300 166.800 52.400 ;
        RECT 167.600 52.300 168.400 52.400 ;
        RECT 166.000 51.700 168.400 52.300 ;
        RECT 166.000 51.600 166.800 51.700 ;
        RECT 167.600 50.800 168.400 51.700 ;
        RECT 169.200 50.200 169.800 53.600 ;
        RECT 168.200 49.400 170.000 50.200 ;
        RECT 168.200 42.200 169.000 49.400 ;
        RECT 174.000 42.200 174.800 59.800 ;
        RECT 177.200 53.800 178.000 59.800 ;
        RECT 183.600 56.600 184.400 59.800 ;
        RECT 185.200 57.000 186.000 59.800 ;
        RECT 186.800 57.000 187.600 59.800 ;
        RECT 188.400 57.000 189.200 59.800 ;
        RECT 191.600 57.000 192.400 59.800 ;
        RECT 194.800 57.000 195.600 59.800 ;
        RECT 196.400 57.000 197.200 59.800 ;
        RECT 198.000 57.000 198.800 59.800 ;
        RECT 199.600 57.000 200.400 59.800 ;
        RECT 181.800 55.800 184.400 56.600 ;
        RECT 201.200 56.600 202.000 59.800 ;
        RECT 187.800 55.800 192.400 56.400 ;
        RECT 181.800 55.200 182.600 55.800 ;
        RECT 179.600 54.400 182.600 55.200 ;
        RECT 177.200 53.000 186.000 53.800 ;
        RECT 187.800 53.400 188.600 55.800 ;
        RECT 191.600 55.600 192.400 55.800 ;
        RECT 193.200 55.600 194.800 56.400 ;
        RECT 197.800 55.600 198.800 56.400 ;
        RECT 201.200 55.800 203.600 56.600 ;
        RECT 190.000 53.600 190.800 55.200 ;
        RECT 191.600 54.800 192.400 55.000 ;
        RECT 191.600 54.200 196.000 54.800 ;
        RECT 195.200 54.000 196.000 54.200 ;
        RECT 177.200 47.400 178.000 53.000 ;
        RECT 186.600 52.600 188.600 53.400 ;
        RECT 192.400 52.600 195.600 53.400 ;
        RECT 198.000 52.800 198.800 55.600 ;
        RECT 202.800 55.200 203.600 55.800 ;
        RECT 202.800 54.600 204.600 55.200 ;
        RECT 203.800 53.400 204.600 54.600 ;
        RECT 207.600 54.600 208.400 59.800 ;
        RECT 209.200 56.000 210.000 59.800 ;
        RECT 212.400 56.000 213.200 59.800 ;
        RECT 215.600 56.000 216.400 59.800 ;
        RECT 209.200 55.200 210.200 56.000 ;
        RECT 212.400 55.800 216.400 56.000 ;
        RECT 217.200 55.800 218.000 59.800 ;
        RECT 218.800 55.800 219.600 59.800 ;
        RECT 220.400 56.000 221.200 59.800 ;
        RECT 223.600 56.000 224.400 59.800 ;
        RECT 220.400 55.800 224.400 56.000 ;
        RECT 212.600 55.400 216.200 55.800 ;
        RECT 207.600 54.000 208.800 54.600 ;
        RECT 203.800 52.600 207.600 53.400 ;
        RECT 208.200 52.000 208.800 54.000 ;
        RECT 208.000 51.400 208.800 52.000 ;
        RECT 206.600 50.800 207.400 51.000 ;
        RECT 180.400 50.200 207.400 50.800 ;
        RECT 180.400 49.600 181.200 50.200 ;
        RECT 183.800 50.000 184.600 50.200 ;
        RECT 208.000 49.600 208.600 51.400 ;
        RECT 209.400 50.800 210.200 55.200 ;
        RECT 213.200 54.400 214.000 54.800 ;
        RECT 217.200 54.400 217.800 55.800 ;
        RECT 219.000 54.400 219.600 55.800 ;
        RECT 220.600 55.400 224.200 55.800 ;
        RECT 222.800 54.400 223.600 54.800 ;
        RECT 212.400 53.800 214.000 54.400 ;
        RECT 212.400 53.600 213.200 53.800 ;
        RECT 215.400 53.600 218.000 54.400 ;
        RECT 218.800 53.600 221.400 54.400 ;
        RECT 222.800 53.800 224.400 54.400 ;
        RECT 223.600 53.600 224.400 53.800 ;
        RECT 225.200 54.300 226.000 59.800 ;
        RECT 226.800 55.600 227.600 57.200 ;
        RECT 228.400 56.000 229.200 59.800 ;
        RECT 231.600 56.000 232.400 59.800 ;
        RECT 228.400 55.800 232.400 56.000 ;
        RECT 233.200 56.300 234.000 59.800 ;
        RECT 234.800 56.300 235.600 56.400 ;
        RECT 228.600 55.400 232.200 55.800 ;
        RECT 233.200 55.700 235.600 56.300 ;
        RECT 236.400 56.000 237.200 59.800 ;
        RECT 229.200 54.400 230.000 54.800 ;
        RECT 233.200 54.400 233.800 55.700 ;
        RECT 234.800 55.600 235.600 55.700 ;
        RECT 236.200 55.200 237.200 56.000 ;
        RECT 228.400 54.300 230.000 54.400 ;
        RECT 225.200 53.800 230.000 54.300 ;
        RECT 225.200 53.700 229.200 53.800 ;
        RECT 214.000 51.600 214.800 53.200 ;
        RECT 215.400 52.400 216.000 53.600 ;
        RECT 215.400 51.600 216.400 52.400 ;
        RECT 220.800 52.300 221.400 53.600 ;
        RECT 217.300 51.700 221.400 52.300 ;
        RECT 186.800 49.400 187.600 49.600 ;
        RECT 182.200 49.000 187.600 49.400 ;
        RECT 181.400 48.800 187.600 49.000 ;
        RECT 188.600 49.000 197.200 49.600 ;
        RECT 178.800 48.000 180.400 48.800 ;
        RECT 181.400 48.200 182.800 48.800 ;
        RECT 188.600 48.200 189.200 49.000 ;
        RECT 196.400 48.800 197.200 49.000 ;
        RECT 199.600 49.000 208.600 49.600 ;
        RECT 199.600 48.800 200.400 49.000 ;
        RECT 179.800 47.600 180.400 48.000 ;
        RECT 183.400 47.600 189.200 48.200 ;
        RECT 189.800 47.600 192.400 48.400 ;
        RECT 177.200 46.800 179.200 47.400 ;
        RECT 179.800 46.800 184.000 47.600 ;
        RECT 178.600 46.200 179.200 46.800 ;
        RECT 178.600 45.600 179.600 46.200 ;
        RECT 178.800 42.200 179.600 45.600 ;
        RECT 182.000 42.200 182.800 46.800 ;
        RECT 185.200 42.200 186.000 45.000 ;
        RECT 186.800 42.200 187.600 45.000 ;
        RECT 188.400 42.200 189.200 47.000 ;
        RECT 191.600 42.200 192.400 47.000 ;
        RECT 194.800 42.200 195.600 48.400 ;
        RECT 202.800 47.600 205.400 48.400 ;
        RECT 198.000 46.800 202.200 47.600 ;
        RECT 196.400 42.200 197.200 45.000 ;
        RECT 198.000 42.200 198.800 45.000 ;
        RECT 199.600 42.200 200.400 45.000 ;
        RECT 202.800 42.200 203.600 47.600 ;
        RECT 208.000 47.400 208.600 49.000 ;
        RECT 206.000 46.800 208.600 47.400 ;
        RECT 209.200 50.000 210.200 50.800 ;
        RECT 215.400 50.200 216.000 51.600 ;
        RECT 217.300 50.400 217.900 51.700 ;
        RECT 217.200 50.200 218.000 50.400 ;
        RECT 209.200 48.300 210.000 50.000 ;
        RECT 215.000 49.600 216.000 50.200 ;
        RECT 216.600 49.600 218.000 50.200 ;
        RECT 218.800 50.200 219.600 50.400 ;
        RECT 220.800 50.200 221.400 51.700 ;
        RECT 222.000 51.600 222.800 53.200 ;
        RECT 218.800 49.600 220.200 50.200 ;
        RECT 220.800 49.600 221.800 50.200 ;
        RECT 210.800 48.300 211.600 48.400 ;
        RECT 209.200 47.700 211.600 48.300 ;
        RECT 206.000 42.200 206.800 46.800 ;
        RECT 209.200 42.200 210.000 47.700 ;
        RECT 210.800 47.600 211.600 47.700 ;
        RECT 215.000 42.200 215.800 49.600 ;
        RECT 216.600 48.400 217.200 49.600 ;
        RECT 216.400 47.600 217.200 48.400 ;
        RECT 219.600 48.400 220.200 49.600 ;
        RECT 219.600 47.600 220.400 48.400 ;
        RECT 221.000 42.200 221.800 49.600 ;
        RECT 225.200 48.300 226.000 53.700 ;
        RECT 228.400 53.600 229.200 53.700 ;
        RECT 231.400 53.600 234.000 54.400 ;
        RECT 230.000 51.600 230.800 53.200 ;
        RECT 231.400 50.200 232.000 53.600 ;
        RECT 236.200 50.800 237.000 55.200 ;
        RECT 238.000 54.600 238.800 59.800 ;
        RECT 244.400 56.600 245.200 59.800 ;
        RECT 246.000 57.000 246.800 59.800 ;
        RECT 247.600 57.000 248.400 59.800 ;
        RECT 249.200 57.000 250.000 59.800 ;
        RECT 250.800 57.000 251.600 59.800 ;
        RECT 254.000 57.000 254.800 59.800 ;
        RECT 257.200 57.000 258.000 59.800 ;
        RECT 258.800 57.000 259.600 59.800 ;
        RECT 260.400 57.000 261.200 59.800 ;
        RECT 242.800 55.800 245.200 56.600 ;
        RECT 262.000 56.600 262.800 59.800 ;
        RECT 242.800 55.200 243.600 55.800 ;
        RECT 237.600 54.000 238.800 54.600 ;
        RECT 241.800 54.600 243.600 55.200 ;
        RECT 247.600 55.600 248.600 56.400 ;
        RECT 251.600 55.600 253.200 56.400 ;
        RECT 254.000 55.800 258.600 56.400 ;
        RECT 262.000 55.800 264.600 56.600 ;
        RECT 254.000 55.600 254.800 55.800 ;
        RECT 237.600 52.000 238.200 54.000 ;
        RECT 241.800 53.400 242.600 54.600 ;
        RECT 238.800 52.600 242.600 53.400 ;
        RECT 247.600 52.800 248.400 55.600 ;
        RECT 254.000 54.800 254.800 55.000 ;
        RECT 250.400 54.200 254.800 54.800 ;
        RECT 250.400 54.000 251.200 54.200 ;
        RECT 255.600 53.600 256.400 55.200 ;
        RECT 257.800 53.400 258.600 55.800 ;
        RECT 263.800 55.200 264.600 55.800 ;
        RECT 263.800 54.400 266.800 55.200 ;
        RECT 268.400 53.800 269.200 59.800 ;
        RECT 270.000 55.200 270.800 59.800 ;
        RECT 270.000 54.600 272.200 55.200 ;
        RECT 250.800 52.600 254.000 53.400 ;
        RECT 257.800 52.600 259.800 53.400 ;
        RECT 260.400 53.000 269.200 53.800 ;
        RECT 237.600 51.400 238.400 52.000 ;
        RECT 233.200 50.200 234.000 50.400 ;
        RECT 231.000 49.600 232.000 50.200 ;
        RECT 232.600 49.600 234.000 50.200 ;
        RECT 236.200 50.000 237.200 50.800 ;
        RECT 226.800 48.300 227.600 48.400 ;
        RECT 225.200 47.700 227.600 48.300 ;
        RECT 225.200 42.200 226.000 47.700 ;
        RECT 226.800 47.600 227.600 47.700 ;
        RECT 231.000 42.200 231.800 49.600 ;
        RECT 232.600 48.400 233.200 49.600 ;
        RECT 232.400 47.600 233.200 48.400 ;
        RECT 236.400 42.200 237.200 50.000 ;
        RECT 237.800 49.600 238.400 51.400 ;
        RECT 239.000 50.800 239.800 51.000 ;
        RECT 239.000 50.200 266.000 50.800 ;
        RECT 261.800 50.000 262.800 50.200 ;
        RECT 265.200 49.600 266.000 50.200 ;
        RECT 237.800 49.000 246.800 49.600 ;
        RECT 237.800 47.400 238.400 49.000 ;
        RECT 246.000 48.800 246.800 49.000 ;
        RECT 249.200 49.000 257.800 49.600 ;
        RECT 249.200 48.800 250.000 49.000 ;
        RECT 241.000 47.600 243.600 48.400 ;
        RECT 237.800 46.800 240.400 47.400 ;
        RECT 239.600 42.200 240.400 46.800 ;
        RECT 242.800 42.200 243.600 47.600 ;
        RECT 244.200 46.800 248.400 47.600 ;
        RECT 246.000 42.200 246.800 45.000 ;
        RECT 247.600 42.200 248.400 45.000 ;
        RECT 249.200 42.200 250.000 45.000 ;
        RECT 250.800 42.200 251.600 48.400 ;
        RECT 254.000 47.600 256.600 48.400 ;
        RECT 257.200 48.200 257.800 49.000 ;
        RECT 258.800 49.400 259.600 49.600 ;
        RECT 258.800 49.000 264.200 49.400 ;
        RECT 258.800 48.800 265.000 49.000 ;
        RECT 263.600 48.200 265.000 48.800 ;
        RECT 257.200 47.600 263.000 48.200 ;
        RECT 266.000 48.000 267.600 48.800 ;
        RECT 266.000 47.600 266.600 48.000 ;
        RECT 254.000 42.200 254.800 47.000 ;
        RECT 257.200 42.200 258.000 47.000 ;
        RECT 262.400 46.800 266.600 47.600 ;
        RECT 268.400 47.400 269.200 53.000 ;
        RECT 271.600 51.600 272.200 54.600 ;
        RECT 273.200 52.400 274.000 59.800 ;
        RECT 271.600 50.800 272.800 51.600 ;
        RECT 271.600 50.200 272.200 50.800 ;
        RECT 273.400 50.200 274.000 52.400 ;
        RECT 267.200 46.800 269.200 47.400 ;
        RECT 270.000 49.600 272.200 50.200 ;
        RECT 258.800 42.200 259.600 45.000 ;
        RECT 260.400 42.200 261.200 45.000 ;
        RECT 263.600 42.200 264.400 46.800 ;
        RECT 267.200 46.200 267.800 46.800 ;
        RECT 266.800 45.600 267.800 46.200 ;
        RECT 266.800 42.200 267.600 45.600 ;
        RECT 270.000 42.200 270.800 49.600 ;
        RECT 273.200 44.300 274.000 50.200 ;
        RECT 281.200 53.800 282.000 59.800 ;
        RECT 287.600 56.600 288.400 59.800 ;
        RECT 289.200 57.000 290.000 59.800 ;
        RECT 290.800 57.000 291.600 59.800 ;
        RECT 292.400 57.000 293.200 59.800 ;
        RECT 295.600 57.000 296.400 59.800 ;
        RECT 298.800 57.000 299.600 59.800 ;
        RECT 300.400 57.000 301.200 59.800 ;
        RECT 302.000 57.000 302.800 59.800 ;
        RECT 303.600 57.000 304.400 59.800 ;
        RECT 285.800 55.800 288.400 56.600 ;
        RECT 305.200 56.600 306.000 59.800 ;
        RECT 291.800 55.800 296.400 56.400 ;
        RECT 285.800 55.200 286.600 55.800 ;
        RECT 283.600 54.400 286.600 55.200 ;
        RECT 281.200 53.000 290.000 53.800 ;
        RECT 291.800 53.400 292.600 55.800 ;
        RECT 295.600 55.600 296.400 55.800 ;
        RECT 297.200 55.600 298.800 56.400 ;
        RECT 301.800 55.600 302.800 56.400 ;
        RECT 305.200 55.800 307.600 56.600 ;
        RECT 294.000 53.600 294.800 55.200 ;
        RECT 295.600 54.800 296.400 55.000 ;
        RECT 295.600 54.200 300.000 54.800 ;
        RECT 299.200 54.000 300.000 54.200 ;
        RECT 281.200 47.400 282.000 53.000 ;
        RECT 290.600 52.600 292.600 53.400 ;
        RECT 296.400 52.600 299.600 53.400 ;
        RECT 302.000 52.800 302.800 55.600 ;
        RECT 306.800 55.200 307.600 55.800 ;
        RECT 306.800 54.600 308.600 55.200 ;
        RECT 307.800 53.400 308.600 54.600 ;
        RECT 311.600 54.600 312.400 59.800 ;
        RECT 313.200 56.000 314.000 59.800 ;
        RECT 313.200 55.200 314.200 56.000 ;
        RECT 311.600 54.000 312.800 54.600 ;
        RECT 307.800 52.600 311.600 53.400 ;
        RECT 312.200 52.000 312.800 54.000 ;
        RECT 312.000 51.400 312.800 52.000 ;
        RECT 310.600 50.800 311.400 51.000 ;
        RECT 284.400 50.200 311.400 50.800 ;
        RECT 284.400 49.600 285.200 50.200 ;
        RECT 287.800 50.000 288.600 50.200 ;
        RECT 312.000 49.600 312.600 51.400 ;
        RECT 313.400 50.800 314.200 55.200 ;
        RECT 290.800 49.400 291.600 49.600 ;
        RECT 286.200 49.000 291.600 49.400 ;
        RECT 285.400 48.800 291.600 49.000 ;
        RECT 292.600 49.000 301.200 49.600 ;
        RECT 282.800 48.000 284.400 48.800 ;
        RECT 285.400 48.200 286.800 48.800 ;
        RECT 292.600 48.200 293.200 49.000 ;
        RECT 300.400 48.800 301.200 49.000 ;
        RECT 303.600 49.000 312.600 49.600 ;
        RECT 303.600 48.800 304.400 49.000 ;
        RECT 283.800 47.600 284.400 48.000 ;
        RECT 287.400 47.600 293.200 48.200 ;
        RECT 293.800 47.600 296.400 48.400 ;
        RECT 281.200 46.800 283.200 47.400 ;
        RECT 283.800 46.800 288.000 47.600 ;
        RECT 282.600 46.200 283.200 46.800 ;
        RECT 282.600 45.600 283.600 46.200 ;
        RECT 279.600 44.300 280.400 44.400 ;
        RECT 273.200 43.700 280.400 44.300 ;
        RECT 273.200 42.200 274.000 43.700 ;
        RECT 279.600 43.600 280.400 43.700 ;
        RECT 282.800 42.200 283.600 45.600 ;
        RECT 286.000 42.200 286.800 46.800 ;
        RECT 289.200 42.200 290.000 45.000 ;
        RECT 290.800 42.200 291.600 45.000 ;
        RECT 292.400 42.200 293.200 47.000 ;
        RECT 295.600 42.200 296.400 47.000 ;
        RECT 298.800 42.200 299.600 48.400 ;
        RECT 306.800 47.600 309.400 48.400 ;
        RECT 302.000 46.800 306.200 47.600 ;
        RECT 300.400 42.200 301.200 45.000 ;
        RECT 302.000 42.200 302.800 45.000 ;
        RECT 303.600 42.200 304.400 45.000 ;
        RECT 306.800 42.200 307.600 47.600 ;
        RECT 312.000 47.400 312.600 49.000 ;
        RECT 310.000 46.800 312.600 47.400 ;
        RECT 313.200 50.000 314.200 50.800 ;
        RECT 310.000 42.200 310.800 46.800 ;
        RECT 313.200 42.200 314.000 50.000 ;
        RECT 318.000 42.200 318.800 59.800 ;
        RECT 319.600 53.800 320.400 59.800 ;
        RECT 326.000 56.600 326.800 59.800 ;
        RECT 327.600 57.000 328.400 59.800 ;
        RECT 329.200 57.000 330.000 59.800 ;
        RECT 330.800 57.000 331.600 59.800 ;
        RECT 334.000 57.000 334.800 59.800 ;
        RECT 337.200 57.000 338.000 59.800 ;
        RECT 338.800 57.000 339.600 59.800 ;
        RECT 340.400 57.000 341.200 59.800 ;
        RECT 342.000 57.000 342.800 59.800 ;
        RECT 324.200 55.800 326.800 56.600 ;
        RECT 343.600 56.600 344.400 59.800 ;
        RECT 330.200 55.800 334.800 56.400 ;
        RECT 324.200 55.200 325.000 55.800 ;
        RECT 322.000 54.400 325.000 55.200 ;
        RECT 319.600 53.000 328.400 53.800 ;
        RECT 330.200 53.400 331.000 55.800 ;
        RECT 334.000 55.600 334.800 55.800 ;
        RECT 335.600 55.600 337.200 56.400 ;
        RECT 340.200 55.600 341.200 56.400 ;
        RECT 343.600 55.800 346.000 56.600 ;
        RECT 332.400 53.600 333.200 55.200 ;
        RECT 334.000 54.800 334.800 55.000 ;
        RECT 334.000 54.200 338.400 54.800 ;
        RECT 337.600 54.000 338.400 54.200 ;
        RECT 319.600 47.400 320.400 53.000 ;
        RECT 329.000 52.600 331.000 53.400 ;
        RECT 334.800 52.600 338.000 53.400 ;
        RECT 340.400 52.800 341.200 55.600 ;
        RECT 345.200 55.200 346.000 55.800 ;
        RECT 345.200 54.600 347.000 55.200 ;
        RECT 346.200 53.400 347.000 54.600 ;
        RECT 350.000 54.600 350.800 59.800 ;
        RECT 351.600 56.000 352.400 59.800 ;
        RECT 356.400 57.800 357.200 59.800 ;
        RECT 351.600 55.200 352.600 56.000 ;
        RECT 354.800 55.600 355.600 57.200 ;
        RECT 356.600 56.300 357.200 57.800 ;
        RECT 358.000 56.300 358.800 56.400 ;
        RECT 356.500 55.700 358.800 56.300 ;
        RECT 350.000 54.000 351.200 54.600 ;
        RECT 346.200 52.600 350.000 53.400 ;
        RECT 321.200 52.200 322.000 52.400 ;
        RECT 321.000 52.000 322.000 52.200 ;
        RECT 326.000 52.000 326.800 52.400 ;
        RECT 343.600 52.000 344.400 52.600 ;
        RECT 350.600 52.000 351.200 54.000 ;
        RECT 321.000 51.400 344.400 52.000 ;
        RECT 350.400 51.400 351.200 52.000 ;
        RECT 351.800 52.300 352.600 55.200 ;
        RECT 356.600 54.400 357.200 55.700 ;
        RECT 358.000 55.600 358.800 55.700 ;
        RECT 359.600 55.600 360.400 57.200 ;
        RECT 356.400 53.600 357.200 54.400 ;
        RECT 354.800 52.300 355.600 52.400 ;
        RECT 351.800 51.700 355.600 52.300 ;
        RECT 350.400 49.600 351.000 51.400 ;
        RECT 351.800 50.800 352.600 51.700 ;
        RECT 354.800 51.600 355.600 51.700 ;
        RECT 329.200 49.400 330.000 49.600 ;
        RECT 324.600 49.000 330.000 49.400 ;
        RECT 323.800 48.800 330.000 49.000 ;
        RECT 331.000 49.000 339.600 49.600 ;
        RECT 321.200 48.000 322.800 48.800 ;
        RECT 323.800 48.200 325.200 48.800 ;
        RECT 331.000 48.200 331.600 49.000 ;
        RECT 338.800 48.800 339.600 49.000 ;
        RECT 342.000 49.000 351.000 49.600 ;
        RECT 342.000 48.800 342.800 49.000 ;
        RECT 322.200 47.600 322.800 48.000 ;
        RECT 325.800 47.600 331.600 48.200 ;
        RECT 332.200 47.600 334.800 48.400 ;
        RECT 319.600 46.800 321.600 47.400 ;
        RECT 322.200 46.800 326.400 47.600 ;
        RECT 321.000 46.200 321.600 46.800 ;
        RECT 321.000 45.600 322.000 46.200 ;
        RECT 321.200 42.200 322.000 45.600 ;
        RECT 324.400 42.200 325.200 46.800 ;
        RECT 327.600 42.200 328.400 45.000 ;
        RECT 329.200 42.200 330.000 45.000 ;
        RECT 330.800 42.200 331.600 47.000 ;
        RECT 334.000 42.200 334.800 47.000 ;
        RECT 337.200 42.200 338.000 48.400 ;
        RECT 345.200 47.600 347.800 48.400 ;
        RECT 340.400 46.800 344.600 47.600 ;
        RECT 338.800 42.200 339.600 45.000 ;
        RECT 340.400 42.200 341.200 45.000 ;
        RECT 342.000 42.200 342.800 45.000 ;
        RECT 345.200 42.200 346.000 47.600 ;
        RECT 350.400 47.400 351.000 49.000 ;
        RECT 348.400 46.800 351.000 47.400 ;
        RECT 351.600 50.000 352.600 50.800 ;
        RECT 356.600 50.200 357.200 53.600 ;
        RECT 361.200 54.300 362.000 59.800 ;
        RECT 362.800 56.000 363.600 59.800 ;
        RECT 366.000 56.000 366.800 59.800 ;
        RECT 362.800 55.800 366.800 56.000 ;
        RECT 367.600 55.800 368.400 59.800 ;
        RECT 369.800 56.400 370.600 59.800 ;
        RECT 369.800 55.800 371.600 56.400 ;
        RECT 363.000 55.400 366.600 55.800 ;
        RECT 363.600 54.400 364.400 54.800 ;
        RECT 367.600 54.400 368.200 55.800 ;
        RECT 362.800 54.300 364.400 54.400 ;
        RECT 361.200 53.800 364.400 54.300 ;
        RECT 361.200 53.700 363.600 53.800 ;
        RECT 358.000 50.800 358.800 52.400 ;
        RECT 348.400 42.200 349.200 46.800 ;
        RECT 351.600 42.200 352.400 50.000 ;
        RECT 356.400 49.400 358.200 50.200 ;
        RECT 357.400 42.200 358.200 49.400 ;
        RECT 361.200 42.200 362.000 53.700 ;
        RECT 362.800 53.600 363.600 53.700 ;
        RECT 365.800 53.600 368.400 54.400 ;
        RECT 364.400 51.600 365.200 53.200 ;
        RECT 365.800 50.200 366.400 53.600 ;
        RECT 370.800 52.300 371.600 55.800 ;
        RECT 372.400 53.600 373.200 55.200 ;
        RECT 374.000 53.800 374.800 59.800 ;
        RECT 380.400 56.600 381.200 59.800 ;
        RECT 382.000 57.000 382.800 59.800 ;
        RECT 383.600 57.000 384.400 59.800 ;
        RECT 385.200 57.000 386.000 59.800 ;
        RECT 388.400 57.000 389.200 59.800 ;
        RECT 391.600 57.000 392.400 59.800 ;
        RECT 393.200 57.000 394.000 59.800 ;
        RECT 394.800 57.000 395.600 59.800 ;
        RECT 396.400 57.000 397.200 59.800 ;
        RECT 378.600 55.800 381.200 56.600 ;
        RECT 398.000 56.600 398.800 59.800 ;
        RECT 384.600 55.800 389.200 56.400 ;
        RECT 378.600 55.200 379.400 55.800 ;
        RECT 376.400 54.400 379.400 55.200 ;
        RECT 367.700 51.700 371.600 52.300 ;
        RECT 367.700 50.400 368.300 51.700 ;
        RECT 367.600 50.200 368.400 50.400 ;
        RECT 365.400 49.600 366.400 50.200 ;
        RECT 367.000 49.600 368.400 50.200 ;
        RECT 365.400 42.200 366.200 49.600 ;
        RECT 367.000 48.400 367.600 49.600 ;
        RECT 369.200 48.800 370.000 50.400 ;
        RECT 366.800 47.600 367.600 48.400 ;
        RECT 370.800 42.200 371.600 51.700 ;
        RECT 374.000 53.000 382.800 53.800 ;
        RECT 384.600 53.400 385.400 55.800 ;
        RECT 388.400 55.600 389.200 55.800 ;
        RECT 390.000 55.600 391.600 56.400 ;
        RECT 394.600 55.600 395.600 56.400 ;
        RECT 398.000 55.800 400.400 56.600 ;
        RECT 386.800 53.600 387.600 55.200 ;
        RECT 388.400 54.800 389.200 55.000 ;
        RECT 388.400 54.200 392.800 54.800 ;
        RECT 392.000 54.000 392.800 54.200 ;
        RECT 374.000 47.400 374.800 53.000 ;
        RECT 383.400 52.600 385.400 53.400 ;
        RECT 389.200 52.600 392.400 53.400 ;
        RECT 394.800 52.800 395.600 55.600 ;
        RECT 399.600 55.200 400.400 55.800 ;
        RECT 399.600 54.600 401.400 55.200 ;
        RECT 400.600 53.400 401.400 54.600 ;
        RECT 404.400 54.600 405.200 59.800 ;
        RECT 406.000 56.000 406.800 59.800 ;
        RECT 413.000 56.000 413.800 59.000 ;
        RECT 417.200 57.000 418.000 59.000 ;
        RECT 406.000 55.200 407.000 56.000 ;
        RECT 404.400 54.000 405.600 54.600 ;
        RECT 400.600 52.600 404.400 53.400 ;
        RECT 375.400 52.000 376.200 52.200 ;
        RECT 377.200 52.000 378.000 52.400 ;
        RECT 380.400 52.000 381.200 52.400 ;
        RECT 398.000 52.000 398.800 52.600 ;
        RECT 405.000 52.000 405.600 54.000 ;
        RECT 375.400 51.400 398.800 52.000 ;
        RECT 404.800 51.400 405.600 52.000 ;
        RECT 404.800 49.600 405.400 51.400 ;
        RECT 406.200 50.800 407.000 55.200 ;
        RECT 412.200 55.400 413.800 56.000 ;
        RECT 412.200 55.000 413.000 55.400 ;
        RECT 412.200 54.400 412.800 55.000 ;
        RECT 417.400 54.800 418.000 57.000 ;
        RECT 409.200 54.300 410.000 54.400 ;
        RECT 410.800 54.300 412.800 54.400 ;
        RECT 409.200 53.700 412.800 54.300 ;
        RECT 413.800 54.200 418.000 54.800 ;
        RECT 413.800 53.800 414.800 54.200 ;
        RECT 409.200 53.600 410.000 53.700 ;
        RECT 410.800 53.600 412.800 53.700 ;
        RECT 410.800 50.800 411.600 52.400 ;
        RECT 383.600 49.400 384.400 49.600 ;
        RECT 379.000 49.000 384.400 49.400 ;
        RECT 378.200 48.800 384.400 49.000 ;
        RECT 385.400 49.000 394.000 49.600 ;
        RECT 375.600 48.000 377.200 48.800 ;
        RECT 378.200 48.200 379.600 48.800 ;
        RECT 385.400 48.200 386.000 49.000 ;
        RECT 393.200 48.800 394.000 49.000 ;
        RECT 396.400 49.000 405.400 49.600 ;
        RECT 396.400 48.800 397.200 49.000 ;
        RECT 376.600 47.600 377.200 48.000 ;
        RECT 380.200 47.600 386.000 48.200 ;
        RECT 386.600 47.600 389.200 48.400 ;
        RECT 374.000 46.800 376.000 47.400 ;
        RECT 376.600 46.800 380.800 47.600 ;
        RECT 375.400 46.200 376.000 46.800 ;
        RECT 375.400 45.600 376.400 46.200 ;
        RECT 375.600 42.200 376.400 45.600 ;
        RECT 378.800 42.200 379.600 46.800 ;
        RECT 382.000 42.200 382.800 45.000 ;
        RECT 383.600 42.200 384.400 45.000 ;
        RECT 385.200 42.200 386.000 47.000 ;
        RECT 388.400 42.200 389.200 47.000 ;
        RECT 391.600 42.200 392.400 48.400 ;
        RECT 399.600 47.600 402.200 48.400 ;
        RECT 394.800 46.800 399.000 47.600 ;
        RECT 393.200 42.200 394.000 45.000 ;
        RECT 394.800 42.200 395.600 45.000 ;
        RECT 396.400 42.200 397.200 45.000 ;
        RECT 399.600 42.200 400.400 47.600 ;
        RECT 404.800 47.400 405.400 49.000 ;
        RECT 402.800 46.800 405.400 47.400 ;
        RECT 406.000 50.000 407.000 50.800 ;
        RECT 402.800 42.200 403.600 46.800 ;
        RECT 406.000 42.200 406.800 50.000 ;
        RECT 412.200 49.800 412.800 53.600 ;
        RECT 413.400 53.000 414.800 53.800 ;
        RECT 414.200 51.000 414.800 53.000 ;
        RECT 415.600 51.600 416.400 53.200 ;
        RECT 417.200 51.600 418.000 53.200 ;
        RECT 414.200 50.400 418.000 51.000 ;
        RECT 412.200 49.200 413.800 49.800 ;
        RECT 413.000 42.200 413.800 49.200 ;
        RECT 417.400 47.000 418.000 50.400 ;
        RECT 417.200 43.000 418.000 47.000 ;
        RECT 418.800 42.200 419.600 59.800 ;
        RECT 420.400 55.600 421.200 57.200 ;
        RECT 432.200 56.000 433.000 59.000 ;
        RECT 436.400 57.000 437.200 59.000 ;
        RECT 431.400 55.400 433.000 56.000 ;
        RECT 431.400 55.000 432.200 55.400 ;
        RECT 431.400 54.400 432.000 55.000 ;
        RECT 436.600 54.800 437.200 57.000 ;
        RECT 430.000 53.600 432.000 54.400 ;
        RECT 433.000 54.200 437.200 54.800 ;
        RECT 433.000 53.800 434.000 54.200 ;
        RECT 425.200 52.300 426.000 52.400 ;
        RECT 430.000 52.300 430.800 52.400 ;
        RECT 425.200 51.700 430.800 52.300 ;
        RECT 425.200 51.600 426.000 51.700 ;
        RECT 430.000 50.800 430.800 51.700 ;
        RECT 431.400 49.800 432.000 53.600 ;
        RECT 432.600 53.000 434.000 53.800 ;
        RECT 433.400 51.000 434.000 53.000 ;
        RECT 434.800 51.600 435.600 53.200 ;
        RECT 436.400 51.600 437.200 53.200 ;
        RECT 433.400 50.400 437.200 51.000 ;
        RECT 431.400 49.200 433.000 49.800 ;
        RECT 432.200 42.200 433.000 49.200 ;
        RECT 436.600 47.000 437.200 50.400 ;
        RECT 436.400 43.000 437.200 47.000 ;
        RECT 438.000 42.200 438.800 59.800 ;
        RECT 439.600 56.300 440.400 57.200 ;
        RECT 442.800 56.300 443.600 59.800 ;
        RECT 439.600 55.700 443.600 56.300 ;
        RECT 439.600 55.600 440.400 55.700 ;
        RECT 442.600 55.200 443.600 55.700 ;
        RECT 442.600 50.800 443.400 55.200 ;
        RECT 444.400 54.600 445.200 59.800 ;
        RECT 450.800 56.600 451.600 59.800 ;
        RECT 452.400 57.000 453.200 59.800 ;
        RECT 454.000 57.000 454.800 59.800 ;
        RECT 455.600 57.000 456.400 59.800 ;
        RECT 457.200 57.000 458.000 59.800 ;
        RECT 460.400 57.000 461.200 59.800 ;
        RECT 463.600 57.000 464.400 59.800 ;
        RECT 465.200 57.000 466.000 59.800 ;
        RECT 466.800 57.000 467.600 59.800 ;
        RECT 449.200 55.800 451.600 56.600 ;
        RECT 468.400 56.600 469.200 59.800 ;
        RECT 449.200 55.200 450.000 55.800 ;
        RECT 444.000 54.000 445.200 54.600 ;
        RECT 448.200 54.600 450.000 55.200 ;
        RECT 454.000 55.600 455.000 56.400 ;
        RECT 458.000 55.600 459.600 56.400 ;
        RECT 460.400 55.800 465.000 56.400 ;
        RECT 468.400 55.800 471.000 56.600 ;
        RECT 460.400 55.600 461.200 55.800 ;
        RECT 444.000 52.000 444.600 54.000 ;
        RECT 448.200 53.400 449.000 54.600 ;
        RECT 445.200 52.600 449.000 53.400 ;
        RECT 454.000 52.800 454.800 55.600 ;
        RECT 460.400 54.800 461.200 55.000 ;
        RECT 456.800 54.200 461.200 54.800 ;
        RECT 456.800 54.000 457.600 54.200 ;
        RECT 462.000 53.600 462.800 55.200 ;
        RECT 464.200 53.400 465.000 55.800 ;
        RECT 470.200 55.200 471.000 55.800 ;
        RECT 470.200 54.400 473.200 55.200 ;
        RECT 474.800 53.800 475.600 59.800 ;
        RECT 479.000 56.400 479.800 59.800 ;
        RECT 478.000 55.800 479.800 56.400 ;
        RECT 485.000 56.000 485.800 59.000 ;
        RECT 489.200 57.000 490.000 59.000 ;
        RECT 457.200 52.600 460.400 53.400 ;
        RECT 464.200 52.600 466.200 53.400 ;
        RECT 466.800 53.000 475.600 53.800 ;
        RECT 476.400 53.600 477.200 55.200 ;
        RECT 450.800 52.000 451.600 52.600 ;
        RECT 468.400 52.000 469.200 52.400 ;
        RECT 473.200 52.200 474.000 52.400 ;
        RECT 473.200 52.000 474.200 52.200 ;
        RECT 444.000 51.400 444.800 52.000 ;
        RECT 450.800 51.400 474.200 52.000 ;
        RECT 442.600 50.000 443.600 50.800 ;
        RECT 442.800 42.200 443.600 50.000 ;
        RECT 444.200 49.600 444.800 51.400 ;
        RECT 444.200 49.000 453.200 49.600 ;
        RECT 444.200 47.400 444.800 49.000 ;
        RECT 452.400 48.800 453.200 49.000 ;
        RECT 455.600 49.000 464.200 49.600 ;
        RECT 455.600 48.800 456.400 49.000 ;
        RECT 447.400 47.600 450.000 48.400 ;
        RECT 444.200 46.800 446.800 47.400 ;
        RECT 446.000 42.200 446.800 46.800 ;
        RECT 449.200 42.200 450.000 47.600 ;
        RECT 450.600 46.800 454.800 47.600 ;
        RECT 452.400 42.200 453.200 45.000 ;
        RECT 454.000 42.200 454.800 45.000 ;
        RECT 455.600 42.200 456.400 45.000 ;
        RECT 457.200 42.200 458.000 48.400 ;
        RECT 460.400 47.600 463.000 48.400 ;
        RECT 463.600 48.200 464.200 49.000 ;
        RECT 465.200 49.400 466.000 49.600 ;
        RECT 465.200 49.000 470.600 49.400 ;
        RECT 465.200 48.800 471.400 49.000 ;
        RECT 470.000 48.200 471.400 48.800 ;
        RECT 463.600 47.600 469.400 48.200 ;
        RECT 472.400 48.000 474.000 48.800 ;
        RECT 472.400 47.600 473.000 48.000 ;
        RECT 460.400 42.200 461.200 47.000 ;
        RECT 463.600 42.200 464.400 47.000 ;
        RECT 468.800 46.800 473.000 47.600 ;
        RECT 474.800 47.400 475.600 53.000 ;
        RECT 473.600 46.800 475.600 47.400 ;
        RECT 465.200 42.200 466.000 45.000 ;
        RECT 466.800 42.200 467.600 45.000 ;
        RECT 470.000 42.200 470.800 46.800 ;
        RECT 473.600 46.200 474.200 46.800 ;
        RECT 473.200 45.600 474.200 46.200 ;
        RECT 473.200 42.200 474.000 45.600 ;
        RECT 478.000 42.200 478.800 55.800 ;
        RECT 484.200 55.400 485.800 56.000 ;
        RECT 484.200 55.000 485.000 55.400 ;
        RECT 484.200 54.400 484.800 55.000 ;
        RECT 489.400 54.800 490.000 57.000 ;
        RECT 482.800 53.600 484.800 54.400 ;
        RECT 485.800 54.200 490.000 54.800 ;
        RECT 490.800 57.000 491.600 59.000 ;
        RECT 490.800 54.800 491.400 57.000 ;
        RECT 495.000 56.000 495.800 59.000 ;
        RECT 500.400 56.000 501.200 59.800 ;
        RECT 503.600 56.000 504.400 59.800 ;
        RECT 495.000 55.400 496.600 56.000 ;
        RECT 500.400 55.800 504.400 56.000 ;
        RECT 505.200 55.800 506.000 59.800 ;
        RECT 506.800 56.000 507.600 59.800 ;
        RECT 510.000 56.000 510.800 59.800 ;
        RECT 506.800 55.800 510.800 56.000 ;
        RECT 511.600 55.800 512.400 59.800 ;
        RECT 514.800 56.000 515.600 59.800 ;
        RECT 500.600 55.400 504.200 55.800 ;
        RECT 495.800 55.000 496.600 55.400 ;
        RECT 490.800 54.200 495.000 54.800 ;
        RECT 485.800 53.800 486.800 54.200 ;
        RECT 484.200 52.400 484.800 53.600 ;
        RECT 485.400 53.000 486.800 53.800 ;
        RECT 494.000 53.800 495.000 54.200 ;
        RECT 496.000 54.400 496.600 55.000 ;
        RECT 501.200 54.400 502.000 54.800 ;
        RECT 505.200 54.400 505.800 55.800 ;
        RECT 507.000 55.400 510.600 55.800 ;
        RECT 507.600 54.400 508.400 54.800 ;
        RECT 511.600 54.400 512.200 55.800 ;
        RECT 514.600 55.200 515.600 56.000 ;
        RECT 496.000 54.300 498.000 54.400 ;
        RECT 482.800 50.800 483.600 52.400 ;
        RECT 484.200 51.600 485.200 52.400 ;
        RECT 479.600 48.800 480.400 50.400 ;
        RECT 484.200 49.800 484.800 51.600 ;
        RECT 486.200 51.000 486.800 53.000 ;
        RECT 487.600 51.600 488.400 53.200 ;
        RECT 489.200 52.300 490.000 53.200 ;
        RECT 490.800 52.300 491.600 53.200 ;
        RECT 489.200 51.700 491.600 52.300 ;
        RECT 489.200 51.600 490.000 51.700 ;
        RECT 490.800 51.600 491.600 51.700 ;
        RECT 492.400 51.600 493.200 53.200 ;
        RECT 494.000 53.000 495.400 53.800 ;
        RECT 496.000 53.700 499.500 54.300 ;
        RECT 496.000 53.600 498.000 53.700 ;
        RECT 494.000 51.000 494.600 53.000 ;
        RECT 486.200 50.400 490.000 51.000 ;
        RECT 484.200 49.200 485.800 49.800 ;
        RECT 485.000 42.200 485.800 49.200 ;
        RECT 489.400 47.000 490.000 50.400 ;
        RECT 489.200 43.000 490.000 47.000 ;
        RECT 490.800 50.400 494.600 51.000 ;
        RECT 490.800 47.000 491.400 50.400 ;
        RECT 496.000 49.800 496.600 53.600 ;
        RECT 497.200 50.800 498.000 52.400 ;
        RECT 498.900 52.300 499.500 53.700 ;
        RECT 500.400 53.800 502.000 54.400 ;
        RECT 500.400 53.600 501.200 53.800 ;
        RECT 503.400 53.600 506.000 54.400 ;
        RECT 506.800 53.800 508.400 54.400 ;
        RECT 506.800 53.600 507.600 53.800 ;
        RECT 509.800 53.600 512.400 54.400 ;
        RECT 502.000 52.300 502.800 53.200 ;
        RECT 498.900 51.700 502.800 52.300 ;
        RECT 502.000 51.600 502.800 51.700 ;
        RECT 503.400 50.200 504.000 53.600 ;
        RECT 508.400 51.600 509.200 53.200 ;
        RECT 505.200 50.200 506.000 50.400 ;
        RECT 509.800 50.200 510.400 53.600 ;
        RECT 514.600 50.800 515.400 55.200 ;
        RECT 516.400 54.600 517.200 59.800 ;
        RECT 522.800 56.600 523.600 59.800 ;
        RECT 524.400 57.000 525.200 59.800 ;
        RECT 526.000 57.000 526.800 59.800 ;
        RECT 527.600 57.000 528.400 59.800 ;
        RECT 529.200 57.000 530.000 59.800 ;
        RECT 532.400 57.000 533.200 59.800 ;
        RECT 535.600 57.000 536.400 59.800 ;
        RECT 537.200 57.000 538.000 59.800 ;
        RECT 538.800 57.000 539.600 59.800 ;
        RECT 521.200 55.800 523.600 56.600 ;
        RECT 540.400 56.600 541.200 59.800 ;
        RECT 521.200 55.200 522.000 55.800 ;
        RECT 516.000 54.000 517.200 54.600 ;
        RECT 520.200 54.600 522.000 55.200 ;
        RECT 526.000 55.600 527.000 56.400 ;
        RECT 530.000 55.600 531.600 56.400 ;
        RECT 532.400 55.800 537.000 56.400 ;
        RECT 540.400 55.800 543.000 56.600 ;
        RECT 532.400 55.600 533.200 55.800 ;
        RECT 516.000 52.000 516.600 54.000 ;
        RECT 520.200 53.400 521.000 54.600 ;
        RECT 517.200 52.600 521.000 53.400 ;
        RECT 526.000 52.800 526.800 55.600 ;
        RECT 532.400 54.800 533.200 55.000 ;
        RECT 528.800 54.200 533.200 54.800 ;
        RECT 528.800 54.000 529.600 54.200 ;
        RECT 534.000 53.600 534.800 55.200 ;
        RECT 536.200 53.400 537.000 55.800 ;
        RECT 542.200 55.200 543.000 55.800 ;
        RECT 542.200 54.400 545.200 55.200 ;
        RECT 546.800 53.800 547.600 59.800 ;
        RECT 529.200 52.600 532.400 53.400 ;
        RECT 536.200 52.600 538.200 53.400 ;
        RECT 538.800 53.000 547.600 53.800 ;
        RECT 522.800 52.000 523.600 52.600 ;
        RECT 534.000 52.000 534.800 52.400 ;
        RECT 540.400 52.000 541.200 52.400 ;
        RECT 542.000 52.000 542.800 52.400 ;
        RECT 545.400 52.000 546.200 52.200 ;
        RECT 516.000 51.400 516.800 52.000 ;
        RECT 522.800 51.400 546.200 52.000 ;
        RECT 511.600 50.300 512.400 50.400 ;
        RECT 513.200 50.300 514.000 50.400 ;
        RECT 511.600 50.200 514.000 50.300 ;
        RECT 495.000 49.200 496.600 49.800 ;
        RECT 503.000 49.600 504.000 50.200 ;
        RECT 504.600 49.600 506.000 50.200 ;
        RECT 509.400 49.600 510.400 50.200 ;
        RECT 511.000 49.700 514.000 50.200 ;
        RECT 514.600 50.000 515.600 50.800 ;
        RECT 511.000 49.600 512.400 49.700 ;
        RECT 513.200 49.600 514.000 49.700 ;
        RECT 490.800 43.000 491.600 47.000 ;
        RECT 495.000 42.200 495.800 49.200 ;
        RECT 503.000 42.200 503.800 49.600 ;
        RECT 504.600 48.400 505.200 49.600 ;
        RECT 504.400 47.600 505.200 48.400 ;
        RECT 509.400 42.200 510.200 49.600 ;
        RECT 511.000 48.400 511.600 49.600 ;
        RECT 510.800 47.600 511.600 48.400 ;
        RECT 514.800 42.200 515.600 50.000 ;
        RECT 516.200 49.600 516.800 51.400 ;
        RECT 516.200 49.000 525.200 49.600 ;
        RECT 516.200 47.400 516.800 49.000 ;
        RECT 524.400 48.800 525.200 49.000 ;
        RECT 527.600 49.000 536.200 49.600 ;
        RECT 527.600 48.800 528.400 49.000 ;
        RECT 519.400 47.600 522.000 48.400 ;
        RECT 516.200 46.800 518.800 47.400 ;
        RECT 518.000 42.200 518.800 46.800 ;
        RECT 521.200 42.200 522.000 47.600 ;
        RECT 522.600 46.800 526.800 47.600 ;
        RECT 524.400 42.200 525.200 45.000 ;
        RECT 526.000 42.200 526.800 45.000 ;
        RECT 527.600 42.200 528.400 45.000 ;
        RECT 529.200 42.200 530.000 48.400 ;
        RECT 532.400 47.600 535.000 48.400 ;
        RECT 535.600 48.200 536.200 49.000 ;
        RECT 537.200 49.400 538.000 49.600 ;
        RECT 537.200 49.000 542.600 49.400 ;
        RECT 537.200 48.800 543.400 49.000 ;
        RECT 542.000 48.200 543.400 48.800 ;
        RECT 535.600 47.600 541.400 48.200 ;
        RECT 544.400 48.000 546.000 48.800 ;
        RECT 544.400 47.600 545.000 48.000 ;
        RECT 532.400 42.200 533.200 47.000 ;
        RECT 535.600 42.200 536.400 47.000 ;
        RECT 540.800 46.800 545.000 47.600 ;
        RECT 546.800 47.400 547.600 53.000 ;
        RECT 545.600 46.800 547.600 47.400 ;
        RECT 537.200 42.200 538.000 45.000 ;
        RECT 538.800 42.200 539.600 45.000 ;
        RECT 542.000 42.200 542.800 46.800 ;
        RECT 545.600 46.200 546.200 46.800 ;
        RECT 545.200 45.600 546.200 46.200 ;
        RECT 545.200 42.200 546.000 45.600 ;
        RECT 2.800 32.000 3.600 39.800 ;
        RECT 6.000 35.200 6.800 39.800 ;
        RECT 2.600 31.200 3.600 32.000 ;
        RECT 4.200 34.600 6.800 35.200 ;
        RECT 4.200 33.000 4.800 34.600 ;
        RECT 9.200 34.400 10.000 39.800 ;
        RECT 12.400 37.000 13.200 39.800 ;
        RECT 14.000 37.000 14.800 39.800 ;
        RECT 15.600 37.000 16.400 39.800 ;
        RECT 10.600 34.400 14.800 35.200 ;
        RECT 7.400 33.600 10.000 34.400 ;
        RECT 17.200 33.600 18.000 39.800 ;
        RECT 20.400 35.000 21.200 39.800 ;
        RECT 23.600 35.000 24.400 39.800 ;
        RECT 25.200 37.000 26.000 39.800 ;
        RECT 26.800 37.000 27.600 39.800 ;
        RECT 30.000 35.200 30.800 39.800 ;
        RECT 33.200 36.400 34.000 39.800 ;
        RECT 33.200 35.800 34.200 36.400 ;
        RECT 33.600 35.200 34.200 35.800 ;
        RECT 28.800 34.400 33.000 35.200 ;
        RECT 33.600 34.600 35.600 35.200 ;
        RECT 20.400 33.600 23.000 34.400 ;
        RECT 23.600 33.800 29.400 34.400 ;
        RECT 32.400 34.000 33.000 34.400 ;
        RECT 12.400 33.000 13.200 33.200 ;
        RECT 4.200 32.400 13.200 33.000 ;
        RECT 15.600 33.000 16.400 33.200 ;
        RECT 23.600 33.000 24.200 33.800 ;
        RECT 30.000 33.200 31.400 33.800 ;
        RECT 32.400 33.200 34.000 34.000 ;
        RECT 15.600 32.400 24.200 33.000 ;
        RECT 25.200 33.000 31.400 33.200 ;
        RECT 25.200 32.600 30.600 33.000 ;
        RECT 25.200 32.400 26.000 32.600 ;
        RECT 2.600 26.800 3.400 31.200 ;
        RECT 4.200 30.600 4.800 32.400 ;
        RECT 4.000 30.000 4.800 30.600 ;
        RECT 10.800 30.000 34.200 30.600 ;
        RECT 4.000 28.000 4.600 30.000 ;
        RECT 10.800 29.400 11.600 30.000 ;
        RECT 28.400 29.600 29.200 30.000 ;
        RECT 31.600 29.600 32.400 30.000 ;
        RECT 33.400 29.800 34.200 30.000 ;
        RECT 5.200 28.600 9.000 29.400 ;
        RECT 4.000 27.400 5.200 28.000 ;
        RECT 2.600 26.000 3.600 26.800 ;
        RECT 2.800 22.200 3.600 26.000 ;
        RECT 4.400 22.200 5.200 27.400 ;
        RECT 8.200 27.400 9.000 28.600 ;
        RECT 8.200 26.800 10.000 27.400 ;
        RECT 9.200 26.200 10.000 26.800 ;
        RECT 14.000 26.400 14.800 29.200 ;
        RECT 17.200 28.600 20.400 29.400 ;
        RECT 24.200 28.600 26.200 29.400 ;
        RECT 34.800 29.000 35.600 34.600 ;
        RECT 38.000 32.000 38.800 39.800 ;
        RECT 41.200 35.200 42.000 39.800 ;
        RECT 16.800 27.800 17.600 28.000 ;
        RECT 16.800 27.200 21.200 27.800 ;
        RECT 20.400 27.000 21.200 27.200 ;
        RECT 22.000 26.800 22.800 28.400 ;
        RECT 9.200 25.400 11.600 26.200 ;
        RECT 14.000 25.600 15.000 26.400 ;
        RECT 18.000 25.600 19.600 26.400 ;
        RECT 20.400 26.200 21.200 26.400 ;
        RECT 24.200 26.200 25.000 28.600 ;
        RECT 26.800 28.200 35.600 29.000 ;
        RECT 30.200 26.800 33.200 27.600 ;
        RECT 30.200 26.200 31.000 26.800 ;
        RECT 20.400 25.600 25.000 26.200 ;
        RECT 10.800 22.200 11.600 25.400 ;
        RECT 28.400 25.400 31.000 26.200 ;
        RECT 12.400 22.200 13.200 25.000 ;
        RECT 14.000 22.200 14.800 25.000 ;
        RECT 15.600 22.200 16.400 25.000 ;
        RECT 17.200 22.200 18.000 25.000 ;
        RECT 20.400 22.200 21.200 25.000 ;
        RECT 23.600 22.200 24.400 25.000 ;
        RECT 25.200 22.200 26.000 25.000 ;
        RECT 26.800 22.200 27.600 25.000 ;
        RECT 28.400 22.200 29.200 25.400 ;
        RECT 34.800 22.200 35.600 28.200 ;
        RECT 37.800 31.200 38.800 32.000 ;
        RECT 39.400 34.600 42.000 35.200 ;
        RECT 39.400 33.000 40.000 34.600 ;
        RECT 44.400 34.400 45.200 39.800 ;
        RECT 47.600 37.000 48.400 39.800 ;
        RECT 49.200 37.000 50.000 39.800 ;
        RECT 50.800 37.000 51.600 39.800 ;
        RECT 45.800 34.400 50.000 35.200 ;
        RECT 42.600 33.600 45.200 34.400 ;
        RECT 52.400 33.600 53.200 39.800 ;
        RECT 55.600 35.000 56.400 39.800 ;
        RECT 58.800 35.000 59.600 39.800 ;
        RECT 60.400 37.000 61.200 39.800 ;
        RECT 62.000 37.000 62.800 39.800 ;
        RECT 65.200 35.200 66.000 39.800 ;
        RECT 68.400 36.400 69.200 39.800 ;
        RECT 68.400 35.800 69.400 36.400 ;
        RECT 68.800 35.200 69.400 35.800 ;
        RECT 64.000 34.400 68.200 35.200 ;
        RECT 68.800 34.600 70.800 35.200 ;
        RECT 55.600 33.600 58.200 34.400 ;
        RECT 58.800 33.800 64.600 34.400 ;
        RECT 67.600 34.000 68.200 34.400 ;
        RECT 47.600 33.000 48.400 33.200 ;
        RECT 39.400 32.400 48.400 33.000 ;
        RECT 50.800 33.000 51.600 33.200 ;
        RECT 58.800 33.000 59.400 33.800 ;
        RECT 65.200 33.200 66.600 33.800 ;
        RECT 67.600 33.200 69.200 34.000 ;
        RECT 50.800 32.400 59.400 33.000 ;
        RECT 60.400 33.000 66.600 33.200 ;
        RECT 60.400 32.600 65.800 33.000 ;
        RECT 60.400 32.400 61.200 32.600 ;
        RECT 37.800 26.800 38.600 31.200 ;
        RECT 39.400 30.600 40.000 32.400 ;
        RECT 39.200 30.000 40.000 30.600 ;
        RECT 46.000 30.000 69.400 30.600 ;
        RECT 39.200 28.000 39.800 30.000 ;
        RECT 46.000 29.400 46.800 30.000 ;
        RECT 63.600 29.600 64.400 30.000 ;
        RECT 66.800 29.600 67.600 30.000 ;
        RECT 68.600 29.800 69.400 30.000 ;
        RECT 40.400 28.600 44.200 29.400 ;
        RECT 39.200 27.400 40.400 28.000 ;
        RECT 37.800 26.000 38.800 26.800 ;
        RECT 38.000 22.200 38.800 26.000 ;
        RECT 39.600 22.200 40.400 27.400 ;
        RECT 43.400 27.400 44.200 28.600 ;
        RECT 43.400 26.800 45.200 27.400 ;
        RECT 44.400 26.200 45.200 26.800 ;
        RECT 49.200 26.400 50.000 29.200 ;
        RECT 52.400 28.600 55.600 29.400 ;
        RECT 59.400 28.600 61.400 29.400 ;
        RECT 70.000 29.000 70.800 34.600 ;
        RECT 74.800 32.400 75.600 39.800 ;
        RECT 73.400 31.800 75.600 32.400 ;
        RECT 73.400 31.200 74.000 31.800 ;
        RECT 72.800 30.400 74.000 31.200 ;
        RECT 78.000 31.200 78.800 39.800 ;
        RECT 81.200 31.200 82.000 39.800 ;
        RECT 84.400 31.200 85.200 39.800 ;
        RECT 87.600 31.200 88.400 39.800 ;
        RECT 92.400 36.400 93.200 39.800 ;
        RECT 92.200 35.800 93.200 36.400 ;
        RECT 92.200 35.200 92.800 35.800 ;
        RECT 95.600 35.200 96.400 39.800 ;
        RECT 98.800 37.000 99.600 39.800 ;
        RECT 100.400 37.000 101.200 39.800 ;
        RECT 90.800 34.600 92.800 35.200 ;
        RECT 78.000 30.400 79.800 31.200 ;
        RECT 81.200 30.400 83.400 31.200 ;
        RECT 84.400 30.400 86.600 31.200 ;
        RECT 87.600 30.400 90.000 31.200 ;
        RECT 52.000 27.800 52.800 28.000 ;
        RECT 52.000 27.200 56.400 27.800 ;
        RECT 55.600 27.000 56.400 27.200 ;
        RECT 57.200 26.800 58.000 28.400 ;
        RECT 44.400 25.400 46.800 26.200 ;
        RECT 49.200 25.600 50.200 26.400 ;
        RECT 53.200 25.600 54.800 26.400 ;
        RECT 55.600 26.200 56.400 26.400 ;
        RECT 59.400 26.200 60.200 28.600 ;
        RECT 62.000 28.200 70.800 29.000 ;
        RECT 65.400 26.800 68.400 27.600 ;
        RECT 65.400 26.200 66.200 26.800 ;
        RECT 55.600 25.600 60.200 26.200 ;
        RECT 46.000 22.200 46.800 25.400 ;
        RECT 63.600 25.400 66.200 26.200 ;
        RECT 47.600 22.200 48.400 25.000 ;
        RECT 49.200 22.200 50.000 25.000 ;
        RECT 50.800 22.200 51.600 25.000 ;
        RECT 52.400 22.200 53.200 25.000 ;
        RECT 55.600 22.200 56.400 25.000 ;
        RECT 58.800 22.200 59.600 25.000 ;
        RECT 60.400 22.200 61.200 25.000 ;
        RECT 62.000 22.200 62.800 25.000 ;
        RECT 63.600 22.200 64.400 25.400 ;
        RECT 70.000 22.200 70.800 28.200 ;
        RECT 73.400 27.400 74.000 30.400 ;
        RECT 74.800 28.800 75.600 30.400 ;
        RECT 79.000 29.000 79.800 30.400 ;
        RECT 82.600 29.000 83.400 30.400 ;
        RECT 85.800 29.000 86.600 30.400 ;
        RECT 79.000 28.200 81.600 29.000 ;
        RECT 82.600 28.200 85.000 29.000 ;
        RECT 85.800 28.200 88.400 29.000 ;
        RECT 79.000 27.600 79.800 28.200 ;
        RECT 82.600 27.600 83.400 28.200 ;
        RECT 85.800 27.600 86.600 28.200 ;
        RECT 89.200 27.600 90.000 30.400 ;
        RECT 73.400 26.800 75.600 27.400 ;
        RECT 74.800 22.200 75.600 26.800 ;
        RECT 78.000 26.800 79.800 27.600 ;
        RECT 81.200 26.800 83.400 27.600 ;
        RECT 84.400 26.800 86.600 27.600 ;
        RECT 87.600 26.800 90.000 27.600 ;
        RECT 90.800 29.000 91.600 34.600 ;
        RECT 93.400 34.400 97.600 35.200 ;
        RECT 102.000 35.000 102.800 39.800 ;
        RECT 105.200 35.000 106.000 39.800 ;
        RECT 93.400 34.000 94.000 34.400 ;
        RECT 92.400 33.200 94.000 34.000 ;
        RECT 97.000 33.800 102.800 34.400 ;
        RECT 95.000 33.200 96.400 33.800 ;
        RECT 95.000 33.000 101.200 33.200 ;
        RECT 95.800 32.600 101.200 33.000 ;
        RECT 100.400 32.400 101.200 32.600 ;
        RECT 102.200 33.000 102.800 33.800 ;
        RECT 103.400 33.600 106.000 34.400 ;
        RECT 108.400 33.600 109.200 39.800 ;
        RECT 110.000 37.000 110.800 39.800 ;
        RECT 111.600 37.000 112.400 39.800 ;
        RECT 113.200 37.000 114.000 39.800 ;
        RECT 111.600 34.400 115.800 35.200 ;
        RECT 116.400 34.400 117.200 39.800 ;
        RECT 119.600 35.200 120.400 39.800 ;
        RECT 119.600 34.600 122.200 35.200 ;
        RECT 116.400 33.600 119.000 34.400 ;
        RECT 110.000 33.000 110.800 33.200 ;
        RECT 102.200 32.400 110.800 33.000 ;
        RECT 113.200 33.000 114.000 33.200 ;
        RECT 121.600 33.000 122.200 34.600 ;
        RECT 113.200 32.400 122.200 33.000 ;
        RECT 121.600 30.600 122.200 32.400 ;
        RECT 122.800 32.000 123.600 39.800 ;
        RECT 134.000 32.000 134.800 39.800 ;
        RECT 137.200 35.200 138.000 39.800 ;
        RECT 122.800 31.200 123.800 32.000 ;
        RECT 92.200 30.000 115.600 30.600 ;
        RECT 121.600 30.000 122.400 30.600 ;
        RECT 92.200 29.800 93.000 30.000 ;
        RECT 94.000 29.600 94.800 30.000 ;
        RECT 97.200 29.600 98.000 30.000 ;
        RECT 114.800 29.400 115.600 30.000 ;
        RECT 90.800 28.200 99.600 29.000 ;
        RECT 100.200 28.600 102.200 29.400 ;
        RECT 106.000 28.600 109.200 29.400 ;
        RECT 78.000 22.200 78.800 26.800 ;
        RECT 81.200 22.200 82.000 26.800 ;
        RECT 84.400 22.200 85.200 26.800 ;
        RECT 87.600 22.200 88.400 26.800 ;
        RECT 90.800 22.200 91.600 28.200 ;
        RECT 93.200 26.800 96.200 27.600 ;
        RECT 95.400 26.200 96.200 26.800 ;
        RECT 101.400 26.200 102.200 28.600 ;
        RECT 103.600 26.800 104.400 28.400 ;
        RECT 108.800 27.800 109.600 28.000 ;
        RECT 105.200 27.200 109.600 27.800 ;
        RECT 105.200 27.000 106.000 27.200 ;
        RECT 111.600 26.400 112.400 29.200 ;
        RECT 117.400 28.600 121.200 29.400 ;
        RECT 117.400 27.400 118.200 28.600 ;
        RECT 121.800 28.000 122.400 30.000 ;
        RECT 105.200 26.200 106.000 26.400 ;
        RECT 95.400 25.400 98.000 26.200 ;
        RECT 101.400 25.600 106.000 26.200 ;
        RECT 106.800 25.600 108.400 26.400 ;
        RECT 111.400 25.600 112.400 26.400 ;
        RECT 116.400 26.800 118.200 27.400 ;
        RECT 121.200 27.400 122.400 28.000 ;
        RECT 116.400 26.200 117.200 26.800 ;
        RECT 97.200 22.200 98.000 25.400 ;
        RECT 114.800 25.400 117.200 26.200 ;
        RECT 98.800 22.200 99.600 25.000 ;
        RECT 100.400 22.200 101.200 25.000 ;
        RECT 102.000 22.200 102.800 25.000 ;
        RECT 105.200 22.200 106.000 25.000 ;
        RECT 108.400 22.200 109.200 25.000 ;
        RECT 110.000 22.200 110.800 25.000 ;
        RECT 111.600 22.200 112.400 25.000 ;
        RECT 113.200 22.200 114.000 25.000 ;
        RECT 114.800 22.200 115.600 25.400 ;
        RECT 121.200 22.200 122.000 27.400 ;
        RECT 123.000 26.800 123.800 31.200 ;
        RECT 122.800 26.000 123.800 26.800 ;
        RECT 133.800 31.200 134.800 32.000 ;
        RECT 135.400 34.600 138.000 35.200 ;
        RECT 135.400 33.000 136.000 34.600 ;
        RECT 140.400 34.400 141.200 39.800 ;
        RECT 143.600 37.000 144.400 39.800 ;
        RECT 145.200 37.000 146.000 39.800 ;
        RECT 146.800 37.000 147.600 39.800 ;
        RECT 141.800 34.400 146.000 35.200 ;
        RECT 138.600 33.600 141.200 34.400 ;
        RECT 148.400 33.600 149.200 39.800 ;
        RECT 151.600 35.000 152.400 39.800 ;
        RECT 154.800 35.000 155.600 39.800 ;
        RECT 156.400 37.000 157.200 39.800 ;
        RECT 158.000 37.000 158.800 39.800 ;
        RECT 161.200 35.200 162.000 39.800 ;
        RECT 164.400 36.400 165.200 39.800 ;
        RECT 164.400 35.800 165.400 36.400 ;
        RECT 164.800 35.200 165.400 35.800 ;
        RECT 160.000 34.400 164.200 35.200 ;
        RECT 164.800 34.600 166.800 35.200 ;
        RECT 151.600 33.600 154.200 34.400 ;
        RECT 154.800 33.800 160.600 34.400 ;
        RECT 163.600 34.000 164.200 34.400 ;
        RECT 143.600 33.000 144.400 33.200 ;
        RECT 135.400 32.400 144.400 33.000 ;
        RECT 146.800 33.000 147.600 33.200 ;
        RECT 154.800 33.000 155.400 33.800 ;
        RECT 161.200 33.200 162.600 33.800 ;
        RECT 163.600 33.200 165.200 34.000 ;
        RECT 146.800 32.400 155.400 33.000 ;
        RECT 156.400 33.000 162.600 33.200 ;
        RECT 156.400 32.600 161.800 33.000 ;
        RECT 156.400 32.400 157.200 32.600 ;
        RECT 133.800 26.800 134.600 31.200 ;
        RECT 135.400 30.600 136.000 32.400 ;
        RECT 159.400 31.800 160.200 32.000 ;
        RECT 162.800 31.800 163.600 32.400 ;
        RECT 136.600 31.200 163.600 31.800 ;
        RECT 136.600 31.000 137.400 31.200 ;
        RECT 135.200 30.000 136.000 30.600 ;
        RECT 135.200 28.000 135.800 30.000 ;
        RECT 136.400 28.600 140.200 29.400 ;
        RECT 135.200 27.400 136.400 28.000 ;
        RECT 133.800 26.000 134.800 26.800 ;
        RECT 122.800 22.200 123.600 26.000 ;
        RECT 134.000 22.200 134.800 26.000 ;
        RECT 135.600 22.200 136.400 27.400 ;
        RECT 139.400 27.400 140.200 28.600 ;
        RECT 139.400 26.800 141.200 27.400 ;
        RECT 140.400 26.200 141.200 26.800 ;
        RECT 145.200 26.400 146.000 29.200 ;
        RECT 148.400 28.600 151.600 29.400 ;
        RECT 155.400 28.600 157.400 29.400 ;
        RECT 166.000 29.000 166.800 34.600 ;
        RECT 169.200 32.000 170.000 39.800 ;
        RECT 172.400 35.200 173.200 39.800 ;
        RECT 148.000 27.800 148.800 28.000 ;
        RECT 148.000 27.200 152.400 27.800 ;
        RECT 151.600 27.000 152.400 27.200 ;
        RECT 153.200 26.800 154.000 28.400 ;
        RECT 140.400 25.400 142.800 26.200 ;
        RECT 145.200 25.600 146.200 26.400 ;
        RECT 149.200 25.600 150.800 26.400 ;
        RECT 151.600 26.200 152.400 26.400 ;
        RECT 155.400 26.200 156.200 28.600 ;
        RECT 158.000 28.200 166.800 29.000 ;
        RECT 161.400 26.800 164.400 27.600 ;
        RECT 161.400 26.200 162.200 26.800 ;
        RECT 151.600 25.600 156.200 26.200 ;
        RECT 142.000 22.200 142.800 25.400 ;
        RECT 159.600 25.400 162.200 26.200 ;
        RECT 143.600 22.200 144.400 25.000 ;
        RECT 145.200 22.200 146.000 25.000 ;
        RECT 146.800 22.200 147.600 25.000 ;
        RECT 148.400 22.200 149.200 25.000 ;
        RECT 151.600 22.200 152.400 25.000 ;
        RECT 154.800 22.200 155.600 25.000 ;
        RECT 156.400 22.200 157.200 25.000 ;
        RECT 158.000 22.200 158.800 25.000 ;
        RECT 159.600 22.200 160.400 25.400 ;
        RECT 166.000 22.200 166.800 28.200 ;
        RECT 169.000 31.200 170.000 32.000 ;
        RECT 170.600 34.600 173.200 35.200 ;
        RECT 170.600 33.000 171.200 34.600 ;
        RECT 175.600 34.400 176.400 39.800 ;
        RECT 178.800 37.000 179.600 39.800 ;
        RECT 180.400 37.000 181.200 39.800 ;
        RECT 182.000 37.000 182.800 39.800 ;
        RECT 177.000 34.400 181.200 35.200 ;
        RECT 173.800 33.600 176.400 34.400 ;
        RECT 183.600 33.600 184.400 39.800 ;
        RECT 186.800 35.000 187.600 39.800 ;
        RECT 190.000 35.000 190.800 39.800 ;
        RECT 191.600 37.000 192.400 39.800 ;
        RECT 193.200 37.000 194.000 39.800 ;
        RECT 196.400 35.200 197.200 39.800 ;
        RECT 199.600 36.400 200.400 39.800 ;
        RECT 199.600 35.800 200.600 36.400 ;
        RECT 200.000 35.200 200.600 35.800 ;
        RECT 195.200 34.400 199.400 35.200 ;
        RECT 200.000 34.600 202.000 35.200 ;
        RECT 186.800 33.600 189.400 34.400 ;
        RECT 190.000 33.800 195.800 34.400 ;
        RECT 198.800 34.000 199.400 34.400 ;
        RECT 178.800 33.000 179.600 33.200 ;
        RECT 170.600 32.400 179.600 33.000 ;
        RECT 182.000 33.000 182.800 33.200 ;
        RECT 190.000 33.000 190.600 33.800 ;
        RECT 196.400 33.200 197.800 33.800 ;
        RECT 198.800 33.200 200.400 34.000 ;
        RECT 182.000 32.400 190.600 33.000 ;
        RECT 191.600 33.000 197.800 33.200 ;
        RECT 191.600 32.600 197.000 33.000 ;
        RECT 191.600 32.400 192.400 32.600 ;
        RECT 169.000 26.800 169.800 31.200 ;
        RECT 170.600 30.600 171.200 32.400 ;
        RECT 194.600 31.800 195.600 32.000 ;
        RECT 198.000 31.800 198.800 32.400 ;
        RECT 171.800 31.200 198.800 31.800 ;
        RECT 171.800 31.000 172.600 31.200 ;
        RECT 170.400 30.000 171.200 30.600 ;
        RECT 170.400 28.000 171.000 30.000 ;
        RECT 171.600 28.600 175.400 29.400 ;
        RECT 170.400 27.400 171.600 28.000 ;
        RECT 169.000 26.000 170.000 26.800 ;
        RECT 169.200 22.200 170.000 26.000 ;
        RECT 170.800 22.200 171.600 27.400 ;
        RECT 174.600 27.400 175.400 28.600 ;
        RECT 174.600 26.800 176.400 27.400 ;
        RECT 175.600 26.200 176.400 26.800 ;
        RECT 180.400 26.400 181.200 29.200 ;
        RECT 183.600 28.600 186.800 29.400 ;
        RECT 190.600 28.600 192.600 29.400 ;
        RECT 201.200 29.000 202.000 34.600 ;
        RECT 183.200 27.800 184.000 28.000 ;
        RECT 183.200 27.200 187.600 27.800 ;
        RECT 186.800 27.000 187.600 27.200 ;
        RECT 188.400 26.800 189.200 28.400 ;
        RECT 175.600 25.400 178.000 26.200 ;
        RECT 180.400 25.600 181.400 26.400 ;
        RECT 184.400 25.600 186.000 26.400 ;
        RECT 186.800 26.200 187.600 26.400 ;
        RECT 190.600 26.200 191.400 28.600 ;
        RECT 193.200 28.200 202.000 29.000 ;
        RECT 196.600 26.800 199.600 27.600 ;
        RECT 196.600 26.200 197.400 26.800 ;
        RECT 186.800 25.600 191.400 26.200 ;
        RECT 177.200 22.200 178.000 25.400 ;
        RECT 194.800 25.400 197.400 26.200 ;
        RECT 178.800 22.200 179.600 25.000 ;
        RECT 180.400 22.200 181.200 25.000 ;
        RECT 182.000 22.200 182.800 25.000 ;
        RECT 183.600 22.200 184.400 25.000 ;
        RECT 186.800 22.200 187.600 25.000 ;
        RECT 190.000 22.200 190.800 25.000 ;
        RECT 191.600 22.200 192.400 25.000 ;
        RECT 193.200 22.200 194.000 25.000 ;
        RECT 194.800 22.200 195.600 25.400 ;
        RECT 201.200 22.200 202.000 28.200 ;
        RECT 202.800 26.800 203.600 28.400 ;
        RECT 204.400 26.200 205.200 39.800 ;
        RECT 208.400 33.600 209.200 34.400 ;
        RECT 206.000 31.600 206.800 33.200 ;
        RECT 208.400 32.400 209.000 33.600 ;
        RECT 209.800 32.400 210.600 39.800 ;
        RECT 214.000 34.300 214.800 34.400 ;
        RECT 215.600 34.300 216.400 39.800 ;
        RECT 214.000 33.700 216.400 34.300 ;
        RECT 214.000 33.600 214.800 33.700 ;
        RECT 207.600 31.800 209.000 32.400 ;
        RECT 209.600 31.800 210.600 32.400 ;
        RECT 207.600 31.600 208.400 31.800 ;
        RECT 206.100 30.300 206.700 31.600 ;
        RECT 209.600 30.300 210.200 31.800 ;
        RECT 206.100 29.700 210.200 30.300 ;
        RECT 209.600 28.400 210.200 29.700 ;
        RECT 210.800 30.300 211.600 30.400 ;
        RECT 214.000 30.300 214.800 30.400 ;
        RECT 210.800 29.700 214.800 30.300 ;
        RECT 210.800 28.800 211.600 29.700 ;
        RECT 214.000 29.600 214.800 29.700 ;
        RECT 215.600 30.300 216.400 33.700 ;
        RECT 219.800 32.400 220.600 39.800 ;
        RECT 226.200 38.400 227.000 39.800 ;
        RECT 225.200 37.600 227.000 38.400 ;
        RECT 221.200 33.600 222.000 34.400 ;
        RECT 221.400 32.400 222.000 33.600 ;
        RECT 226.200 32.400 227.000 37.600 ;
        RECT 227.600 33.600 228.400 34.400 ;
        RECT 227.800 32.400 228.400 33.600 ;
        RECT 218.800 31.600 220.800 32.400 ;
        RECT 221.400 31.800 222.800 32.400 ;
        RECT 226.200 31.800 227.200 32.400 ;
        RECT 227.800 32.300 229.200 32.400 ;
        RECT 230.000 32.300 230.800 32.400 ;
        RECT 227.800 31.800 230.800 32.300 ;
        RECT 231.600 32.000 232.400 39.800 ;
        RECT 234.800 35.200 235.600 39.800 ;
        RECT 222.000 31.600 222.800 31.800 ;
        RECT 218.800 30.300 219.600 30.400 ;
        RECT 215.600 29.700 219.600 30.300 ;
        RECT 207.600 27.600 210.200 28.400 ;
        RECT 212.400 28.200 213.200 28.400 ;
        RECT 211.600 27.600 213.200 28.200 ;
        RECT 207.800 26.200 208.400 27.600 ;
        RECT 211.600 27.200 212.400 27.600 ;
        RECT 209.400 26.200 213.000 26.600 ;
        RECT 204.400 25.600 206.200 26.200 ;
        RECT 205.400 22.200 206.200 25.600 ;
        RECT 207.600 22.200 208.400 26.200 ;
        RECT 209.200 26.000 213.200 26.200 ;
        RECT 209.200 22.200 210.000 26.000 ;
        RECT 212.400 22.200 213.200 26.000 ;
        RECT 214.000 24.800 214.800 26.400 ;
        RECT 215.600 22.200 216.400 29.700 ;
        RECT 218.800 28.800 219.600 29.700 ;
        RECT 220.200 28.400 220.800 31.600 ;
        RECT 222.000 30.300 222.800 30.400 ;
        RECT 225.200 30.300 226.000 30.400 ;
        RECT 222.000 29.700 226.000 30.300 ;
        RECT 222.000 29.600 222.800 29.700 ;
        RECT 225.200 28.800 226.000 29.700 ;
        RECT 226.600 28.400 227.200 31.800 ;
        RECT 228.400 31.700 230.800 31.800 ;
        RECT 228.400 31.600 229.200 31.700 ;
        RECT 230.000 31.600 230.800 31.700 ;
        RECT 231.400 31.200 232.400 32.000 ;
        RECT 233.000 34.600 235.600 35.200 ;
        RECT 233.000 33.000 233.600 34.600 ;
        RECT 238.000 34.400 238.800 39.800 ;
        RECT 241.200 37.000 242.000 39.800 ;
        RECT 242.800 37.000 243.600 39.800 ;
        RECT 244.400 37.000 245.200 39.800 ;
        RECT 239.400 34.400 243.600 35.200 ;
        RECT 236.200 33.600 238.800 34.400 ;
        RECT 246.000 33.600 246.800 39.800 ;
        RECT 249.200 35.000 250.000 39.800 ;
        RECT 252.400 35.000 253.200 39.800 ;
        RECT 254.000 37.000 254.800 39.800 ;
        RECT 255.600 37.000 256.400 39.800 ;
        RECT 258.800 35.200 259.600 39.800 ;
        RECT 262.000 36.400 262.800 39.800 ;
        RECT 262.000 35.800 263.000 36.400 ;
        RECT 262.400 35.200 263.000 35.800 ;
        RECT 257.600 34.400 261.800 35.200 ;
        RECT 262.400 34.600 264.400 35.200 ;
        RECT 249.200 33.600 251.800 34.400 ;
        RECT 252.400 33.800 258.200 34.400 ;
        RECT 261.200 34.000 261.800 34.400 ;
        RECT 241.200 33.000 242.000 33.200 ;
        RECT 233.000 32.400 242.000 33.000 ;
        RECT 244.400 33.000 245.200 33.200 ;
        RECT 252.400 33.000 253.000 33.800 ;
        RECT 258.800 33.200 260.200 33.800 ;
        RECT 261.200 33.200 262.800 34.000 ;
        RECT 244.400 32.400 253.000 33.000 ;
        RECT 254.000 33.000 260.200 33.200 ;
        RECT 254.000 32.600 259.400 33.000 ;
        RECT 254.000 32.400 254.800 32.600 ;
        RECT 217.200 28.200 218.000 28.400 ;
        RECT 217.200 27.600 218.800 28.200 ;
        RECT 220.200 27.600 222.800 28.400 ;
        RECT 223.600 28.200 224.400 28.400 ;
        RECT 223.600 27.600 225.200 28.200 ;
        RECT 226.600 27.600 229.200 28.400 ;
        RECT 218.000 27.200 218.800 27.600 ;
        RECT 217.400 26.200 221.000 26.600 ;
        RECT 222.000 26.200 222.600 27.600 ;
        RECT 224.400 27.200 225.200 27.600 ;
        RECT 223.800 26.200 227.400 26.600 ;
        RECT 228.400 26.200 229.000 27.600 ;
        RECT 231.400 26.800 232.200 31.200 ;
        RECT 233.000 30.600 233.600 32.400 ;
        RECT 260.400 32.300 261.200 32.400 ;
        RECT 262.000 32.300 262.800 32.400 ;
        RECT 257.000 31.800 257.800 32.000 ;
        RECT 260.400 31.800 262.800 32.300 ;
        RECT 234.200 31.700 262.800 31.800 ;
        RECT 234.200 31.200 261.200 31.700 ;
        RECT 262.000 31.600 262.800 31.700 ;
        RECT 234.200 31.000 235.000 31.200 ;
        RECT 232.800 30.000 233.600 30.600 ;
        RECT 232.800 28.000 233.400 30.000 ;
        RECT 234.000 28.600 237.800 29.400 ;
        RECT 232.800 27.400 234.000 28.000 ;
        RECT 217.200 26.000 221.200 26.200 ;
        RECT 217.200 22.200 218.000 26.000 ;
        RECT 220.400 22.200 221.200 26.000 ;
        RECT 222.000 22.200 222.800 26.200 ;
        RECT 223.600 26.000 227.600 26.200 ;
        RECT 223.600 22.200 224.400 26.000 ;
        RECT 226.800 22.200 227.600 26.000 ;
        RECT 228.400 22.200 229.200 26.200 ;
        RECT 231.400 26.000 232.400 26.800 ;
        RECT 231.600 22.200 232.400 26.000 ;
        RECT 233.200 22.200 234.000 27.400 ;
        RECT 237.000 27.400 237.800 28.600 ;
        RECT 237.000 26.800 238.800 27.400 ;
        RECT 238.000 26.200 238.800 26.800 ;
        RECT 242.800 26.400 243.600 29.200 ;
        RECT 246.000 28.600 249.200 29.400 ;
        RECT 253.000 28.600 255.000 29.400 ;
        RECT 263.600 29.000 264.400 34.600 ;
        RECT 245.600 27.800 246.400 28.000 ;
        RECT 245.600 27.200 250.000 27.800 ;
        RECT 249.200 27.000 250.000 27.200 ;
        RECT 250.800 26.800 251.600 28.400 ;
        RECT 238.000 25.400 240.400 26.200 ;
        RECT 242.800 25.600 243.800 26.400 ;
        RECT 246.800 25.600 248.400 26.400 ;
        RECT 249.200 26.200 250.000 26.400 ;
        RECT 253.000 26.200 253.800 28.600 ;
        RECT 255.600 28.200 264.400 29.000 ;
        RECT 259.000 26.800 262.000 27.600 ;
        RECT 259.000 26.200 259.800 26.800 ;
        RECT 249.200 25.600 253.800 26.200 ;
        RECT 239.600 22.200 240.400 25.400 ;
        RECT 257.200 25.400 259.800 26.200 ;
        RECT 241.200 22.200 242.000 25.000 ;
        RECT 242.800 22.200 243.600 25.000 ;
        RECT 244.400 22.200 245.200 25.000 ;
        RECT 246.000 22.200 246.800 25.000 ;
        RECT 249.200 22.200 250.000 25.000 ;
        RECT 252.400 22.200 253.200 25.000 ;
        RECT 254.000 22.200 254.800 25.000 ;
        RECT 255.600 22.200 256.400 25.000 ;
        RECT 257.200 22.200 258.000 25.400 ;
        RECT 263.600 22.200 264.400 28.200 ;
        RECT 266.800 28.300 267.600 39.800 ;
        RECT 271.000 32.400 271.800 39.800 ;
        RECT 272.400 33.600 273.200 34.400 ;
        RECT 272.600 32.400 273.200 33.600 ;
        RECT 282.000 33.600 282.800 34.400 ;
        RECT 282.000 32.400 282.600 33.600 ;
        RECT 283.400 32.400 284.200 39.800 ;
        RECT 271.000 31.800 272.000 32.400 ;
        RECT 272.600 31.800 274.000 32.400 ;
        RECT 270.000 28.800 270.800 30.400 ;
        RECT 271.400 28.400 272.000 31.800 ;
        RECT 273.200 31.600 274.000 31.800 ;
        RECT 281.200 31.800 282.600 32.400 ;
        RECT 283.200 31.800 284.200 32.400 ;
        RECT 289.200 32.000 290.000 39.800 ;
        RECT 292.400 35.200 293.200 39.800 ;
        RECT 281.200 31.600 282.000 31.800 ;
        RECT 273.300 30.300 273.900 31.600 ;
        RECT 283.200 30.300 283.800 31.800 ;
        RECT 289.000 31.200 290.000 32.000 ;
        RECT 290.600 34.600 293.200 35.200 ;
        RECT 290.600 33.000 291.200 34.600 ;
        RECT 295.600 34.400 296.400 39.800 ;
        RECT 298.800 37.000 299.600 39.800 ;
        RECT 300.400 37.000 301.200 39.800 ;
        RECT 302.000 37.000 302.800 39.800 ;
        RECT 297.000 34.400 301.200 35.200 ;
        RECT 293.800 33.600 296.400 34.400 ;
        RECT 303.600 33.600 304.400 39.800 ;
        RECT 306.800 35.000 307.600 39.800 ;
        RECT 310.000 35.000 310.800 39.800 ;
        RECT 311.600 37.000 312.400 39.800 ;
        RECT 313.200 37.000 314.000 39.800 ;
        RECT 316.400 35.200 317.200 39.800 ;
        RECT 319.600 36.400 320.400 39.800 ;
        RECT 319.600 35.800 320.600 36.400 ;
        RECT 320.000 35.200 320.600 35.800 ;
        RECT 315.200 34.400 319.400 35.200 ;
        RECT 320.000 34.600 322.000 35.200 ;
        RECT 306.800 33.600 309.400 34.400 ;
        RECT 310.000 33.800 315.800 34.400 ;
        RECT 318.800 34.000 319.400 34.400 ;
        RECT 298.800 33.000 299.600 33.200 ;
        RECT 290.600 32.400 299.600 33.000 ;
        RECT 302.000 33.000 302.800 33.200 ;
        RECT 310.000 33.000 310.600 33.800 ;
        RECT 316.400 33.200 317.800 33.800 ;
        RECT 318.800 33.200 320.400 34.000 ;
        RECT 302.000 32.400 310.600 33.000 ;
        RECT 311.600 33.000 317.800 33.200 ;
        RECT 311.600 32.600 317.000 33.000 ;
        RECT 311.600 32.400 312.400 32.600 ;
        RECT 273.300 29.700 283.800 30.300 ;
        RECT 283.200 28.400 283.800 29.700 ;
        RECT 284.400 30.300 285.200 30.400 ;
        RECT 287.600 30.300 288.400 30.400 ;
        RECT 284.400 29.700 288.400 30.300 ;
        RECT 284.400 28.800 285.200 29.700 ;
        RECT 287.600 29.600 288.400 29.700 ;
        RECT 268.400 28.300 269.200 28.400 ;
        RECT 266.800 28.200 269.200 28.300 ;
        RECT 266.800 27.700 270.000 28.200 ;
        RECT 265.200 24.800 266.000 26.400 ;
        RECT 266.800 22.200 267.600 27.700 ;
        RECT 268.400 27.600 270.000 27.700 ;
        RECT 271.400 27.600 274.000 28.400 ;
        RECT 281.200 27.600 283.800 28.400 ;
        RECT 286.000 28.200 286.800 28.400 ;
        RECT 285.200 27.600 286.800 28.200 ;
        RECT 269.200 27.200 270.000 27.600 ;
        RECT 268.600 26.200 272.200 26.600 ;
        RECT 273.200 26.200 273.800 27.600 ;
        RECT 281.400 26.200 282.000 27.600 ;
        RECT 285.200 27.200 286.000 27.600 ;
        RECT 289.000 26.800 289.800 31.200 ;
        RECT 290.600 30.600 291.200 32.400 ;
        RECT 314.600 31.800 315.600 32.000 ;
        RECT 318.000 31.800 318.800 32.400 ;
        RECT 291.800 31.200 318.800 31.800 ;
        RECT 291.800 31.000 292.600 31.200 ;
        RECT 290.400 30.000 291.200 30.600 ;
        RECT 290.400 28.000 291.000 30.000 ;
        RECT 291.600 28.600 295.400 29.400 ;
        RECT 290.400 27.400 291.600 28.000 ;
        RECT 283.000 26.200 286.600 26.600 ;
        RECT 268.400 26.000 272.400 26.200 ;
        RECT 268.400 22.200 269.200 26.000 ;
        RECT 271.600 22.200 272.400 26.000 ;
        RECT 273.200 22.200 274.000 26.200 ;
        RECT 281.200 22.200 282.000 26.200 ;
        RECT 282.800 26.000 286.800 26.200 ;
        RECT 289.000 26.000 290.000 26.800 ;
        RECT 282.800 22.200 283.600 26.000 ;
        RECT 286.000 22.200 286.800 26.000 ;
        RECT 289.200 22.200 290.000 26.000 ;
        RECT 290.800 22.200 291.600 27.400 ;
        RECT 294.600 27.400 295.400 28.600 ;
        RECT 294.600 26.800 296.400 27.400 ;
        RECT 295.600 26.200 296.400 26.800 ;
        RECT 300.400 26.400 301.200 29.200 ;
        RECT 303.600 28.600 306.800 29.400 ;
        RECT 310.600 28.600 312.600 29.400 ;
        RECT 321.200 29.000 322.000 34.600 ;
        RECT 324.400 32.000 325.200 39.800 ;
        RECT 327.600 35.200 328.400 39.800 ;
        RECT 303.200 27.800 304.000 28.000 ;
        RECT 303.200 27.200 307.600 27.800 ;
        RECT 306.800 27.000 307.600 27.200 ;
        RECT 308.400 26.800 309.200 28.400 ;
        RECT 295.600 25.400 298.000 26.200 ;
        RECT 300.400 25.600 301.400 26.400 ;
        RECT 304.400 25.600 306.000 26.400 ;
        RECT 306.800 26.200 307.600 26.400 ;
        RECT 310.600 26.200 311.400 28.600 ;
        RECT 313.200 28.200 322.000 29.000 ;
        RECT 316.600 26.800 319.600 27.600 ;
        RECT 316.600 26.200 317.400 26.800 ;
        RECT 306.800 25.600 311.400 26.200 ;
        RECT 297.200 22.200 298.000 25.400 ;
        RECT 314.800 25.400 317.400 26.200 ;
        RECT 298.800 22.200 299.600 25.000 ;
        RECT 300.400 22.200 301.200 25.000 ;
        RECT 302.000 22.200 302.800 25.000 ;
        RECT 303.600 22.200 304.400 25.000 ;
        RECT 306.800 22.200 307.600 25.000 ;
        RECT 310.000 22.200 310.800 25.000 ;
        RECT 311.600 22.200 312.400 25.000 ;
        RECT 313.200 22.200 314.000 25.000 ;
        RECT 314.800 22.200 315.600 25.400 ;
        RECT 321.200 22.200 322.000 28.200 ;
        RECT 324.200 31.200 325.200 32.000 ;
        RECT 325.800 34.600 328.400 35.200 ;
        RECT 325.800 33.000 326.400 34.600 ;
        RECT 330.800 34.400 331.600 39.800 ;
        RECT 334.000 37.000 334.800 39.800 ;
        RECT 335.600 37.000 336.400 39.800 ;
        RECT 337.200 37.000 338.000 39.800 ;
        RECT 332.200 34.400 336.400 35.200 ;
        RECT 329.000 33.600 331.600 34.400 ;
        RECT 338.800 33.600 339.600 39.800 ;
        RECT 342.000 35.000 342.800 39.800 ;
        RECT 345.200 35.000 346.000 39.800 ;
        RECT 346.800 37.000 347.600 39.800 ;
        RECT 348.400 37.000 349.200 39.800 ;
        RECT 351.600 35.200 352.400 39.800 ;
        RECT 354.800 36.400 355.600 39.800 ;
        RECT 354.800 35.800 355.800 36.400 ;
        RECT 355.200 35.200 355.800 35.800 ;
        RECT 350.400 34.400 354.600 35.200 ;
        RECT 355.200 34.600 357.200 35.200 ;
        RECT 342.000 33.600 344.600 34.400 ;
        RECT 345.200 33.800 351.000 34.400 ;
        RECT 354.000 34.000 354.600 34.400 ;
        RECT 334.000 33.000 334.800 33.200 ;
        RECT 325.800 32.400 334.800 33.000 ;
        RECT 337.200 33.000 338.000 33.200 ;
        RECT 345.200 33.000 345.800 33.800 ;
        RECT 351.600 33.200 353.000 33.800 ;
        RECT 354.000 33.200 355.600 34.000 ;
        RECT 337.200 32.400 345.800 33.000 ;
        RECT 346.800 33.000 353.000 33.200 ;
        RECT 346.800 32.600 352.200 33.000 ;
        RECT 346.800 32.400 347.600 32.600 ;
        RECT 324.200 26.800 325.000 31.200 ;
        RECT 325.800 30.600 326.400 32.400 ;
        RECT 325.600 30.000 326.400 30.600 ;
        RECT 332.400 30.000 355.800 30.600 ;
        RECT 325.600 28.000 326.200 30.000 ;
        RECT 332.400 29.400 333.200 30.000 ;
        RECT 343.600 29.600 344.400 30.000 ;
        RECT 350.000 29.600 350.800 30.000 ;
        RECT 355.000 29.800 355.800 30.000 ;
        RECT 326.800 28.600 330.600 29.400 ;
        RECT 325.600 27.400 326.800 28.000 ;
        RECT 324.200 26.000 325.200 26.800 ;
        RECT 324.400 22.200 325.200 26.000 ;
        RECT 326.000 22.200 326.800 27.400 ;
        RECT 329.800 27.400 330.600 28.600 ;
        RECT 329.800 26.800 331.600 27.400 ;
        RECT 330.800 26.200 331.600 26.800 ;
        RECT 335.600 26.400 336.400 29.200 ;
        RECT 338.800 28.600 342.000 29.400 ;
        RECT 345.800 28.600 347.800 29.400 ;
        RECT 356.400 29.000 357.200 34.600 ;
        RECT 359.600 31.200 360.400 39.800 ;
        RECT 362.800 31.200 363.600 39.800 ;
        RECT 366.000 31.200 366.800 39.800 ;
        RECT 369.200 31.200 370.000 39.800 ;
        RECT 374.000 36.400 374.800 39.800 ;
        RECT 373.800 35.800 374.800 36.400 ;
        RECT 373.800 35.200 374.400 35.800 ;
        RECT 377.200 35.200 378.000 39.800 ;
        RECT 380.400 37.000 381.200 39.800 ;
        RECT 382.000 37.000 382.800 39.800 ;
        RECT 338.400 27.800 339.200 28.000 ;
        RECT 338.400 27.200 342.800 27.800 ;
        RECT 342.000 27.000 342.800 27.200 ;
        RECT 343.600 26.800 344.400 28.400 ;
        RECT 330.800 25.400 333.200 26.200 ;
        RECT 335.600 25.600 336.600 26.400 ;
        RECT 339.600 25.600 341.200 26.400 ;
        RECT 342.000 26.200 342.800 26.400 ;
        RECT 345.800 26.200 346.600 28.600 ;
        RECT 348.400 28.200 357.200 29.000 ;
        RECT 351.800 26.800 354.800 27.600 ;
        RECT 351.800 26.200 352.600 26.800 ;
        RECT 342.000 25.600 346.600 26.200 ;
        RECT 332.400 22.200 333.200 25.400 ;
        RECT 350.000 25.400 352.600 26.200 ;
        RECT 334.000 22.200 334.800 25.000 ;
        RECT 335.600 22.200 336.400 25.000 ;
        RECT 337.200 22.200 338.000 25.000 ;
        RECT 338.800 22.200 339.600 25.000 ;
        RECT 342.000 22.200 342.800 25.000 ;
        RECT 345.200 22.200 346.000 25.000 ;
        RECT 346.800 22.200 347.600 25.000 ;
        RECT 348.400 22.200 349.200 25.000 ;
        RECT 350.000 22.200 350.800 25.400 ;
        RECT 356.400 22.200 357.200 28.200 ;
        RECT 358.000 30.400 360.400 31.200 ;
        RECT 361.400 30.400 363.600 31.200 ;
        RECT 364.600 30.400 366.800 31.200 ;
        RECT 368.200 30.400 370.000 31.200 ;
        RECT 372.400 34.600 374.400 35.200 ;
        RECT 358.000 27.600 358.800 30.400 ;
        RECT 361.400 29.000 362.200 30.400 ;
        RECT 364.600 29.000 365.400 30.400 ;
        RECT 368.200 29.000 369.000 30.400 ;
        RECT 359.600 28.200 362.200 29.000 ;
        RECT 363.000 28.200 365.400 29.000 ;
        RECT 366.400 28.200 369.000 29.000 ;
        RECT 361.400 27.600 362.200 28.200 ;
        RECT 364.600 27.600 365.400 28.200 ;
        RECT 368.200 27.600 369.000 28.200 ;
        RECT 372.400 29.000 373.200 34.600 ;
        RECT 375.000 34.400 379.200 35.200 ;
        RECT 383.600 35.000 384.400 39.800 ;
        RECT 386.800 35.000 387.600 39.800 ;
        RECT 375.000 34.000 375.600 34.400 ;
        RECT 374.000 33.200 375.600 34.000 ;
        RECT 378.600 33.800 384.400 34.400 ;
        RECT 376.600 33.200 378.000 33.800 ;
        RECT 376.600 33.000 382.800 33.200 ;
        RECT 377.400 32.600 382.800 33.000 ;
        RECT 382.000 32.400 382.800 32.600 ;
        RECT 383.800 33.000 384.400 33.800 ;
        RECT 385.000 33.600 387.600 34.400 ;
        RECT 390.000 33.600 390.800 39.800 ;
        RECT 391.600 37.000 392.400 39.800 ;
        RECT 393.200 37.000 394.000 39.800 ;
        RECT 394.800 37.000 395.600 39.800 ;
        RECT 393.200 34.400 397.400 35.200 ;
        RECT 398.000 34.400 398.800 39.800 ;
        RECT 401.200 35.200 402.000 39.800 ;
        RECT 401.200 34.600 403.800 35.200 ;
        RECT 398.000 33.600 400.600 34.400 ;
        RECT 391.600 33.000 392.400 33.200 ;
        RECT 383.800 32.400 392.400 33.000 ;
        RECT 394.800 33.000 395.600 33.200 ;
        RECT 403.200 33.000 403.800 34.600 ;
        RECT 394.800 32.400 403.800 33.000 ;
        RECT 403.200 30.600 403.800 32.400 ;
        RECT 404.400 32.000 405.200 39.800 ;
        RECT 409.200 38.300 410.000 39.800 ;
        RECT 414.000 38.300 414.800 38.400 ;
        RECT 409.200 37.700 414.800 38.300 ;
        RECT 404.400 31.200 405.400 32.000 ;
        RECT 373.800 30.000 397.200 30.600 ;
        RECT 403.200 30.000 404.000 30.600 ;
        RECT 373.800 29.800 374.600 30.000 ;
        RECT 377.200 29.600 378.000 30.000 ;
        RECT 378.800 29.600 379.600 30.000 ;
        RECT 396.400 29.400 397.200 30.000 ;
        RECT 372.400 28.200 381.200 29.000 ;
        RECT 381.800 28.600 383.800 29.400 ;
        RECT 387.600 28.600 390.800 29.400 ;
        RECT 358.000 26.800 360.400 27.600 ;
        RECT 361.400 26.800 363.600 27.600 ;
        RECT 364.600 26.800 366.800 27.600 ;
        RECT 368.200 26.800 370.000 27.600 ;
        RECT 359.600 22.200 360.400 26.800 ;
        RECT 362.800 22.200 363.600 26.800 ;
        RECT 366.000 22.200 366.800 26.800 ;
        RECT 369.200 22.200 370.000 26.800 ;
        RECT 372.400 22.200 373.200 28.200 ;
        RECT 374.800 26.800 377.800 27.600 ;
        RECT 377.000 26.200 377.800 26.800 ;
        RECT 383.000 26.200 383.800 28.600 ;
        RECT 385.200 26.800 386.000 28.400 ;
        RECT 390.400 27.800 391.200 28.000 ;
        RECT 386.800 27.200 391.200 27.800 ;
        RECT 386.800 27.000 387.600 27.200 ;
        RECT 393.200 26.400 394.000 29.200 ;
        RECT 399.000 28.600 402.800 29.400 ;
        RECT 399.000 27.400 399.800 28.600 ;
        RECT 403.400 28.000 404.000 30.000 ;
        RECT 386.800 26.200 387.600 26.400 ;
        RECT 377.000 25.400 379.600 26.200 ;
        RECT 383.000 25.600 387.600 26.200 ;
        RECT 388.400 25.600 390.000 26.400 ;
        RECT 393.000 25.600 394.000 26.400 ;
        RECT 398.000 26.800 399.800 27.400 ;
        RECT 402.800 27.400 404.000 28.000 ;
        RECT 398.000 26.200 398.800 26.800 ;
        RECT 378.800 22.200 379.600 25.400 ;
        RECT 396.400 25.400 398.800 26.200 ;
        RECT 380.400 22.200 381.200 25.000 ;
        RECT 382.000 22.200 382.800 25.000 ;
        RECT 383.600 22.200 384.400 25.000 ;
        RECT 386.800 22.200 387.600 25.000 ;
        RECT 390.000 22.200 390.800 25.000 ;
        RECT 391.600 22.200 392.400 25.000 ;
        RECT 393.200 22.200 394.000 25.000 ;
        RECT 394.800 22.200 395.600 25.000 ;
        RECT 396.400 22.200 397.200 25.400 ;
        RECT 402.800 22.200 403.600 27.400 ;
        RECT 404.600 26.800 405.400 31.200 ;
        RECT 404.400 26.000 405.400 26.800 ;
        RECT 404.400 22.200 405.200 26.000 ;
        RECT 407.600 24.800 408.400 26.400 ;
        RECT 409.200 22.200 410.000 37.700 ;
        RECT 414.000 37.600 414.800 37.700 ;
        RECT 418.800 36.400 419.600 39.800 ;
        RECT 418.600 35.800 419.600 36.400 ;
        RECT 418.600 35.200 419.200 35.800 ;
        RECT 422.000 35.200 422.800 39.800 ;
        RECT 425.200 37.000 426.000 39.800 ;
        RECT 426.800 37.000 427.600 39.800 ;
        RECT 417.200 34.600 419.200 35.200 ;
        RECT 417.200 29.000 418.000 34.600 ;
        RECT 419.800 34.400 424.000 35.200 ;
        RECT 428.400 35.000 429.200 39.800 ;
        RECT 431.600 35.000 432.400 39.800 ;
        RECT 419.800 34.000 420.400 34.400 ;
        RECT 418.800 33.200 420.400 34.000 ;
        RECT 423.400 33.800 429.200 34.400 ;
        RECT 421.400 33.200 422.800 33.800 ;
        RECT 421.400 33.000 427.600 33.200 ;
        RECT 422.200 32.600 427.600 33.000 ;
        RECT 426.800 32.400 427.600 32.600 ;
        RECT 428.600 33.000 429.200 33.800 ;
        RECT 429.800 33.600 432.400 34.400 ;
        RECT 434.800 33.600 435.600 39.800 ;
        RECT 436.400 37.000 437.200 39.800 ;
        RECT 438.000 37.000 438.800 39.800 ;
        RECT 439.600 37.000 440.400 39.800 ;
        RECT 438.000 34.400 442.200 35.200 ;
        RECT 442.800 34.400 443.600 39.800 ;
        RECT 446.000 35.200 446.800 39.800 ;
        RECT 446.000 34.600 448.600 35.200 ;
        RECT 442.800 33.600 445.400 34.400 ;
        RECT 436.400 33.000 437.200 33.200 ;
        RECT 428.600 32.400 437.200 33.000 ;
        RECT 439.600 33.000 440.400 33.200 ;
        RECT 448.000 33.000 448.600 34.600 ;
        RECT 439.600 32.400 448.600 33.000 ;
        RECT 448.000 30.600 448.600 32.400 ;
        RECT 449.200 32.000 450.000 39.800 ;
        RECT 449.200 31.200 450.200 32.000 ;
        RECT 418.600 30.000 442.000 30.600 ;
        RECT 448.000 30.000 448.800 30.600 ;
        RECT 418.600 29.800 419.400 30.000 ;
        RECT 420.400 29.600 421.200 30.000 ;
        RECT 423.600 29.600 424.400 30.000 ;
        RECT 441.200 29.400 442.000 30.000 ;
        RECT 417.200 28.200 426.000 29.000 ;
        RECT 426.600 28.600 428.600 29.400 ;
        RECT 432.400 28.600 435.600 29.400 ;
        RECT 417.200 22.200 418.000 28.200 ;
        RECT 419.600 26.800 422.600 27.600 ;
        RECT 421.800 26.200 422.600 26.800 ;
        RECT 427.800 26.200 428.600 28.600 ;
        RECT 430.000 26.800 430.800 28.400 ;
        RECT 435.200 27.800 436.000 28.000 ;
        RECT 431.600 27.200 436.000 27.800 ;
        RECT 431.600 27.000 432.400 27.200 ;
        RECT 438.000 26.400 438.800 29.200 ;
        RECT 443.800 28.600 447.600 29.400 ;
        RECT 443.800 27.400 444.600 28.600 ;
        RECT 448.200 28.000 448.800 30.000 ;
        RECT 431.600 26.200 432.400 26.400 ;
        RECT 421.800 25.400 424.400 26.200 ;
        RECT 427.800 25.600 432.400 26.200 ;
        RECT 433.200 25.600 434.800 26.400 ;
        RECT 437.800 25.600 438.800 26.400 ;
        RECT 442.800 26.800 444.600 27.400 ;
        RECT 447.600 27.400 448.800 28.000 ;
        RECT 442.800 26.200 443.600 26.800 ;
        RECT 423.600 22.200 424.400 25.400 ;
        RECT 441.200 25.400 443.600 26.200 ;
        RECT 425.200 22.200 426.000 25.000 ;
        RECT 426.800 22.200 427.600 25.000 ;
        RECT 428.400 22.200 429.200 25.000 ;
        RECT 431.600 22.200 432.400 25.000 ;
        RECT 434.800 22.200 435.600 25.000 ;
        RECT 436.400 22.200 437.200 25.000 ;
        RECT 438.000 22.200 438.800 25.000 ;
        RECT 439.600 22.200 440.400 25.000 ;
        RECT 441.200 22.200 442.000 25.400 ;
        RECT 447.600 22.200 448.400 27.400 ;
        RECT 449.400 26.800 450.200 31.200 ;
        RECT 449.200 26.000 450.200 26.800 ;
        RECT 452.400 31.200 453.200 39.800 ;
        RECT 456.600 35.800 457.800 39.800 ;
        RECT 461.200 35.800 462.000 39.800 ;
        RECT 465.600 36.400 466.400 39.800 ;
        RECT 465.600 35.800 467.600 36.400 ;
        RECT 457.200 35.000 458.000 35.800 ;
        RECT 461.400 35.200 462.000 35.800 ;
        RECT 460.600 34.600 464.200 35.200 ;
        RECT 466.800 35.000 467.600 35.800 ;
        RECT 460.600 34.400 461.400 34.600 ;
        RECT 463.400 34.400 464.200 34.600 ;
        RECT 456.400 33.200 457.800 34.000 ;
        RECT 457.200 32.200 457.800 33.200 ;
        RECT 459.400 33.000 461.600 33.600 ;
        RECT 459.400 32.800 460.200 33.000 ;
        RECT 457.200 31.600 459.600 32.200 ;
        RECT 452.400 30.600 456.600 31.200 ;
        RECT 452.400 27.200 453.200 30.600 ;
        RECT 455.800 30.400 456.600 30.600 ;
        RECT 459.000 30.400 459.600 31.600 ;
        RECT 461.000 31.800 461.600 33.000 ;
        RECT 462.200 33.000 463.000 33.200 ;
        RECT 466.800 33.000 467.600 33.200 ;
        RECT 462.200 32.400 467.600 33.000 ;
        RECT 461.000 31.400 465.800 31.800 ;
        RECT 470.000 31.400 470.800 39.800 ;
        RECT 461.000 31.200 470.800 31.400 ;
        RECT 465.000 31.000 470.800 31.200 ;
        RECT 465.200 30.800 470.800 31.000 ;
        RECT 454.200 29.800 455.000 30.000 ;
        RECT 454.200 29.200 458.000 29.800 ;
        RECT 458.800 29.600 459.600 30.400 ;
        RECT 463.600 30.200 464.400 30.400 ;
        RECT 463.600 29.600 468.600 30.200 ;
        RECT 457.200 29.000 458.000 29.200 ;
        RECT 459.000 28.400 459.600 29.600 ;
        RECT 465.200 29.400 466.000 29.600 ;
        RECT 467.800 29.400 468.600 29.600 ;
        RECT 466.200 28.400 467.000 28.600 ;
        RECT 459.000 27.800 470.000 28.400 ;
        RECT 459.400 27.600 460.200 27.800 ;
        RECT 452.400 26.600 456.400 27.200 ;
        RECT 449.200 22.200 450.000 26.000 ;
        RECT 452.400 22.200 453.200 26.600 ;
        RECT 455.400 26.400 456.400 26.600 ;
        RECT 455.600 26.300 456.400 26.400 ;
        RECT 458.800 26.300 459.600 26.400 ;
        RECT 455.600 25.700 459.600 26.300 ;
        RECT 458.800 25.600 459.600 25.700 ;
        RECT 465.200 25.600 465.800 27.800 ;
        RECT 468.400 27.600 470.000 27.800 ;
        RECT 473.200 28.300 474.000 39.800 ;
        RECT 477.400 32.400 478.200 39.800 ;
        RECT 478.800 33.600 479.600 34.400 ;
        RECT 479.000 32.400 479.600 33.600 ;
        RECT 477.400 31.800 478.400 32.400 ;
        RECT 479.000 31.800 480.400 32.400 ;
        RECT 482.800 32.000 483.600 39.800 ;
        RECT 486.000 35.200 486.800 39.800 ;
        RECT 476.400 28.800 477.200 30.400 ;
        RECT 477.800 28.400 478.400 31.800 ;
        RECT 479.600 31.600 480.400 31.800 ;
        RECT 482.600 31.200 483.600 32.000 ;
        RECT 484.200 34.600 486.800 35.200 ;
        RECT 484.200 33.000 484.800 34.600 ;
        RECT 489.200 34.400 490.000 39.800 ;
        RECT 492.400 37.000 493.200 39.800 ;
        RECT 494.000 37.000 494.800 39.800 ;
        RECT 495.600 37.000 496.400 39.800 ;
        RECT 490.600 34.400 494.800 35.200 ;
        RECT 487.400 33.600 490.000 34.400 ;
        RECT 497.200 33.600 498.000 39.800 ;
        RECT 500.400 35.000 501.200 39.800 ;
        RECT 503.600 35.000 504.400 39.800 ;
        RECT 505.200 37.000 506.000 39.800 ;
        RECT 506.800 37.000 507.600 39.800 ;
        RECT 510.000 35.200 510.800 39.800 ;
        RECT 513.200 36.400 514.000 39.800 ;
        RECT 520.200 38.400 521.000 39.800 ;
        RECT 519.600 37.600 521.000 38.400 ;
        RECT 513.200 35.800 514.200 36.400 ;
        RECT 513.600 35.200 514.200 35.800 ;
        RECT 508.800 34.400 513.000 35.200 ;
        RECT 513.600 34.600 515.600 35.200 ;
        RECT 500.400 33.600 503.000 34.400 ;
        RECT 503.600 33.800 509.400 34.400 ;
        RECT 512.400 34.000 513.000 34.400 ;
        RECT 492.400 33.000 493.200 33.200 ;
        RECT 484.200 32.400 493.200 33.000 ;
        RECT 495.600 33.000 496.400 33.200 ;
        RECT 503.600 33.000 504.200 33.800 ;
        RECT 510.000 33.200 511.400 33.800 ;
        RECT 512.400 33.200 514.000 34.000 ;
        RECT 495.600 32.400 504.200 33.000 ;
        RECT 505.200 33.000 511.400 33.200 ;
        RECT 505.200 32.600 510.600 33.000 ;
        RECT 505.200 32.400 506.000 32.600 ;
        RECT 474.800 28.300 475.600 28.400 ;
        RECT 473.200 28.200 475.600 28.300 ;
        RECT 473.200 27.700 476.400 28.200 ;
        RECT 463.400 25.400 464.200 25.600 ;
        RECT 457.200 24.200 458.000 25.000 ;
        RECT 461.400 24.800 464.200 25.400 ;
        RECT 465.200 24.800 466.000 25.600 ;
        RECT 461.400 24.200 462.000 24.800 ;
        RECT 466.800 24.200 467.600 25.000 ;
        RECT 456.600 23.600 458.000 24.200 ;
        RECT 456.600 22.200 457.800 23.600 ;
        RECT 461.200 22.200 462.000 24.200 ;
        RECT 465.600 23.600 467.600 24.200 ;
        RECT 465.600 22.200 466.400 23.600 ;
        RECT 470.000 22.200 470.800 27.000 ;
        RECT 471.600 24.800 472.400 26.400 ;
        RECT 473.200 22.200 474.000 27.700 ;
        RECT 474.800 27.600 476.400 27.700 ;
        RECT 477.800 27.600 480.400 28.400 ;
        RECT 475.600 27.200 476.400 27.600 ;
        RECT 475.000 26.200 478.600 26.600 ;
        RECT 479.600 26.200 480.200 27.600 ;
        RECT 482.600 26.800 483.400 31.200 ;
        RECT 484.200 30.600 484.800 32.400 ;
        RECT 484.000 30.000 484.800 30.600 ;
        RECT 490.800 30.000 514.200 30.600 ;
        RECT 484.000 28.000 484.600 30.000 ;
        RECT 490.800 29.400 491.600 30.000 ;
        RECT 508.400 29.600 509.200 30.000 ;
        RECT 510.000 29.600 510.800 30.000 ;
        RECT 513.400 29.800 514.200 30.000 ;
        RECT 485.200 28.600 489.000 29.400 ;
        RECT 484.000 27.400 485.200 28.000 ;
        RECT 474.800 26.000 478.800 26.200 ;
        RECT 474.800 22.200 475.600 26.000 ;
        RECT 478.000 22.200 478.800 26.000 ;
        RECT 479.600 22.200 480.400 26.200 ;
        RECT 482.600 26.000 483.600 26.800 ;
        RECT 482.800 22.200 483.600 26.000 ;
        RECT 484.400 22.200 485.200 27.400 ;
        RECT 488.200 27.400 489.000 28.600 ;
        RECT 488.200 26.800 490.000 27.400 ;
        RECT 489.200 26.200 490.000 26.800 ;
        RECT 494.000 26.400 494.800 29.200 ;
        RECT 497.200 28.600 500.400 29.400 ;
        RECT 504.200 28.600 506.200 29.400 ;
        RECT 514.800 29.000 515.600 34.600 ;
        RECT 520.200 32.800 521.000 37.600 ;
        RECT 524.400 35.000 525.200 39.000 ;
        RECT 519.400 32.200 521.000 32.800 ;
        RECT 518.000 29.600 518.800 31.200 ;
        RECT 496.800 27.800 497.600 28.000 ;
        RECT 496.800 27.200 501.200 27.800 ;
        RECT 500.400 27.000 501.200 27.200 ;
        RECT 502.000 26.800 502.800 28.400 ;
        RECT 489.200 25.400 491.600 26.200 ;
        RECT 494.000 25.600 495.000 26.400 ;
        RECT 498.000 25.600 499.600 26.400 ;
        RECT 500.400 26.200 501.200 26.400 ;
        RECT 504.200 26.200 505.000 28.600 ;
        RECT 506.800 28.200 515.600 29.000 ;
        RECT 519.400 28.400 520.000 32.200 ;
        RECT 524.600 31.600 525.200 35.000 ;
        RECT 521.400 31.000 525.200 31.600 ;
        RECT 526.000 35.000 526.800 39.000 ;
        RECT 530.200 38.400 531.000 39.800 ;
        RECT 530.200 37.600 531.600 38.400 ;
        RECT 526.000 31.600 526.600 35.000 ;
        RECT 530.200 32.800 531.000 37.600 ;
        RECT 530.200 32.200 531.800 32.800 ;
        RECT 526.000 31.000 529.800 31.600 ;
        RECT 521.400 29.000 522.000 31.000 ;
        RECT 510.200 26.800 513.200 27.600 ;
        RECT 510.200 26.200 511.000 26.800 ;
        RECT 500.400 25.600 505.000 26.200 ;
        RECT 490.800 22.200 491.600 25.400 ;
        RECT 508.400 25.400 511.000 26.200 ;
        RECT 492.400 22.200 493.200 25.000 ;
        RECT 494.000 22.200 494.800 25.000 ;
        RECT 495.600 22.200 496.400 25.000 ;
        RECT 497.200 22.200 498.000 25.000 ;
        RECT 500.400 22.200 501.200 25.000 ;
        RECT 503.600 22.200 504.400 25.000 ;
        RECT 505.200 22.200 506.000 25.000 ;
        RECT 506.800 22.200 507.600 25.000 ;
        RECT 508.400 22.200 509.200 25.400 ;
        RECT 514.800 22.200 515.600 28.200 ;
        RECT 518.000 27.600 520.000 28.400 ;
        RECT 520.600 28.200 522.000 29.000 ;
        RECT 522.800 28.800 523.600 30.400 ;
        RECT 524.400 30.300 525.200 30.400 ;
        RECT 526.000 30.300 526.800 30.400 ;
        RECT 524.400 29.700 526.800 30.300 ;
        RECT 524.400 28.800 525.200 29.700 ;
        RECT 526.000 28.800 526.800 29.700 ;
        RECT 527.600 28.800 528.400 30.400 ;
        RECT 529.200 29.000 529.800 31.000 ;
        RECT 519.400 27.000 520.000 27.600 ;
        RECT 521.000 27.800 522.000 28.200 ;
        RECT 529.200 28.200 530.600 29.000 ;
        RECT 531.200 28.400 531.800 32.200 ;
        RECT 537.200 31.200 538.000 39.800 ;
        RECT 540.400 31.200 541.200 39.800 ;
        RECT 543.600 31.200 544.400 39.800 ;
        RECT 546.800 31.200 547.600 39.800 ;
        RECT 532.400 29.600 533.200 31.200 ;
        RECT 537.200 30.400 539.000 31.200 ;
        RECT 540.400 30.400 542.600 31.200 ;
        RECT 543.600 30.400 545.800 31.200 ;
        RECT 546.800 30.400 549.200 31.200 ;
        RECT 538.200 29.000 539.000 30.400 ;
        RECT 541.800 29.000 542.600 30.400 ;
        RECT 545.000 29.000 545.800 30.400 ;
        RECT 529.200 27.800 530.200 28.200 ;
        RECT 521.000 27.200 525.200 27.800 ;
        RECT 519.400 26.600 520.200 27.000 ;
        RECT 519.400 26.000 521.000 26.600 ;
        RECT 520.200 23.000 521.000 26.000 ;
        RECT 524.600 25.000 525.200 27.200 ;
        RECT 524.400 23.000 525.200 25.000 ;
        RECT 526.000 27.200 530.200 27.800 ;
        RECT 531.200 27.600 533.200 28.400 ;
        RECT 538.200 28.200 540.800 29.000 ;
        RECT 541.800 28.200 544.200 29.000 ;
        RECT 545.000 28.200 547.600 29.000 ;
        RECT 538.200 27.600 539.000 28.200 ;
        RECT 541.800 27.600 542.600 28.200 ;
        RECT 545.000 27.600 545.800 28.200 ;
        RECT 548.400 27.600 549.200 30.400 ;
        RECT 526.000 25.000 526.600 27.200 ;
        RECT 531.200 27.000 531.800 27.600 ;
        RECT 531.000 26.600 531.800 27.000 ;
        RECT 530.200 26.000 531.800 26.600 ;
        RECT 537.200 26.800 539.000 27.600 ;
        RECT 540.400 26.800 542.600 27.600 ;
        RECT 543.600 26.800 545.800 27.600 ;
        RECT 546.800 26.800 549.200 27.600 ;
        RECT 526.000 23.000 526.800 25.000 ;
        RECT 530.200 23.000 531.000 26.000 ;
        RECT 537.200 22.200 538.000 26.800 ;
        RECT 540.400 22.200 541.200 26.800 ;
        RECT 543.600 22.200 544.400 26.800 ;
        RECT 546.800 22.200 547.600 26.800 ;
        RECT 2.800 16.000 3.600 19.800 ;
        RECT 2.600 15.200 3.600 16.000 ;
        RECT 2.600 10.800 3.400 15.200 ;
        RECT 4.400 14.600 5.200 19.800 ;
        RECT 10.800 16.600 11.600 19.800 ;
        RECT 12.400 17.000 13.200 19.800 ;
        RECT 14.000 17.000 14.800 19.800 ;
        RECT 15.600 17.000 16.400 19.800 ;
        RECT 17.200 17.000 18.000 19.800 ;
        RECT 20.400 17.000 21.200 19.800 ;
        RECT 23.600 17.000 24.400 19.800 ;
        RECT 25.200 17.000 26.000 19.800 ;
        RECT 26.800 17.000 27.600 19.800 ;
        RECT 9.200 15.800 11.600 16.600 ;
        RECT 28.400 16.600 29.200 19.800 ;
        RECT 9.200 15.200 10.000 15.800 ;
        RECT 4.000 14.000 5.200 14.600 ;
        RECT 8.200 14.600 10.000 15.200 ;
        RECT 14.000 15.600 15.000 16.400 ;
        RECT 18.000 15.600 19.600 16.400 ;
        RECT 20.400 15.800 25.000 16.400 ;
        RECT 28.400 15.800 31.000 16.600 ;
        RECT 20.400 15.600 21.200 15.800 ;
        RECT 4.000 12.000 4.600 14.000 ;
        RECT 8.200 13.400 9.000 14.600 ;
        RECT 5.200 12.600 9.000 13.400 ;
        RECT 14.000 12.800 14.800 15.600 ;
        RECT 20.400 14.800 21.200 15.000 ;
        RECT 16.800 14.200 21.200 14.800 ;
        RECT 16.800 14.000 17.600 14.200 ;
        RECT 22.000 13.600 22.800 15.200 ;
        RECT 24.200 13.400 25.000 15.800 ;
        RECT 30.200 15.200 31.000 15.800 ;
        RECT 30.200 14.400 33.200 15.200 ;
        RECT 34.800 13.800 35.600 19.800 ;
        RECT 17.200 12.600 20.400 13.400 ;
        RECT 24.200 12.600 26.200 13.400 ;
        RECT 26.800 13.000 35.600 13.800 ;
        RECT 10.800 12.000 11.600 12.600 ;
        RECT 28.400 12.000 29.200 12.400 ;
        RECT 31.600 12.000 32.400 12.400 ;
        RECT 33.400 12.000 34.200 12.200 ;
        RECT 4.000 11.400 4.800 12.000 ;
        RECT 10.800 11.400 34.200 12.000 ;
        RECT 2.600 10.000 3.600 10.800 ;
        RECT 2.800 2.200 3.600 10.000 ;
        RECT 4.200 9.600 4.800 11.400 ;
        RECT 4.200 9.000 13.200 9.600 ;
        RECT 4.200 7.400 4.800 9.000 ;
        RECT 12.400 8.800 13.200 9.000 ;
        RECT 15.600 9.000 24.200 9.600 ;
        RECT 15.600 8.800 16.400 9.000 ;
        RECT 7.400 7.600 10.000 8.400 ;
        RECT 4.200 6.800 6.800 7.400 ;
        RECT 6.000 2.200 6.800 6.800 ;
        RECT 9.200 2.200 10.000 7.600 ;
        RECT 10.600 6.800 14.800 7.600 ;
        RECT 12.400 2.200 13.200 5.000 ;
        RECT 14.000 2.200 14.800 5.000 ;
        RECT 15.600 2.200 16.400 5.000 ;
        RECT 17.200 2.200 18.000 8.400 ;
        RECT 20.400 7.600 23.000 8.400 ;
        RECT 23.600 8.200 24.200 9.000 ;
        RECT 25.200 9.400 26.000 9.600 ;
        RECT 25.200 9.000 30.600 9.400 ;
        RECT 25.200 8.800 31.400 9.000 ;
        RECT 30.000 8.200 31.400 8.800 ;
        RECT 23.600 7.600 29.400 8.200 ;
        RECT 32.400 8.000 34.000 8.800 ;
        RECT 32.400 7.600 33.000 8.000 ;
        RECT 20.400 2.200 21.200 7.000 ;
        RECT 23.600 2.200 24.400 7.000 ;
        RECT 28.800 6.800 33.000 7.600 ;
        RECT 34.800 7.400 35.600 13.000 ;
        RECT 33.600 6.800 35.600 7.400 ;
        RECT 36.400 13.800 37.200 19.800 ;
        RECT 42.800 16.600 43.600 19.800 ;
        RECT 44.400 17.000 45.200 19.800 ;
        RECT 46.000 17.000 46.800 19.800 ;
        RECT 47.600 17.000 48.400 19.800 ;
        RECT 50.800 17.000 51.600 19.800 ;
        RECT 54.000 17.000 54.800 19.800 ;
        RECT 55.600 17.000 56.400 19.800 ;
        RECT 57.200 17.000 58.000 19.800 ;
        RECT 58.800 17.000 59.600 19.800 ;
        RECT 41.000 15.800 43.600 16.600 ;
        RECT 60.400 16.600 61.200 19.800 ;
        RECT 47.000 15.800 51.600 16.400 ;
        RECT 41.000 15.200 41.800 15.800 ;
        RECT 38.800 14.400 41.800 15.200 ;
        RECT 36.400 13.000 45.200 13.800 ;
        RECT 47.000 13.400 47.800 15.800 ;
        RECT 50.800 15.600 51.600 15.800 ;
        RECT 52.400 15.600 54.000 16.400 ;
        RECT 57.000 15.600 58.000 16.400 ;
        RECT 60.400 15.800 62.800 16.600 ;
        RECT 49.200 13.600 50.000 15.200 ;
        RECT 50.800 14.800 51.600 15.000 ;
        RECT 50.800 14.200 55.200 14.800 ;
        RECT 54.400 14.000 55.200 14.200 ;
        RECT 36.400 7.400 37.200 13.000 ;
        RECT 45.800 12.600 47.800 13.400 ;
        RECT 51.600 12.600 54.800 13.400 ;
        RECT 57.200 12.800 58.000 15.600 ;
        RECT 62.000 15.200 62.800 15.800 ;
        RECT 62.000 14.600 63.800 15.200 ;
        RECT 63.000 13.400 63.800 14.600 ;
        RECT 66.800 14.600 67.600 19.800 ;
        RECT 68.400 16.000 69.200 19.800 ;
        RECT 72.200 16.800 73.000 19.800 ;
        RECT 68.400 15.200 69.400 16.000 ;
        RECT 66.800 14.000 68.000 14.600 ;
        RECT 63.000 12.600 66.800 13.400 ;
        RECT 37.800 12.000 38.600 12.200 ;
        RECT 42.800 12.000 43.600 12.400 ;
        RECT 60.400 12.000 61.200 12.600 ;
        RECT 67.400 12.000 68.000 14.000 ;
        RECT 37.800 11.400 61.200 12.000 ;
        RECT 67.200 11.400 68.000 12.000 ;
        RECT 67.200 9.600 67.800 11.400 ;
        RECT 68.600 10.800 69.400 15.200 ;
        RECT 71.600 15.800 73.000 16.800 ;
        RECT 76.400 15.800 77.200 19.800 ;
        RECT 78.000 15.800 78.800 19.800 ;
        RECT 82.200 16.800 83.000 19.800 ;
        RECT 82.200 15.800 83.600 16.800 ;
        RECT 71.600 12.400 72.200 15.800 ;
        RECT 76.400 15.600 77.000 15.800 ;
        RECT 75.200 15.200 77.000 15.600 ;
        RECT 72.800 15.000 77.000 15.200 ;
        RECT 78.200 15.600 78.800 15.800 ;
        RECT 78.200 15.200 80.000 15.600 ;
        RECT 78.200 15.000 82.400 15.200 ;
        RECT 72.800 14.600 75.800 15.000 ;
        RECT 79.400 14.600 82.400 15.000 ;
        RECT 72.800 14.400 73.600 14.600 ;
        RECT 81.600 14.400 82.400 14.600 ;
        RECT 70.000 12.300 70.800 12.400 ;
        RECT 71.600 12.300 72.400 12.400 ;
        RECT 70.000 11.700 72.400 12.300 ;
        RECT 70.000 11.600 70.800 11.700 ;
        RECT 71.600 11.600 72.400 11.700 ;
        RECT 46.000 9.400 46.800 9.600 ;
        RECT 41.400 9.000 46.800 9.400 ;
        RECT 40.600 8.800 46.800 9.000 ;
        RECT 47.800 9.000 56.400 9.600 ;
        RECT 38.000 8.000 39.600 8.800 ;
        RECT 40.600 8.200 42.000 8.800 ;
        RECT 47.800 8.200 48.400 9.000 ;
        RECT 55.600 8.800 56.400 9.000 ;
        RECT 58.800 9.000 67.800 9.600 ;
        RECT 58.800 8.800 59.600 9.000 ;
        RECT 39.000 7.600 39.600 8.000 ;
        RECT 42.600 7.600 48.400 8.200 ;
        RECT 49.000 7.600 51.600 8.400 ;
        RECT 36.400 6.800 38.400 7.400 ;
        RECT 39.000 6.800 43.200 7.600 ;
        RECT 25.200 2.200 26.000 5.000 ;
        RECT 26.800 2.200 27.600 5.000 ;
        RECT 30.000 2.200 30.800 6.800 ;
        RECT 33.600 6.200 34.200 6.800 ;
        RECT 33.200 5.600 34.200 6.200 ;
        RECT 37.800 6.200 38.400 6.800 ;
        RECT 37.800 5.600 38.800 6.200 ;
        RECT 33.200 2.200 34.000 5.600 ;
        RECT 38.000 2.200 38.800 5.600 ;
        RECT 41.200 2.200 42.000 6.800 ;
        RECT 44.400 2.200 45.200 5.000 ;
        RECT 46.000 2.200 46.800 5.000 ;
        RECT 47.600 2.200 48.400 7.000 ;
        RECT 50.800 2.200 51.600 7.000 ;
        RECT 54.000 2.200 54.800 8.400 ;
        RECT 62.000 7.600 64.600 8.400 ;
        RECT 57.200 6.800 61.400 7.600 ;
        RECT 55.600 2.200 56.400 5.000 ;
        RECT 57.200 2.200 58.000 5.000 ;
        RECT 58.800 2.200 59.600 5.000 ;
        RECT 62.000 2.200 62.800 7.600 ;
        RECT 67.200 7.400 67.800 9.000 ;
        RECT 65.200 6.800 67.800 7.400 ;
        RECT 68.400 10.000 69.400 10.800 ;
        RECT 71.600 10.200 72.200 11.600 ;
        RECT 73.000 11.000 73.600 14.400 ;
        RECT 76.400 14.300 77.200 14.400 ;
        RECT 78.000 14.300 78.800 14.400 ;
        RECT 76.400 13.700 78.800 14.300 ;
        RECT 80.000 13.800 80.800 14.000 ;
        RECT 76.400 12.800 77.200 13.700 ;
        RECT 78.000 12.800 78.800 13.700 ;
        RECT 79.800 13.200 80.800 13.800 ;
        RECT 79.800 12.400 80.400 13.200 ;
        RECT 79.600 11.600 80.400 12.400 ;
        RECT 81.600 11.000 82.200 14.400 ;
        RECT 83.000 12.400 83.600 15.800 ;
        RECT 82.800 11.600 83.600 12.400 ;
        RECT 73.000 10.400 75.400 11.000 ;
        RECT 65.200 2.200 66.000 6.800 ;
        RECT 68.400 2.200 69.200 10.000 ;
        RECT 71.600 2.200 72.400 10.200 ;
        RECT 74.800 6.200 75.400 10.400 ;
        RECT 79.800 10.400 82.200 11.000 ;
        RECT 79.800 6.200 80.400 10.400 ;
        RECT 83.000 10.200 83.600 11.600 ;
        RECT 74.800 2.200 75.600 6.200 ;
        RECT 79.600 2.200 80.400 6.200 ;
        RECT 82.800 2.200 83.600 10.200 ;
        RECT 84.400 13.800 85.200 19.800 ;
        RECT 90.800 16.600 91.600 19.800 ;
        RECT 92.400 17.000 93.200 19.800 ;
        RECT 94.000 17.000 94.800 19.800 ;
        RECT 95.600 17.000 96.400 19.800 ;
        RECT 98.800 17.000 99.600 19.800 ;
        RECT 102.000 17.000 102.800 19.800 ;
        RECT 103.600 17.000 104.400 19.800 ;
        RECT 105.200 17.000 106.000 19.800 ;
        RECT 106.800 17.000 107.600 19.800 ;
        RECT 89.000 15.800 91.600 16.600 ;
        RECT 108.400 16.600 109.200 19.800 ;
        RECT 95.000 15.800 99.600 16.400 ;
        RECT 89.000 15.200 89.800 15.800 ;
        RECT 86.800 14.400 89.800 15.200 ;
        RECT 84.400 13.000 93.200 13.800 ;
        RECT 95.000 13.400 95.800 15.800 ;
        RECT 98.800 15.600 99.600 15.800 ;
        RECT 100.400 15.600 102.000 16.400 ;
        RECT 105.000 15.600 106.000 16.400 ;
        RECT 108.400 15.800 110.800 16.600 ;
        RECT 97.200 13.600 98.000 15.200 ;
        RECT 98.800 14.800 99.600 15.000 ;
        RECT 98.800 14.200 103.200 14.800 ;
        RECT 102.400 14.000 103.200 14.200 ;
        RECT 84.400 7.400 85.200 13.000 ;
        RECT 93.800 12.600 95.800 13.400 ;
        RECT 99.600 12.600 102.800 13.400 ;
        RECT 105.200 12.800 106.000 15.600 ;
        RECT 110.000 15.200 110.800 15.800 ;
        RECT 110.000 14.600 111.800 15.200 ;
        RECT 111.000 13.400 111.800 14.600 ;
        RECT 114.800 14.600 115.600 19.800 ;
        RECT 116.400 16.000 117.200 19.800 ;
        RECT 121.200 17.600 122.000 19.800 ;
        RECT 116.400 15.200 117.400 16.000 ;
        RECT 119.600 15.600 120.400 17.200 ;
        RECT 114.800 14.000 116.000 14.600 ;
        RECT 111.000 12.600 114.800 13.400 ;
        RECT 85.800 12.000 86.600 12.200 ;
        RECT 90.800 12.000 91.600 12.400 ;
        RECT 108.400 12.000 109.200 12.600 ;
        RECT 115.400 12.000 116.000 14.000 ;
        RECT 85.800 11.400 109.200 12.000 ;
        RECT 115.200 11.400 116.000 12.000 ;
        RECT 115.200 9.600 115.800 11.400 ;
        RECT 116.600 10.800 117.400 15.200 ;
        RECT 121.400 14.400 122.000 17.600 ;
        RECT 130.800 15.800 131.600 19.800 ;
        RECT 132.400 16.000 133.200 19.800 ;
        RECT 135.600 16.000 136.400 19.800 ;
        RECT 138.800 16.000 139.600 19.800 ;
        RECT 132.400 15.800 136.400 16.000 ;
        RECT 131.000 14.400 131.600 15.800 ;
        RECT 132.600 15.400 136.200 15.800 ;
        RECT 138.600 15.200 139.600 16.000 ;
        RECT 134.800 14.400 135.600 14.800 ;
        RECT 121.200 13.600 122.000 14.400 ;
        RECT 130.800 13.600 133.400 14.400 ;
        RECT 134.800 13.800 136.400 14.400 ;
        RECT 135.600 13.600 136.400 13.800 ;
        RECT 94.000 9.400 94.800 9.600 ;
        RECT 89.400 9.000 94.800 9.400 ;
        RECT 88.600 8.800 94.800 9.000 ;
        RECT 95.800 9.000 104.400 9.600 ;
        RECT 86.000 8.000 87.600 8.800 ;
        RECT 88.600 8.200 90.000 8.800 ;
        RECT 95.800 8.200 96.400 9.000 ;
        RECT 103.600 8.800 104.400 9.000 ;
        RECT 106.800 9.000 115.800 9.600 ;
        RECT 106.800 8.800 107.600 9.000 ;
        RECT 87.000 7.600 87.600 8.000 ;
        RECT 90.600 7.600 96.400 8.200 ;
        RECT 97.000 7.600 99.600 8.400 ;
        RECT 84.400 6.800 86.400 7.400 ;
        RECT 87.000 6.800 91.200 7.600 ;
        RECT 85.800 6.200 86.400 6.800 ;
        RECT 85.800 5.600 86.800 6.200 ;
        RECT 86.000 2.200 86.800 5.600 ;
        RECT 89.200 2.200 90.000 6.800 ;
        RECT 92.400 2.200 93.200 5.000 ;
        RECT 94.000 2.200 94.800 5.000 ;
        RECT 95.600 2.200 96.400 7.000 ;
        RECT 98.800 2.200 99.600 7.000 ;
        RECT 102.000 2.200 102.800 8.400 ;
        RECT 110.000 7.600 112.600 8.400 ;
        RECT 105.200 6.800 109.400 7.600 ;
        RECT 103.600 2.200 104.400 5.000 ;
        RECT 105.200 2.200 106.000 5.000 ;
        RECT 106.800 2.200 107.600 5.000 ;
        RECT 110.000 2.200 110.800 7.600 ;
        RECT 115.200 7.400 115.800 9.000 ;
        RECT 113.200 6.800 115.800 7.400 ;
        RECT 116.400 10.000 117.400 10.800 ;
        RECT 121.400 10.200 122.000 13.600 ;
        RECT 122.800 12.300 123.600 12.400 ;
        RECT 132.800 12.300 133.400 13.600 ;
        RECT 122.800 11.700 133.400 12.300 ;
        RECT 122.800 10.800 123.600 11.700 ;
        RECT 130.800 10.200 131.600 10.400 ;
        RECT 132.800 10.200 133.400 11.700 ;
        RECT 134.000 12.300 134.800 13.200 ;
        RECT 138.600 12.300 139.400 15.200 ;
        RECT 140.400 14.600 141.200 19.800 ;
        RECT 146.800 16.600 147.600 19.800 ;
        RECT 148.400 17.000 149.200 19.800 ;
        RECT 150.000 17.000 150.800 19.800 ;
        RECT 151.600 17.000 152.400 19.800 ;
        RECT 153.200 17.000 154.000 19.800 ;
        RECT 156.400 17.000 157.200 19.800 ;
        RECT 159.600 17.000 160.400 19.800 ;
        RECT 161.200 17.000 162.000 19.800 ;
        RECT 162.800 17.000 163.600 19.800 ;
        RECT 145.200 15.800 147.600 16.600 ;
        RECT 164.400 16.600 165.200 19.800 ;
        RECT 145.200 15.200 146.000 15.800 ;
        RECT 134.000 11.700 139.400 12.300 ;
        RECT 134.000 11.600 134.800 11.700 ;
        RECT 138.600 10.800 139.400 11.700 ;
        RECT 140.000 14.000 141.200 14.600 ;
        RECT 144.200 14.600 146.000 15.200 ;
        RECT 150.000 15.600 151.000 16.400 ;
        RECT 154.000 15.600 155.600 16.400 ;
        RECT 156.400 15.800 161.000 16.400 ;
        RECT 164.400 15.800 167.000 16.600 ;
        RECT 156.400 15.600 157.200 15.800 ;
        RECT 140.000 12.000 140.600 14.000 ;
        RECT 144.200 13.400 145.000 14.600 ;
        RECT 141.200 12.600 145.000 13.400 ;
        RECT 150.000 12.800 150.800 15.600 ;
        RECT 156.400 14.800 157.200 15.000 ;
        RECT 152.800 14.200 157.200 14.800 ;
        RECT 152.800 14.000 153.600 14.200 ;
        RECT 158.000 13.600 158.800 15.200 ;
        RECT 160.200 13.400 161.000 15.800 ;
        RECT 166.200 15.200 167.000 15.800 ;
        RECT 166.200 14.400 169.200 15.200 ;
        RECT 170.800 13.800 171.600 19.800 ;
        RECT 175.600 15.200 176.400 19.800 ;
        RECT 153.200 12.600 156.400 13.400 ;
        RECT 160.200 12.600 162.200 13.400 ;
        RECT 162.800 13.000 171.600 13.800 ;
        RECT 146.800 12.000 147.600 12.600 ;
        RECT 164.400 12.000 165.200 12.400 ;
        RECT 166.000 12.000 166.800 12.400 ;
        RECT 169.400 12.000 170.200 12.200 ;
        RECT 140.000 11.400 140.800 12.000 ;
        RECT 146.800 11.400 170.200 12.000 ;
        RECT 113.200 2.200 114.000 6.800 ;
        RECT 116.400 2.200 117.200 10.000 ;
        RECT 121.200 9.400 123.000 10.200 ;
        RECT 130.800 9.600 132.200 10.200 ;
        RECT 132.800 9.600 133.800 10.200 ;
        RECT 138.600 10.000 139.600 10.800 ;
        RECT 122.200 2.200 123.000 9.400 ;
        RECT 131.600 8.400 132.200 9.600 ;
        RECT 131.600 7.600 132.400 8.400 ;
        RECT 133.000 2.200 133.800 9.600 ;
        RECT 138.800 2.200 139.600 10.000 ;
        RECT 140.200 9.600 140.800 11.400 ;
        RECT 140.200 9.000 149.200 9.600 ;
        RECT 140.200 7.400 140.800 9.000 ;
        RECT 148.400 8.800 149.200 9.000 ;
        RECT 151.600 9.000 160.200 9.600 ;
        RECT 151.600 8.800 152.400 9.000 ;
        RECT 143.400 7.600 146.000 8.400 ;
        RECT 140.200 6.800 142.800 7.400 ;
        RECT 142.000 2.200 142.800 6.800 ;
        RECT 145.200 2.200 146.000 7.600 ;
        RECT 146.600 6.800 150.800 7.600 ;
        RECT 148.400 2.200 149.200 5.000 ;
        RECT 150.000 2.200 150.800 5.000 ;
        RECT 151.600 2.200 152.400 5.000 ;
        RECT 153.200 2.200 154.000 8.400 ;
        RECT 156.400 7.600 159.000 8.400 ;
        RECT 159.600 8.200 160.200 9.000 ;
        RECT 161.200 9.400 162.000 9.600 ;
        RECT 161.200 9.000 166.600 9.400 ;
        RECT 161.200 8.800 167.400 9.000 ;
        RECT 166.000 8.200 167.400 8.800 ;
        RECT 159.600 7.600 165.400 8.200 ;
        RECT 168.400 8.000 170.000 8.800 ;
        RECT 168.400 7.600 169.000 8.000 ;
        RECT 156.400 2.200 157.200 7.000 ;
        RECT 159.600 2.200 160.400 7.000 ;
        RECT 164.800 6.800 169.000 7.600 ;
        RECT 170.800 7.400 171.600 13.000 ;
        RECT 174.200 14.600 176.400 15.200 ;
        RECT 177.200 15.200 178.000 19.800 ;
        RECT 177.200 14.600 179.400 15.200 ;
        RECT 174.200 11.600 174.800 14.600 ;
        RECT 173.600 10.800 174.800 11.600 ;
        RECT 174.200 10.200 174.800 10.800 ;
        RECT 178.800 11.600 179.400 14.600 ;
        RECT 182.000 13.800 182.800 19.800 ;
        RECT 188.400 16.600 189.200 19.800 ;
        RECT 190.000 17.000 190.800 19.800 ;
        RECT 191.600 17.000 192.400 19.800 ;
        RECT 193.200 17.000 194.000 19.800 ;
        RECT 196.400 17.000 197.200 19.800 ;
        RECT 199.600 17.000 200.400 19.800 ;
        RECT 201.200 17.000 202.000 19.800 ;
        RECT 202.800 17.000 203.600 19.800 ;
        RECT 204.400 17.000 205.200 19.800 ;
        RECT 186.600 15.800 189.200 16.600 ;
        RECT 206.000 16.600 206.800 19.800 ;
        RECT 192.600 15.800 197.200 16.400 ;
        RECT 186.600 15.200 187.400 15.800 ;
        RECT 184.400 14.400 187.400 15.200 ;
        RECT 182.000 13.000 190.800 13.800 ;
        RECT 192.600 13.400 193.400 15.800 ;
        RECT 196.400 15.600 197.200 15.800 ;
        RECT 198.000 15.600 199.600 16.400 ;
        RECT 202.600 15.600 203.600 16.400 ;
        RECT 206.000 15.800 208.400 16.600 ;
        RECT 194.800 13.600 195.600 15.200 ;
        RECT 196.400 14.800 197.200 15.000 ;
        RECT 196.400 14.200 200.800 14.800 ;
        RECT 200.000 14.000 200.800 14.200 ;
        RECT 178.800 10.800 180.000 11.600 ;
        RECT 178.800 10.200 179.400 10.800 ;
        RECT 174.200 9.600 176.400 10.200 ;
        RECT 169.600 6.800 171.600 7.400 ;
        RECT 161.200 2.200 162.000 5.000 ;
        RECT 162.800 2.200 163.600 5.000 ;
        RECT 166.000 2.200 166.800 6.800 ;
        RECT 169.600 6.200 170.200 6.800 ;
        RECT 169.200 5.600 170.200 6.200 ;
        RECT 169.200 2.200 170.000 5.600 ;
        RECT 175.600 2.200 176.400 9.600 ;
        RECT 177.200 9.600 179.400 10.200 ;
        RECT 177.200 2.200 178.000 9.600 ;
        RECT 182.000 7.400 182.800 13.000 ;
        RECT 191.400 12.600 193.400 13.400 ;
        RECT 197.200 12.600 200.400 13.400 ;
        RECT 202.800 12.800 203.600 15.600 ;
        RECT 207.600 15.200 208.400 15.800 ;
        RECT 207.600 14.600 209.400 15.200 ;
        RECT 208.600 13.400 209.400 14.600 ;
        RECT 212.400 14.600 213.200 19.800 ;
        RECT 214.000 16.300 214.800 19.800 ;
        RECT 217.200 16.300 218.000 17.200 ;
        RECT 214.000 15.700 218.000 16.300 ;
        RECT 214.000 15.200 215.000 15.700 ;
        RECT 217.200 15.600 218.000 15.700 ;
        RECT 212.400 14.000 213.600 14.600 ;
        RECT 208.600 12.600 212.400 13.400 ;
        RECT 213.000 12.000 213.600 14.000 ;
        RECT 212.800 11.400 213.600 12.000 ;
        RECT 211.400 10.800 212.200 11.000 ;
        RECT 185.200 10.200 212.200 10.800 ;
        RECT 185.200 9.600 186.000 10.200 ;
        RECT 188.600 10.000 189.400 10.200 ;
        RECT 212.800 9.600 213.400 11.400 ;
        RECT 214.200 10.800 215.000 15.200 ;
        RECT 217.200 14.300 218.000 14.400 ;
        RECT 218.800 14.300 219.600 19.800 ;
        RECT 220.400 16.000 221.200 19.800 ;
        RECT 223.600 16.000 224.400 19.800 ;
        RECT 220.400 15.800 224.400 16.000 ;
        RECT 225.200 15.800 226.000 19.800 ;
        RECT 226.800 16.000 227.600 19.800 ;
        RECT 230.000 16.000 230.800 19.800 ;
        RECT 226.800 15.800 230.800 16.000 ;
        RECT 231.600 15.800 232.400 19.800 ;
        RECT 235.800 18.400 236.600 19.800 ;
        RECT 234.800 17.600 236.600 18.400 ;
        RECT 235.800 16.400 236.600 17.600 ;
        RECT 234.800 15.800 236.600 16.400 ;
        RECT 238.000 16.000 238.800 19.800 ;
        RECT 241.200 16.000 242.000 19.800 ;
        RECT 238.000 15.800 242.000 16.000 ;
        RECT 242.800 15.800 243.600 19.800 ;
        RECT 244.400 16.000 245.200 19.800 ;
        RECT 247.600 16.000 248.400 19.800 ;
        RECT 244.400 15.800 248.400 16.000 ;
        RECT 249.200 15.800 250.000 19.800 ;
        RECT 250.800 15.800 251.600 19.800 ;
        RECT 252.400 16.000 253.200 19.800 ;
        RECT 255.600 16.000 256.400 19.800 ;
        RECT 252.400 15.800 256.400 16.000 ;
        RECT 257.200 15.800 258.000 19.800 ;
        RECT 258.800 16.000 259.600 19.800 ;
        RECT 262.000 16.000 262.800 19.800 ;
        RECT 258.800 15.800 262.800 16.000 ;
        RECT 220.600 15.400 224.200 15.800 ;
        RECT 221.200 14.400 222.000 14.800 ;
        RECT 225.200 14.400 225.800 15.800 ;
        RECT 227.000 15.400 230.600 15.800 ;
        RECT 227.600 14.400 228.400 14.800 ;
        RECT 231.600 14.400 232.200 15.800 ;
        RECT 220.400 14.300 222.000 14.400 ;
        RECT 217.200 13.800 222.000 14.300 ;
        RECT 217.200 13.700 221.200 13.800 ;
        RECT 217.200 13.600 218.000 13.700 ;
        RECT 191.600 9.400 192.400 9.600 ;
        RECT 187.000 9.000 192.400 9.400 ;
        RECT 186.200 8.800 192.400 9.000 ;
        RECT 193.400 9.000 202.000 9.600 ;
        RECT 183.600 8.000 185.200 8.800 ;
        RECT 186.200 8.200 187.600 8.800 ;
        RECT 193.400 8.200 194.000 9.000 ;
        RECT 201.200 8.800 202.000 9.000 ;
        RECT 204.400 9.000 213.400 9.600 ;
        RECT 204.400 8.800 205.200 9.000 ;
        RECT 184.600 7.600 185.200 8.000 ;
        RECT 188.200 7.600 194.000 8.200 ;
        RECT 194.600 7.600 197.200 8.400 ;
        RECT 182.000 6.800 184.000 7.400 ;
        RECT 184.600 6.800 188.800 7.600 ;
        RECT 183.400 6.200 184.000 6.800 ;
        RECT 183.400 5.600 184.400 6.200 ;
        RECT 183.600 2.200 184.400 5.600 ;
        RECT 186.800 2.200 187.600 6.800 ;
        RECT 190.000 2.200 190.800 5.000 ;
        RECT 191.600 2.200 192.400 5.000 ;
        RECT 193.200 2.200 194.000 7.000 ;
        RECT 196.400 2.200 197.200 7.000 ;
        RECT 199.600 2.200 200.400 8.400 ;
        RECT 207.600 7.600 210.200 8.400 ;
        RECT 202.800 6.800 207.000 7.600 ;
        RECT 201.200 2.200 202.000 5.000 ;
        RECT 202.800 2.200 203.600 5.000 ;
        RECT 204.400 2.200 205.200 5.000 ;
        RECT 207.600 2.200 208.400 7.600 ;
        RECT 212.800 7.400 213.400 9.000 ;
        RECT 210.800 6.800 213.400 7.400 ;
        RECT 214.000 10.000 215.000 10.800 ;
        RECT 210.800 2.200 211.600 6.800 ;
        RECT 214.000 2.200 214.800 10.000 ;
        RECT 218.800 2.200 219.600 13.700 ;
        RECT 220.400 13.600 221.200 13.700 ;
        RECT 223.400 13.600 226.000 14.400 ;
        RECT 226.800 13.800 228.400 14.400 ;
        RECT 226.800 13.600 227.600 13.800 ;
        RECT 229.800 13.600 232.400 14.400 ;
        RECT 233.200 13.600 234.000 15.200 ;
        RECT 222.000 11.600 222.800 13.200 ;
        RECT 223.400 10.200 224.000 13.600 ;
        RECT 225.200 12.300 226.000 12.400 ;
        RECT 228.400 12.300 229.200 13.200 ;
        RECT 225.200 11.700 229.200 12.300 ;
        RECT 225.200 11.600 226.000 11.700 ;
        RECT 228.400 11.600 229.200 11.700 ;
        RECT 225.200 10.200 226.000 10.400 ;
        RECT 229.800 10.200 230.400 13.600 ;
        RECT 231.600 10.200 232.400 10.400 ;
        RECT 223.000 9.600 224.000 10.200 ;
        RECT 224.600 9.600 226.000 10.200 ;
        RECT 229.400 9.600 230.400 10.200 ;
        RECT 231.000 9.600 232.400 10.200 ;
        RECT 223.000 2.200 223.800 9.600 ;
        RECT 224.600 8.400 225.200 9.600 ;
        RECT 229.400 8.400 230.200 9.600 ;
        RECT 231.000 8.400 231.600 9.600 ;
        RECT 224.400 7.600 225.200 8.400 ;
        RECT 228.400 7.600 230.200 8.400 ;
        RECT 230.800 7.600 231.600 8.400 ;
        RECT 229.400 2.200 230.200 7.600 ;
        RECT 234.800 2.200 235.600 15.800 ;
        RECT 238.200 15.400 241.800 15.800 ;
        RECT 238.800 14.400 239.600 14.800 ;
        RECT 242.800 14.400 243.400 15.800 ;
        RECT 244.600 15.400 248.200 15.800 ;
        RECT 245.200 14.400 246.000 14.800 ;
        RECT 249.200 14.400 249.800 15.800 ;
        RECT 251.000 14.400 251.600 15.800 ;
        RECT 252.600 15.400 256.200 15.800 ;
        RECT 254.800 14.400 255.600 14.800 ;
        RECT 257.400 14.400 258.000 15.800 ;
        RECT 259.000 15.400 262.600 15.800 ;
        RECT 261.200 14.400 262.000 14.800 ;
        RECT 238.000 13.800 239.600 14.400 ;
        RECT 238.000 13.600 238.800 13.800 ;
        RECT 241.000 13.600 243.600 14.400 ;
        RECT 244.400 13.800 246.000 14.400 ;
        RECT 244.400 13.600 245.200 13.800 ;
        RECT 247.400 13.600 250.000 14.400 ;
        RECT 250.800 13.600 253.400 14.400 ;
        RECT 254.800 13.800 256.400 14.400 ;
        RECT 255.600 13.600 256.400 13.800 ;
        RECT 257.200 13.600 259.800 14.400 ;
        RECT 261.200 13.800 262.800 14.400 ;
        RECT 262.000 13.600 262.800 13.800 ;
        RECT 239.600 11.600 240.400 13.200 ;
        RECT 236.400 8.800 237.200 10.400 ;
        RECT 241.000 10.200 241.600 13.600 ;
        RECT 246.000 11.600 246.800 13.200 ;
        RECT 247.400 12.300 248.000 13.600 ;
        RECT 247.400 11.700 251.500 12.300 ;
        RECT 242.800 10.200 243.600 10.400 ;
        RECT 247.400 10.200 248.000 11.700 ;
        RECT 250.900 10.400 251.500 11.700 ;
        RECT 249.200 10.200 250.000 10.400 ;
        RECT 240.600 9.600 241.600 10.200 ;
        RECT 242.200 9.600 243.600 10.200 ;
        RECT 247.000 9.600 248.000 10.200 ;
        RECT 248.600 9.600 250.000 10.200 ;
        RECT 250.800 10.200 251.600 10.400 ;
        RECT 252.800 10.200 253.400 13.600 ;
        RECT 254.000 11.600 254.800 13.200 ;
        RECT 255.600 12.300 256.400 12.400 ;
        RECT 259.200 12.300 259.800 13.600 ;
        RECT 255.600 11.700 259.800 12.300 ;
        RECT 255.600 11.600 256.400 11.700 ;
        RECT 257.200 10.200 258.000 10.400 ;
        RECT 259.200 10.200 259.800 11.700 ;
        RECT 260.400 12.300 261.200 13.200 ;
        RECT 262.000 12.300 262.800 12.400 ;
        RECT 260.400 11.700 262.800 12.300 ;
        RECT 260.400 11.600 261.200 11.700 ;
        RECT 262.000 11.600 262.800 11.700 ;
        RECT 250.800 9.600 252.200 10.200 ;
        RECT 252.800 9.600 253.800 10.200 ;
        RECT 257.200 9.600 258.600 10.200 ;
        RECT 259.200 9.600 260.200 10.200 ;
        RECT 240.600 8.400 241.400 9.600 ;
        RECT 242.200 8.400 242.800 9.600 ;
        RECT 239.600 7.600 241.400 8.400 ;
        RECT 242.000 7.600 242.800 8.400 ;
        RECT 240.600 2.200 241.400 7.600 ;
        RECT 247.000 2.200 247.800 9.600 ;
        RECT 248.600 8.400 249.200 9.600 ;
        RECT 248.400 7.600 249.200 8.400 ;
        RECT 251.600 8.400 252.200 9.600 ;
        RECT 253.000 8.400 253.800 9.600 ;
        RECT 258.000 8.400 258.600 9.600 ;
        RECT 251.600 7.600 252.400 8.400 ;
        RECT 253.000 7.600 254.800 8.400 ;
        RECT 258.000 7.600 258.800 8.400 ;
        RECT 253.000 2.200 253.800 7.600 ;
        RECT 259.400 2.200 260.200 9.600 ;
        RECT 263.600 2.200 264.400 19.800 ;
        RECT 265.200 15.600 266.000 17.200 ;
        RECT 266.800 15.600 267.600 17.200 ;
        RECT 265.200 10.300 266.000 10.400 ;
        RECT 268.400 10.300 269.200 19.800 ;
        RECT 270.000 16.000 270.800 19.800 ;
        RECT 273.200 16.000 274.000 19.800 ;
        RECT 270.000 15.800 274.000 16.000 ;
        RECT 274.800 15.800 275.600 19.800 ;
        RECT 282.800 16.000 283.600 19.800 ;
        RECT 286.000 16.000 286.800 19.800 ;
        RECT 282.800 15.800 286.800 16.000 ;
        RECT 287.600 15.800 288.400 19.800 ;
        RECT 290.800 16.000 291.600 19.800 ;
        RECT 270.200 15.400 273.800 15.800 ;
        RECT 270.800 14.400 271.600 14.800 ;
        RECT 274.800 14.400 275.400 15.800 ;
        RECT 283.000 15.400 286.600 15.800 ;
        RECT 283.600 14.400 284.400 14.800 ;
        RECT 287.600 14.400 288.200 15.800 ;
        RECT 290.600 15.200 291.600 16.000 ;
        RECT 270.000 13.800 271.600 14.400 ;
        RECT 273.000 14.300 275.600 14.400 ;
        RECT 278.000 14.300 278.800 14.400 ;
        RECT 270.000 13.600 270.800 13.800 ;
        RECT 273.000 13.700 278.800 14.300 ;
        RECT 273.000 13.600 275.600 13.700 ;
        RECT 278.000 13.600 278.800 13.700 ;
        RECT 279.600 14.300 280.400 14.400 ;
        RECT 282.800 14.300 284.400 14.400 ;
        RECT 279.600 13.800 284.400 14.300 ;
        RECT 279.600 13.700 283.600 13.800 ;
        RECT 279.600 13.600 280.400 13.700 ;
        RECT 282.800 13.600 283.600 13.700 ;
        RECT 285.800 13.600 288.400 14.400 ;
        RECT 271.600 11.600 272.400 13.200 ;
        RECT 265.200 9.700 269.200 10.300 ;
        RECT 273.000 10.200 273.600 13.600 ;
        RECT 281.200 12.300 282.000 12.400 ;
        RECT 284.400 12.300 285.200 13.200 ;
        RECT 274.900 11.700 285.200 12.300 ;
        RECT 274.900 10.400 275.500 11.700 ;
        RECT 281.200 11.600 282.000 11.700 ;
        RECT 284.400 11.600 285.200 11.700 ;
        RECT 274.800 10.200 275.600 10.400 ;
        RECT 285.800 10.200 286.400 13.600 ;
        RECT 290.600 10.800 291.400 15.200 ;
        RECT 292.400 14.600 293.200 19.800 ;
        RECT 298.800 16.600 299.600 19.800 ;
        RECT 300.400 17.000 301.200 19.800 ;
        RECT 302.000 17.000 302.800 19.800 ;
        RECT 303.600 17.000 304.400 19.800 ;
        RECT 305.200 17.000 306.000 19.800 ;
        RECT 308.400 17.000 309.200 19.800 ;
        RECT 311.600 17.000 312.400 19.800 ;
        RECT 313.200 17.000 314.000 19.800 ;
        RECT 314.800 17.000 315.600 19.800 ;
        RECT 297.200 15.800 299.600 16.600 ;
        RECT 316.400 16.600 317.200 19.800 ;
        RECT 297.200 15.200 298.000 15.800 ;
        RECT 292.000 14.000 293.200 14.600 ;
        RECT 296.200 14.600 298.000 15.200 ;
        RECT 302.000 15.600 303.000 16.400 ;
        RECT 306.000 15.600 307.600 16.400 ;
        RECT 308.400 15.800 313.000 16.400 ;
        RECT 316.400 15.800 319.000 16.600 ;
        RECT 308.400 15.600 309.200 15.800 ;
        RECT 292.000 12.000 292.600 14.000 ;
        RECT 296.200 13.400 297.000 14.600 ;
        RECT 293.200 12.600 297.000 13.400 ;
        RECT 302.000 12.800 302.800 15.600 ;
        RECT 308.400 14.800 309.200 15.000 ;
        RECT 304.800 14.200 309.200 14.800 ;
        RECT 304.800 14.000 305.600 14.200 ;
        RECT 310.000 13.600 310.800 15.200 ;
        RECT 312.200 13.400 313.000 15.800 ;
        RECT 318.200 15.200 319.000 15.800 ;
        RECT 318.200 14.400 321.200 15.200 ;
        RECT 322.800 13.800 323.600 19.800 ;
        RECT 324.400 15.800 325.200 19.800 ;
        RECT 328.600 16.800 329.400 19.800 ;
        RECT 328.600 15.800 330.000 16.800 ;
        RECT 330.800 15.800 331.600 19.800 ;
        RECT 335.000 18.400 335.800 19.800 ;
        RECT 335.000 17.600 336.400 18.400 ;
        RECT 335.000 16.800 335.800 17.600 ;
        RECT 335.000 15.800 336.400 16.800 ;
        RECT 338.800 16.000 339.600 19.800 ;
        RECT 324.600 15.600 325.200 15.800 ;
        RECT 324.600 15.200 326.400 15.600 ;
        RECT 324.600 15.000 328.800 15.200 ;
        RECT 325.800 14.600 328.800 15.000 ;
        RECT 328.000 14.400 328.800 14.600 ;
        RECT 305.200 12.600 308.400 13.400 ;
        RECT 312.200 12.600 314.200 13.400 ;
        RECT 314.800 13.000 323.600 13.800 ;
        RECT 292.000 11.400 292.800 12.000 ;
        RECT 287.600 10.200 288.400 10.400 ;
        RECT 265.200 9.600 266.000 9.700 ;
        RECT 268.400 2.200 269.200 9.700 ;
        RECT 272.600 9.600 273.600 10.200 ;
        RECT 274.200 9.600 275.600 10.200 ;
        RECT 285.400 9.600 286.400 10.200 ;
        RECT 287.000 9.600 288.400 10.200 ;
        RECT 290.600 10.000 291.600 10.800 ;
        RECT 272.600 2.200 273.400 9.600 ;
        RECT 274.200 8.400 274.800 9.600 ;
        RECT 274.000 7.600 274.800 8.400 ;
        RECT 285.400 2.200 286.200 9.600 ;
        RECT 287.000 8.400 287.600 9.600 ;
        RECT 286.800 7.600 287.600 8.400 ;
        RECT 290.800 2.200 291.600 10.000 ;
        RECT 292.200 9.600 292.800 11.400 ;
        RECT 293.400 10.800 294.200 11.000 ;
        RECT 293.400 10.300 320.400 10.800 ;
        RECT 321.200 10.300 322.000 10.400 ;
        RECT 293.400 10.200 322.000 10.300 ;
        RECT 316.200 10.000 317.000 10.200 ;
        RECT 319.600 9.700 322.000 10.200 ;
        RECT 319.600 9.600 320.400 9.700 ;
        RECT 321.200 9.600 322.000 9.700 ;
        RECT 292.200 9.000 301.200 9.600 ;
        RECT 292.200 7.400 292.800 9.000 ;
        RECT 300.400 8.800 301.200 9.000 ;
        RECT 303.600 9.000 312.200 9.600 ;
        RECT 303.600 8.800 304.400 9.000 ;
        RECT 295.400 7.600 298.000 8.400 ;
        RECT 292.200 6.800 294.800 7.400 ;
        RECT 294.000 2.200 294.800 6.800 ;
        RECT 297.200 2.200 298.000 7.600 ;
        RECT 298.600 6.800 302.800 7.600 ;
        RECT 300.400 2.200 301.200 5.000 ;
        RECT 302.000 2.200 302.800 5.000 ;
        RECT 303.600 2.200 304.400 5.000 ;
        RECT 305.200 2.200 306.000 8.400 ;
        RECT 308.400 7.600 311.000 8.400 ;
        RECT 311.600 8.200 312.200 9.000 ;
        RECT 313.200 9.400 314.000 9.600 ;
        RECT 313.200 9.000 318.600 9.400 ;
        RECT 313.200 8.800 319.400 9.000 ;
        RECT 318.000 8.200 319.400 8.800 ;
        RECT 311.600 7.600 317.400 8.200 ;
        RECT 320.400 8.000 322.000 8.800 ;
        RECT 320.400 7.600 321.000 8.000 ;
        RECT 308.400 2.200 309.200 7.000 ;
        RECT 311.600 2.200 312.400 7.000 ;
        RECT 316.800 6.800 321.000 7.600 ;
        RECT 322.800 7.400 323.600 13.000 ;
        RECT 324.400 12.800 325.200 14.400 ;
        RECT 328.000 11.000 328.600 14.400 ;
        RECT 329.400 12.400 330.000 15.800 ;
        RECT 331.000 15.600 331.600 15.800 ;
        RECT 331.000 15.200 332.800 15.600 ;
        RECT 331.000 15.000 335.200 15.200 ;
        RECT 332.200 14.600 335.200 15.000 ;
        RECT 334.400 14.400 335.200 14.600 ;
        RECT 330.800 12.800 331.600 14.400 ;
        RECT 332.800 13.800 333.600 14.000 ;
        RECT 332.600 13.200 333.600 13.800 ;
        RECT 332.600 12.400 333.200 13.200 ;
        RECT 329.200 11.600 330.000 12.400 ;
        RECT 332.400 11.600 333.200 12.400 ;
        RECT 321.600 6.800 323.600 7.400 ;
        RECT 326.200 10.400 328.600 11.000 ;
        RECT 313.200 2.200 314.000 5.000 ;
        RECT 314.800 2.200 315.600 5.000 ;
        RECT 318.000 2.200 318.800 6.800 ;
        RECT 321.600 6.200 322.200 6.800 ;
        RECT 326.200 6.200 326.800 10.400 ;
        RECT 329.400 10.200 330.000 11.600 ;
        RECT 334.400 11.000 335.000 14.400 ;
        RECT 335.800 12.400 336.400 15.800 ;
        RECT 335.600 11.600 336.400 12.400 ;
        RECT 321.200 5.600 322.200 6.200 ;
        RECT 321.200 2.200 322.000 5.600 ;
        RECT 326.000 2.200 326.800 6.200 ;
        RECT 329.200 2.200 330.000 10.200 ;
        RECT 332.600 10.400 335.000 11.000 ;
        RECT 332.600 6.200 333.200 10.400 ;
        RECT 335.800 10.200 336.400 11.600 ;
        RECT 332.400 2.200 333.200 6.200 ;
        RECT 335.600 2.200 336.400 10.200 ;
        RECT 338.600 15.200 339.600 16.000 ;
        RECT 338.600 10.800 339.400 15.200 ;
        RECT 340.400 14.600 341.200 19.800 ;
        RECT 346.800 16.600 347.600 19.800 ;
        RECT 348.400 17.000 349.200 19.800 ;
        RECT 350.000 17.000 350.800 19.800 ;
        RECT 351.600 17.000 352.400 19.800 ;
        RECT 353.200 17.000 354.000 19.800 ;
        RECT 356.400 17.000 357.200 19.800 ;
        RECT 359.600 17.000 360.400 19.800 ;
        RECT 361.200 17.000 362.000 19.800 ;
        RECT 362.800 17.000 363.600 19.800 ;
        RECT 345.200 15.800 347.600 16.600 ;
        RECT 364.400 16.600 365.200 19.800 ;
        RECT 345.200 15.200 346.000 15.800 ;
        RECT 340.000 14.000 341.200 14.600 ;
        RECT 344.200 14.600 346.000 15.200 ;
        RECT 350.000 15.600 351.000 16.400 ;
        RECT 354.000 15.600 355.600 16.400 ;
        RECT 356.400 15.800 361.000 16.400 ;
        RECT 364.400 15.800 367.000 16.600 ;
        RECT 356.400 15.600 357.200 15.800 ;
        RECT 340.000 12.000 340.600 14.000 ;
        RECT 344.200 13.400 345.000 14.600 ;
        RECT 341.200 12.600 345.000 13.400 ;
        RECT 350.000 12.800 350.800 15.600 ;
        RECT 356.400 14.800 357.200 15.000 ;
        RECT 352.800 14.200 357.200 14.800 ;
        RECT 352.800 14.000 353.600 14.200 ;
        RECT 358.000 13.600 358.800 15.200 ;
        RECT 360.200 13.400 361.000 15.800 ;
        RECT 366.200 15.200 367.000 15.800 ;
        RECT 366.200 14.400 369.200 15.200 ;
        RECT 370.800 13.800 371.600 19.800 ;
        RECT 375.600 15.200 376.400 19.800 ;
        RECT 353.200 12.600 356.400 13.400 ;
        RECT 360.200 12.600 362.200 13.400 ;
        RECT 362.800 13.000 371.600 13.800 ;
        RECT 346.800 12.000 347.600 12.600 ;
        RECT 364.400 12.000 365.200 12.400 ;
        RECT 367.600 12.000 368.400 12.400 ;
        RECT 369.400 12.000 370.200 12.200 ;
        RECT 340.000 11.400 340.800 12.000 ;
        RECT 346.800 11.400 370.200 12.000 ;
        RECT 338.600 10.000 339.600 10.800 ;
        RECT 338.800 2.200 339.600 10.000 ;
        RECT 340.200 9.600 340.800 11.400 ;
        RECT 340.200 9.000 349.200 9.600 ;
        RECT 340.200 7.400 340.800 9.000 ;
        RECT 348.400 8.800 349.200 9.000 ;
        RECT 351.600 9.000 360.200 9.600 ;
        RECT 351.600 8.800 352.400 9.000 ;
        RECT 343.400 7.600 346.000 8.400 ;
        RECT 340.200 6.800 342.800 7.400 ;
        RECT 342.000 2.200 342.800 6.800 ;
        RECT 345.200 2.200 346.000 7.600 ;
        RECT 346.600 6.800 350.800 7.600 ;
        RECT 348.400 2.200 349.200 5.000 ;
        RECT 350.000 2.200 350.800 5.000 ;
        RECT 351.600 2.200 352.400 5.000 ;
        RECT 353.200 2.200 354.000 8.400 ;
        RECT 356.400 7.600 359.000 8.400 ;
        RECT 359.600 8.200 360.200 9.000 ;
        RECT 361.200 9.400 362.000 9.600 ;
        RECT 361.200 9.000 366.600 9.400 ;
        RECT 361.200 8.800 367.400 9.000 ;
        RECT 366.000 8.200 367.400 8.800 ;
        RECT 359.600 7.600 365.400 8.200 ;
        RECT 368.400 8.000 370.000 8.800 ;
        RECT 368.400 7.600 369.000 8.000 ;
        RECT 356.400 2.200 357.200 7.000 ;
        RECT 359.600 2.200 360.400 7.000 ;
        RECT 364.800 6.800 369.000 7.600 ;
        RECT 370.800 7.400 371.600 13.000 ;
        RECT 374.200 14.600 376.400 15.200 ;
        RECT 377.200 15.400 378.000 19.800 ;
        RECT 381.400 18.400 382.600 19.800 ;
        RECT 381.400 17.800 382.800 18.400 ;
        RECT 386.000 17.800 386.800 19.800 ;
        RECT 390.400 18.400 391.200 19.800 ;
        RECT 390.400 17.800 392.400 18.400 ;
        RECT 382.000 17.000 382.800 17.800 ;
        RECT 386.200 17.200 386.800 17.800 ;
        RECT 386.200 16.600 389.000 17.200 ;
        RECT 388.200 16.400 389.000 16.600 ;
        RECT 390.000 16.400 390.800 17.200 ;
        RECT 391.600 17.000 392.400 17.800 ;
        RECT 380.200 15.400 381.000 15.600 ;
        RECT 377.200 14.800 381.000 15.400 ;
        RECT 374.200 11.600 374.800 14.600 ;
        RECT 375.600 12.300 376.400 13.200 ;
        RECT 377.200 12.300 378.000 14.800 ;
        RECT 384.200 14.200 385.000 14.400 ;
        RECT 386.800 14.200 387.600 14.400 ;
        RECT 390.000 14.200 390.600 16.400 ;
        RECT 394.800 15.000 395.600 19.800 ;
        RECT 393.200 14.200 394.800 14.400 ;
        RECT 383.800 13.600 394.800 14.200 ;
        RECT 396.400 13.800 397.200 19.800 ;
        RECT 402.800 16.600 403.600 19.800 ;
        RECT 404.400 17.000 405.200 19.800 ;
        RECT 406.000 17.000 406.800 19.800 ;
        RECT 407.600 17.000 408.400 19.800 ;
        RECT 410.800 17.000 411.600 19.800 ;
        RECT 414.000 17.000 414.800 19.800 ;
        RECT 415.600 17.000 416.400 19.800 ;
        RECT 417.200 17.000 418.000 19.800 ;
        RECT 418.800 17.000 419.600 19.800 ;
        RECT 401.000 15.800 403.600 16.600 ;
        RECT 420.400 16.600 421.200 19.800 ;
        RECT 407.000 15.800 411.600 16.400 ;
        RECT 401.000 15.200 401.800 15.800 ;
        RECT 398.800 14.400 401.800 15.200 ;
        RECT 382.000 12.800 382.800 13.000 ;
        RECT 375.600 11.700 378.000 12.300 ;
        RECT 379.000 12.200 382.800 12.800 ;
        RECT 379.000 12.000 379.800 12.200 ;
        RECT 375.600 11.600 376.400 11.700 ;
        RECT 373.600 10.800 374.800 11.600 ;
        RECT 374.200 10.200 374.800 10.800 ;
        RECT 377.200 11.400 378.000 11.700 ;
        RECT 380.600 11.400 381.400 11.600 ;
        RECT 377.200 10.800 381.400 11.400 ;
        RECT 374.200 9.600 376.400 10.200 ;
        RECT 369.600 6.800 371.600 7.400 ;
        RECT 361.200 2.200 362.000 5.000 ;
        RECT 362.800 2.200 363.600 5.000 ;
        RECT 366.000 2.200 366.800 6.800 ;
        RECT 369.600 6.200 370.200 6.800 ;
        RECT 369.200 5.600 370.200 6.200 ;
        RECT 369.200 2.200 370.000 5.600 ;
        RECT 375.600 2.200 376.400 9.600 ;
        RECT 377.200 2.200 378.000 10.800 ;
        RECT 383.800 10.400 384.400 13.600 ;
        RECT 391.000 13.400 391.800 13.600 ;
        RECT 396.400 13.000 405.200 13.800 ;
        RECT 407.000 13.400 407.800 15.800 ;
        RECT 410.800 15.600 411.600 15.800 ;
        RECT 412.400 15.600 414.000 16.400 ;
        RECT 417.000 15.600 418.000 16.400 ;
        RECT 420.400 15.800 422.800 16.600 ;
        RECT 409.200 13.600 410.000 15.200 ;
        RECT 410.800 14.800 411.600 15.000 ;
        RECT 410.800 14.200 415.200 14.800 ;
        RECT 414.400 14.000 415.200 14.200 ;
        RECT 390.000 12.400 390.800 12.600 ;
        RECT 392.600 12.400 393.400 12.600 ;
        RECT 388.400 11.800 393.400 12.400 ;
        RECT 388.400 11.600 389.200 11.800 ;
        RECT 390.000 11.000 395.600 11.200 ;
        RECT 389.800 10.800 395.600 11.000 ;
        RECT 382.000 9.800 384.400 10.400 ;
        RECT 385.800 10.600 395.600 10.800 ;
        RECT 385.800 10.200 390.600 10.600 ;
        RECT 382.000 8.800 382.600 9.800 ;
        RECT 381.200 8.000 382.600 8.800 ;
        RECT 384.200 9.000 385.000 9.200 ;
        RECT 385.800 9.000 386.400 10.200 ;
        RECT 384.200 8.400 386.400 9.000 ;
        RECT 387.000 9.000 392.400 9.600 ;
        RECT 387.000 8.800 387.800 9.000 ;
        RECT 391.600 8.800 392.400 9.000 ;
        RECT 385.400 7.400 386.200 7.600 ;
        RECT 388.200 7.400 389.000 7.600 ;
        RECT 382.000 6.200 382.800 7.000 ;
        RECT 385.400 6.800 389.000 7.400 ;
        RECT 386.200 6.200 386.800 6.800 ;
        RECT 391.600 6.200 392.400 7.000 ;
        RECT 381.400 2.200 382.600 6.200 ;
        RECT 386.000 2.200 386.800 6.200 ;
        RECT 390.400 5.600 392.400 6.200 ;
        RECT 390.400 2.200 391.200 5.600 ;
        RECT 394.800 2.200 395.600 10.600 ;
        RECT 396.400 7.400 397.200 13.000 ;
        RECT 405.800 12.600 407.800 13.400 ;
        RECT 411.600 12.600 414.800 13.400 ;
        RECT 417.200 12.800 418.000 15.600 ;
        RECT 422.000 15.200 422.800 15.800 ;
        RECT 422.000 14.600 423.800 15.200 ;
        RECT 423.000 13.400 423.800 14.600 ;
        RECT 426.800 14.600 427.600 19.800 ;
        RECT 428.400 16.000 429.200 19.800 ;
        RECT 428.400 15.200 429.400 16.000 ;
        RECT 426.800 14.000 428.000 14.600 ;
        RECT 423.000 12.600 426.800 13.400 ;
        RECT 397.800 12.000 398.600 12.200 ;
        RECT 399.600 12.000 400.400 12.400 ;
        RECT 402.800 12.000 403.600 12.400 ;
        RECT 420.400 12.000 421.200 12.600 ;
        RECT 427.400 12.000 428.000 14.000 ;
        RECT 397.800 11.400 421.200 12.000 ;
        RECT 427.200 11.400 428.000 12.000 ;
        RECT 427.200 9.600 427.800 11.400 ;
        RECT 428.600 10.800 429.400 15.200 ;
        RECT 438.000 15.000 438.800 19.800 ;
        RECT 442.400 18.400 443.200 19.800 ;
        RECT 441.200 17.800 443.200 18.400 ;
        RECT 446.800 17.800 447.600 19.800 ;
        RECT 451.000 18.400 452.200 19.800 ;
        RECT 450.800 17.800 452.200 18.400 ;
        RECT 441.200 17.000 442.000 17.800 ;
        RECT 446.800 17.200 447.400 17.800 ;
        RECT 442.800 16.400 443.600 17.200 ;
        RECT 444.600 16.600 447.400 17.200 ;
        RECT 450.800 17.000 451.600 17.800 ;
        RECT 444.600 16.400 445.400 16.600 ;
        RECT 438.800 14.200 440.400 14.400 ;
        RECT 443.000 14.200 443.600 16.400 ;
        RECT 452.600 15.400 453.400 15.600 ;
        RECT 455.600 15.400 456.400 19.800 ;
        RECT 452.600 14.800 456.400 15.400 ;
        RECT 448.600 14.200 449.400 14.400 ;
        RECT 438.800 13.600 449.800 14.200 ;
        RECT 441.800 13.400 442.600 13.600 ;
        RECT 440.200 12.400 441.000 12.600 ;
        RECT 442.800 12.400 443.600 12.600 ;
        RECT 449.200 12.400 449.800 13.600 ;
        RECT 450.800 12.800 451.600 13.000 ;
        RECT 440.200 11.800 445.200 12.400 ;
        RECT 444.400 11.600 445.200 11.800 ;
        RECT 449.200 11.600 450.000 12.400 ;
        RECT 450.800 12.200 454.600 12.800 ;
        RECT 453.800 12.000 454.600 12.200 ;
        RECT 455.600 12.300 456.400 14.800 ;
        RECT 457.200 15.200 458.000 19.800 ;
        RECT 462.000 15.200 462.800 19.800 ;
        RECT 457.200 14.600 459.400 15.200 ;
        RECT 462.000 14.600 464.200 15.200 ;
        RECT 457.200 12.300 458.000 13.200 ;
        RECT 455.600 11.700 458.000 12.300 ;
        RECT 406.000 9.400 406.800 9.600 ;
        RECT 401.400 9.000 406.800 9.400 ;
        RECT 400.600 8.800 406.800 9.000 ;
        RECT 407.800 9.000 416.400 9.600 ;
        RECT 398.000 8.000 399.600 8.800 ;
        RECT 400.600 8.200 402.000 8.800 ;
        RECT 407.800 8.200 408.400 9.000 ;
        RECT 415.600 8.800 416.400 9.000 ;
        RECT 418.800 9.000 427.800 9.600 ;
        RECT 418.800 8.800 419.600 9.000 ;
        RECT 399.000 7.600 399.600 8.000 ;
        RECT 402.600 7.600 408.400 8.200 ;
        RECT 409.000 7.600 411.600 8.400 ;
        RECT 396.400 6.800 398.400 7.400 ;
        RECT 399.000 6.800 403.200 7.600 ;
        RECT 397.800 6.200 398.400 6.800 ;
        RECT 397.800 5.600 398.800 6.200 ;
        RECT 398.000 2.200 398.800 5.600 ;
        RECT 401.200 2.200 402.000 6.800 ;
        RECT 404.400 2.200 405.200 5.000 ;
        RECT 406.000 2.200 406.800 5.000 ;
        RECT 407.600 2.200 408.400 7.000 ;
        RECT 410.800 2.200 411.600 7.000 ;
        RECT 414.000 2.200 414.800 8.400 ;
        RECT 422.000 7.600 424.600 8.400 ;
        RECT 417.200 6.800 421.400 7.600 ;
        RECT 415.600 2.200 416.400 5.000 ;
        RECT 417.200 2.200 418.000 5.000 ;
        RECT 418.800 2.200 419.600 5.000 ;
        RECT 422.000 2.200 422.800 7.600 ;
        RECT 427.200 7.400 427.800 9.000 ;
        RECT 425.200 6.800 427.800 7.400 ;
        RECT 428.400 10.000 429.400 10.800 ;
        RECT 438.000 11.000 443.600 11.200 ;
        RECT 438.000 10.800 443.800 11.000 ;
        RECT 438.000 10.600 447.800 10.800 ;
        RECT 425.200 2.200 426.000 6.800 ;
        RECT 428.400 2.200 429.200 10.000 ;
        RECT 438.000 2.200 438.800 10.600 ;
        RECT 443.000 10.200 447.800 10.600 ;
        RECT 441.200 9.000 446.600 9.600 ;
        RECT 441.200 8.800 442.000 9.000 ;
        RECT 445.800 8.800 446.600 9.000 ;
        RECT 447.200 9.000 447.800 10.200 ;
        RECT 449.200 10.400 449.800 11.600 ;
        RECT 452.200 11.400 453.000 11.600 ;
        RECT 455.600 11.400 456.400 11.700 ;
        RECT 457.200 11.600 458.000 11.700 ;
        RECT 458.800 11.600 459.400 14.600 ;
        RECT 462.000 11.600 462.800 13.200 ;
        RECT 463.600 11.600 464.200 14.600 ;
        RECT 466.800 13.800 467.600 19.800 ;
        RECT 473.200 16.600 474.000 19.800 ;
        RECT 474.800 17.000 475.600 19.800 ;
        RECT 476.400 17.000 477.200 19.800 ;
        RECT 478.000 17.000 478.800 19.800 ;
        RECT 481.200 17.000 482.000 19.800 ;
        RECT 484.400 17.000 485.200 19.800 ;
        RECT 486.000 17.000 486.800 19.800 ;
        RECT 487.600 17.000 488.400 19.800 ;
        RECT 489.200 17.000 490.000 19.800 ;
        RECT 471.400 15.800 474.000 16.600 ;
        RECT 490.800 16.600 491.600 19.800 ;
        RECT 477.400 15.800 482.000 16.400 ;
        RECT 471.400 15.200 472.200 15.800 ;
        RECT 469.200 14.400 472.200 15.200 ;
        RECT 466.800 13.000 475.600 13.800 ;
        RECT 477.400 13.400 478.200 15.800 ;
        RECT 481.200 15.600 482.000 15.800 ;
        RECT 482.800 15.600 484.400 16.400 ;
        RECT 487.400 15.600 488.400 16.400 ;
        RECT 490.800 15.800 493.200 16.600 ;
        RECT 479.600 13.600 480.400 15.200 ;
        RECT 481.200 14.800 482.000 15.000 ;
        RECT 481.200 14.200 485.600 14.800 ;
        RECT 484.800 14.000 485.600 14.200 ;
        RECT 452.200 10.800 456.400 11.400 ;
        RECT 449.200 9.800 451.600 10.400 ;
        RECT 448.600 9.000 449.400 9.200 ;
        RECT 447.200 8.400 449.400 9.000 ;
        RECT 451.000 8.800 451.600 9.800 ;
        RECT 451.000 8.000 452.400 8.800 ;
        RECT 444.600 7.400 445.400 7.600 ;
        RECT 447.400 7.400 448.200 7.600 ;
        RECT 441.200 6.200 442.000 7.000 ;
        RECT 444.600 6.800 448.200 7.400 ;
        RECT 446.800 6.200 447.400 6.800 ;
        RECT 450.800 6.200 451.600 7.000 ;
        RECT 441.200 5.600 443.200 6.200 ;
        RECT 442.400 2.200 443.200 5.600 ;
        RECT 446.800 2.200 447.600 6.200 ;
        RECT 451.000 2.200 452.200 6.200 ;
        RECT 455.600 2.200 456.400 10.800 ;
        RECT 458.800 10.800 460.000 11.600 ;
        RECT 463.600 10.800 464.800 11.600 ;
        RECT 458.800 10.200 459.400 10.800 ;
        RECT 463.600 10.200 464.200 10.800 ;
        RECT 457.200 9.600 459.400 10.200 ;
        RECT 462.000 9.600 464.200 10.200 ;
        RECT 457.200 2.200 458.000 9.600 ;
        RECT 462.000 2.200 462.800 9.600 ;
        RECT 466.800 7.400 467.600 13.000 ;
        RECT 476.200 12.600 478.200 13.400 ;
        RECT 482.000 12.600 485.200 13.400 ;
        RECT 487.600 12.800 488.400 15.600 ;
        RECT 492.400 15.200 493.200 15.800 ;
        RECT 492.400 14.600 494.200 15.200 ;
        RECT 493.400 13.400 494.200 14.600 ;
        RECT 497.200 14.600 498.000 19.800 ;
        RECT 498.800 16.000 499.600 19.800 ;
        RECT 498.800 15.200 499.800 16.000 ;
        RECT 502.000 15.600 502.800 17.200 ;
        RECT 497.200 14.000 498.400 14.600 ;
        RECT 493.400 12.600 497.200 13.400 ;
        RECT 468.200 12.000 469.000 12.200 ;
        RECT 473.200 12.000 474.000 12.400 ;
        RECT 490.800 12.000 491.600 12.600 ;
        RECT 497.800 12.000 498.400 14.000 ;
        RECT 468.200 11.400 491.600 12.000 ;
        RECT 497.600 11.400 498.400 12.000 ;
        RECT 497.600 9.600 498.200 11.400 ;
        RECT 499.000 10.800 499.800 15.200 ;
        RECT 476.400 9.400 477.200 9.600 ;
        RECT 471.800 9.000 477.200 9.400 ;
        RECT 471.000 8.800 477.200 9.000 ;
        RECT 478.200 9.000 486.800 9.600 ;
        RECT 468.400 8.000 470.000 8.800 ;
        RECT 471.000 8.200 472.400 8.800 ;
        RECT 478.200 8.200 478.800 9.000 ;
        RECT 486.000 8.800 486.800 9.000 ;
        RECT 489.200 9.000 498.200 9.600 ;
        RECT 489.200 8.800 490.000 9.000 ;
        RECT 469.400 7.600 470.000 8.000 ;
        RECT 473.000 7.600 478.800 8.200 ;
        RECT 479.400 7.600 482.000 8.400 ;
        RECT 466.800 6.800 468.800 7.400 ;
        RECT 469.400 6.800 473.600 7.600 ;
        RECT 468.200 6.200 468.800 6.800 ;
        RECT 468.200 5.600 469.200 6.200 ;
        RECT 468.400 2.200 469.200 5.600 ;
        RECT 471.600 2.200 472.400 6.800 ;
        RECT 474.800 2.200 475.600 5.000 ;
        RECT 476.400 2.200 477.200 5.000 ;
        RECT 478.000 2.200 478.800 7.000 ;
        RECT 481.200 2.200 482.000 7.000 ;
        RECT 484.400 2.200 485.200 8.400 ;
        RECT 492.400 7.600 495.000 8.400 ;
        RECT 487.600 6.800 491.800 7.600 ;
        RECT 486.000 2.200 486.800 5.000 ;
        RECT 487.600 2.200 488.400 5.000 ;
        RECT 489.200 2.200 490.000 5.000 ;
        RECT 492.400 2.200 493.200 7.600 ;
        RECT 497.600 7.400 498.200 9.000 ;
        RECT 495.600 6.800 498.200 7.400 ;
        RECT 498.800 10.000 499.800 10.800 ;
        RECT 495.600 2.200 496.400 6.800 ;
        RECT 498.800 2.200 499.600 10.000 ;
        RECT 503.600 2.200 504.400 19.800 ;
        RECT 505.200 13.800 506.000 19.800 ;
        RECT 511.600 16.600 512.400 19.800 ;
        RECT 513.200 17.000 514.000 19.800 ;
        RECT 514.800 17.000 515.600 19.800 ;
        RECT 516.400 17.000 517.200 19.800 ;
        RECT 519.600 17.000 520.400 19.800 ;
        RECT 522.800 17.000 523.600 19.800 ;
        RECT 524.400 17.000 525.200 19.800 ;
        RECT 526.000 17.000 526.800 19.800 ;
        RECT 527.600 17.000 528.400 19.800 ;
        RECT 509.800 15.800 512.400 16.600 ;
        RECT 529.200 16.600 530.000 19.800 ;
        RECT 515.800 15.800 520.400 16.400 ;
        RECT 509.800 15.200 510.600 15.800 ;
        RECT 507.600 14.400 510.600 15.200 ;
        RECT 505.200 13.000 514.000 13.800 ;
        RECT 515.800 13.400 516.600 15.800 ;
        RECT 519.600 15.600 520.400 15.800 ;
        RECT 521.200 15.600 522.800 16.400 ;
        RECT 525.800 15.600 526.800 16.400 ;
        RECT 529.200 15.800 531.600 16.600 ;
        RECT 518.000 13.600 518.800 15.200 ;
        RECT 519.600 14.800 520.400 15.000 ;
        RECT 519.600 14.200 524.000 14.800 ;
        RECT 523.200 14.000 524.000 14.200 ;
        RECT 505.200 7.400 506.000 13.000 ;
        RECT 514.600 12.600 516.600 13.400 ;
        RECT 520.400 12.600 523.600 13.400 ;
        RECT 526.000 12.800 526.800 15.600 ;
        RECT 530.800 15.200 531.600 15.800 ;
        RECT 530.800 14.600 532.600 15.200 ;
        RECT 531.800 13.400 532.600 14.600 ;
        RECT 535.600 14.600 536.400 19.800 ;
        RECT 537.200 16.000 538.000 19.800 ;
        RECT 537.200 15.200 538.200 16.000 ;
        RECT 535.600 14.000 536.800 14.600 ;
        RECT 531.800 12.600 535.600 13.400 ;
        RECT 506.600 12.000 507.400 12.200 ;
        RECT 510.000 12.000 510.800 12.400 ;
        RECT 511.600 12.000 512.400 12.400 ;
        RECT 529.200 12.000 530.000 12.600 ;
        RECT 536.200 12.000 536.800 14.000 ;
        RECT 506.600 11.400 530.000 12.000 ;
        RECT 536.000 11.400 536.800 12.000 ;
        RECT 537.400 12.300 538.200 15.200 ;
        RECT 540.400 15.200 541.200 19.800 ;
        RECT 545.200 15.200 546.000 19.800 ;
        RECT 540.400 14.600 542.600 15.200 ;
        RECT 545.200 14.600 547.400 15.200 ;
        RECT 540.400 12.300 541.200 13.200 ;
        RECT 537.400 11.700 541.200 12.300 ;
        RECT 536.000 9.600 536.600 11.400 ;
        RECT 537.400 10.800 538.200 11.700 ;
        RECT 540.400 11.600 541.200 11.700 ;
        RECT 542.000 11.600 542.600 14.600 ;
        RECT 545.200 11.600 546.000 13.200 ;
        RECT 546.800 11.600 547.400 14.600 ;
        RECT 514.800 9.400 515.600 9.600 ;
        RECT 510.200 9.000 515.600 9.400 ;
        RECT 509.400 8.800 515.600 9.000 ;
        RECT 516.600 9.000 525.200 9.600 ;
        RECT 506.800 8.000 508.400 8.800 ;
        RECT 509.400 8.200 510.800 8.800 ;
        RECT 516.600 8.200 517.200 9.000 ;
        RECT 524.400 8.800 525.200 9.000 ;
        RECT 527.600 9.000 536.600 9.600 ;
        RECT 527.600 8.800 528.400 9.000 ;
        RECT 507.800 7.600 508.400 8.000 ;
        RECT 511.400 7.600 517.200 8.200 ;
        RECT 517.800 7.600 520.400 8.400 ;
        RECT 505.200 6.800 507.200 7.400 ;
        RECT 507.800 6.800 512.000 7.600 ;
        RECT 506.600 6.200 507.200 6.800 ;
        RECT 506.600 5.600 507.600 6.200 ;
        RECT 506.800 2.200 507.600 5.600 ;
        RECT 510.000 2.200 510.800 6.800 ;
        RECT 513.200 2.200 514.000 5.000 ;
        RECT 514.800 2.200 515.600 5.000 ;
        RECT 516.400 2.200 517.200 7.000 ;
        RECT 519.600 2.200 520.400 7.000 ;
        RECT 522.800 2.200 523.600 8.400 ;
        RECT 530.800 7.600 533.400 8.400 ;
        RECT 526.000 6.800 530.200 7.600 ;
        RECT 524.400 2.200 525.200 5.000 ;
        RECT 526.000 2.200 526.800 5.000 ;
        RECT 527.600 2.200 528.400 5.000 ;
        RECT 530.800 2.200 531.600 7.600 ;
        RECT 536.000 7.400 536.600 9.000 ;
        RECT 534.000 6.800 536.600 7.400 ;
        RECT 537.200 10.000 538.200 10.800 ;
        RECT 542.000 10.800 543.200 11.600 ;
        RECT 546.800 10.800 548.000 11.600 ;
        RECT 542.000 10.200 542.600 10.800 ;
        RECT 546.800 10.200 547.400 10.800 ;
        RECT 534.000 2.200 534.800 6.800 ;
        RECT 537.200 2.200 538.000 10.000 ;
        RECT 540.400 9.600 542.600 10.200 ;
        RECT 545.200 9.600 547.400 10.200 ;
        RECT 540.400 2.200 541.200 9.600 ;
        RECT 545.200 2.200 546.000 9.600 ;
      LAYER via1 ;
        RECT 18.800 375.600 19.600 376.400 ;
        RECT 20.400 374.200 21.200 375.000 ;
        RECT 28.400 371.600 29.200 372.400 ;
        RECT 31.600 371.600 32.400 372.400 ;
        RECT 14.000 366.800 14.800 367.600 ;
        RECT 17.200 366.200 18.000 367.000 ;
        RECT 12.400 364.200 13.200 365.000 ;
        RECT 14.000 364.200 14.800 365.000 ;
        RECT 15.600 364.200 16.400 365.000 ;
        RECT 20.400 366.200 21.200 367.000 ;
        RECT 23.600 366.200 24.400 367.000 ;
        RECT 44.400 373.000 45.200 373.800 ;
        RECT 54.000 372.600 54.800 373.400 ;
        RECT 38.000 371.600 38.800 372.400 ;
        RECT 60.400 371.600 61.200 372.400 ;
        RECT 46.000 368.800 46.800 369.600 ;
        RECT 50.800 367.600 51.600 368.400 ;
        RECT 25.200 364.200 26.000 365.000 ;
        RECT 26.800 364.200 27.600 365.000 ;
        RECT 47.600 366.200 48.400 367.000 ;
        RECT 44.400 364.200 45.200 365.000 ;
        RECT 46.000 364.200 46.800 365.000 ;
        RECT 50.800 366.200 51.600 367.000 ;
        RECT 54.000 366.200 54.800 367.000 ;
        RECT 55.600 364.200 56.400 365.000 ;
        RECT 57.200 364.200 58.000 365.000 ;
        RECT 58.800 364.200 59.600 365.000 ;
        RECT 89.200 375.600 90.000 376.400 ;
        RECT 90.800 374.200 91.600 375.000 ;
        RECT 100.400 371.600 101.200 372.400 ;
        RECT 68.400 363.600 69.200 364.400 ;
        RECT 73.200 367.600 74.000 368.400 ;
        RECT 84.400 366.800 85.200 367.600 ;
        RECT 87.600 366.200 88.400 367.000 ;
        RECT 82.800 364.200 83.600 365.000 ;
        RECT 84.400 364.200 85.200 365.000 ;
        RECT 86.000 364.200 86.800 365.000 ;
        RECT 90.800 366.200 91.600 367.000 ;
        RECT 94.000 366.200 94.800 367.000 ;
        RECT 130.800 375.600 131.600 376.400 ;
        RECT 132.400 374.200 133.200 375.000 ;
        RECT 140.400 371.600 141.200 372.400 ;
        RECT 95.600 364.200 96.400 365.000 ;
        RECT 97.200 364.200 98.000 365.000 ;
        RECT 114.800 365.600 115.600 366.400 ;
        RECT 126.000 366.800 126.800 367.600 ;
        RECT 129.200 366.200 130.000 367.000 ;
        RECT 124.400 364.200 125.200 365.000 ;
        RECT 126.000 364.200 126.800 365.000 ;
        RECT 127.600 364.200 128.400 365.000 ;
        RECT 132.400 366.200 133.200 367.000 ;
        RECT 135.600 366.200 136.400 367.000 ;
        RECT 156.400 373.000 157.200 373.800 ;
        RECT 166.000 372.600 166.800 373.400 ;
        RECT 153.200 371.600 154.000 372.400 ;
        RECT 172.400 371.600 173.200 372.400 ;
        RECT 158.000 368.800 158.800 369.600 ;
        RECT 162.800 367.600 163.600 368.400 ;
        RECT 137.200 364.200 138.000 365.000 ;
        RECT 138.800 364.200 139.600 365.000 ;
        RECT 159.600 366.200 160.400 367.000 ;
        RECT 156.400 364.200 157.200 365.000 ;
        RECT 158.000 364.200 158.800 365.000 ;
        RECT 162.800 366.200 163.600 367.000 ;
        RECT 166.000 366.200 166.800 367.000 ;
        RECT 167.600 364.200 168.400 365.000 ;
        RECT 169.200 364.200 170.000 365.000 ;
        RECT 170.800 364.200 171.600 365.000 ;
        RECT 191.600 373.000 192.400 373.800 ;
        RECT 201.200 372.600 202.000 373.400 ;
        RECT 186.800 371.600 187.600 372.400 ;
        RECT 193.200 368.800 194.000 369.600 ;
        RECT 198.000 367.600 198.800 368.400 ;
        RECT 194.800 366.200 195.600 367.000 ;
        RECT 191.600 364.200 192.400 365.000 ;
        RECT 193.200 364.200 194.000 365.000 ;
        RECT 198.000 366.200 198.800 367.000 ;
        RECT 201.200 366.200 202.000 367.000 ;
        RECT 202.800 364.200 203.600 365.000 ;
        RECT 204.400 364.200 205.200 365.000 ;
        RECT 206.000 364.200 206.800 365.000 ;
        RECT 215.600 369.600 216.400 370.400 ;
        RECT 218.800 369.600 219.600 370.400 ;
        RECT 236.400 369.600 237.200 370.400 ;
        RECT 233.200 367.600 234.000 368.400 ;
        RECT 249.200 375.600 250.000 376.400 ;
        RECT 242.800 373.600 243.600 374.400 ;
        RECT 270.000 375.600 270.800 376.400 ;
        RECT 271.600 374.200 272.400 375.000 ;
        RECT 302.000 375.600 302.800 376.400 ;
        RECT 295.600 373.600 296.400 374.400 ;
        RECT 281.200 371.600 282.000 372.400 ;
        RECT 250.800 369.600 251.600 370.400 ;
        RECT 254.000 363.600 254.800 364.400 ;
        RECT 265.200 366.800 266.000 367.600 ;
        RECT 268.400 366.200 269.200 367.000 ;
        RECT 263.600 364.200 264.400 365.000 ;
        RECT 265.200 364.200 266.000 365.000 ;
        RECT 266.800 364.200 267.600 365.000 ;
        RECT 271.600 366.200 272.400 367.000 ;
        RECT 274.800 366.200 275.600 367.000 ;
        RECT 276.400 364.200 277.200 365.000 ;
        RECT 278.000 364.200 278.800 365.000 ;
        RECT 303.600 369.600 304.400 370.400 ;
        RECT 318.000 371.600 318.800 372.400 ;
        RECT 322.800 371.600 323.600 372.400 ;
        RECT 305.200 363.600 306.000 364.400 ;
        RECT 332.400 369.600 333.200 370.400 ;
        RECT 334.000 369.600 334.800 370.400 ;
        RECT 327.600 365.600 328.400 366.400 ;
        RECT 337.200 369.600 338.000 370.400 ;
        RECT 346.800 373.600 347.600 374.400 ;
        RECT 356.400 373.000 357.200 373.800 ;
        RECT 366.000 372.600 366.800 373.400 ;
        RECT 388.400 377.600 389.200 378.400 ;
        RECT 358.000 368.800 358.800 369.600 ;
        RECT 362.800 367.600 363.600 368.400 ;
        RECT 359.600 366.200 360.400 367.000 ;
        RECT 356.400 364.200 357.200 365.000 ;
        RECT 358.000 364.200 358.800 365.000 ;
        RECT 362.800 366.200 363.600 367.000 ;
        RECT 366.000 366.200 366.800 367.000 ;
        RECT 367.600 364.200 368.400 365.000 ;
        RECT 369.200 364.200 370.000 365.000 ;
        RECT 370.800 364.200 371.600 365.000 ;
        RECT 386.800 371.600 387.600 372.400 ;
        RECT 402.800 373.000 403.600 373.800 ;
        RECT 380.400 363.600 381.200 364.400 ;
        RECT 412.400 372.600 413.200 373.400 ;
        RECT 399.600 371.600 400.400 372.400 ;
        RECT 427.000 373.600 427.800 374.400 ;
        RECT 404.400 368.800 405.200 369.600 ;
        RECT 409.200 367.600 410.000 368.400 ;
        RECT 406.000 366.200 406.800 367.000 ;
        RECT 402.800 364.200 403.600 365.000 ;
        RECT 404.400 364.200 405.200 365.000 ;
        RECT 409.200 366.200 410.000 367.000 ;
        RECT 412.400 366.200 413.200 367.000 ;
        RECT 414.000 364.200 414.800 365.000 ;
        RECT 415.600 364.200 416.400 365.000 ;
        RECT 417.200 364.200 418.000 365.000 ;
        RECT 437.800 371.600 438.600 372.400 ;
        RECT 454.000 375.600 454.800 376.400 ;
        RECT 455.600 374.200 456.400 375.000 ;
        RECT 463.600 371.600 464.400 372.400 ;
        RECT 449.200 366.800 450.000 367.600 ;
        RECT 452.400 366.200 453.200 367.000 ;
        RECT 447.600 364.200 448.400 365.000 ;
        RECT 449.200 364.200 450.000 365.000 ;
        RECT 450.800 364.200 451.600 365.000 ;
        RECT 455.600 366.200 456.400 367.000 ;
        RECT 458.800 366.200 459.600 367.000 ;
        RECT 479.600 373.000 480.400 373.800 ;
        RECT 489.200 372.600 490.000 373.400 ;
        RECT 474.800 371.600 475.600 372.400 ;
        RECT 495.600 371.600 496.400 372.400 ;
        RECT 481.200 368.800 482.000 369.600 ;
        RECT 486.000 367.600 486.800 368.400 ;
        RECT 460.400 364.200 461.200 365.000 ;
        RECT 462.000 364.200 462.800 365.000 ;
        RECT 482.800 366.200 483.600 367.000 ;
        RECT 479.600 364.200 480.400 365.000 ;
        RECT 481.200 364.200 482.000 365.000 ;
        RECT 486.000 366.200 486.800 367.000 ;
        RECT 489.200 366.200 490.000 367.000 ;
        RECT 490.800 364.200 491.600 365.000 ;
        RECT 492.400 364.200 493.200 365.000 ;
        RECT 494.000 364.200 494.800 365.000 ;
        RECT 529.200 375.600 530.000 376.400 ;
        RECT 530.800 374.200 531.600 375.000 ;
        RECT 521.200 371.600 522.000 372.400 ;
        RECT 542.000 371.600 542.800 372.400 ;
        RECT 510.000 369.600 510.800 370.400 ;
        RECT 503.600 363.600 504.400 364.400 ;
        RECT 513.200 363.600 514.000 364.400 ;
        RECT 524.400 366.800 525.200 367.600 ;
        RECT 527.600 366.200 528.400 367.000 ;
        RECT 522.800 364.200 523.600 365.000 ;
        RECT 524.400 364.200 525.200 365.000 ;
        RECT 526.000 364.200 526.800 365.000 ;
        RECT 530.800 366.200 531.600 367.000 ;
        RECT 534.000 366.200 534.800 367.000 ;
        RECT 535.600 364.200 536.400 365.000 ;
        RECT 537.200 364.200 538.000 365.000 ;
        RECT 546.800 363.600 547.600 364.400 ;
        RECT 14.000 354.400 14.800 355.200 ;
        RECT 17.200 355.000 18.000 355.800 ;
        RECT 12.400 352.400 13.200 353.200 ;
        RECT 2.800 343.600 3.600 344.400 ;
        RECT 22.000 347.600 22.800 348.400 ;
        RECT 18.800 345.600 19.600 346.400 ;
        RECT 12.400 344.200 13.200 345.000 ;
        RECT 14.000 344.200 14.800 345.000 ;
        RECT 15.600 344.200 16.400 345.000 ;
        RECT 17.200 344.200 18.000 345.000 ;
        RECT 20.400 344.200 21.200 345.000 ;
        RECT 23.600 344.200 24.400 345.000 ;
        RECT 25.200 344.200 26.000 345.000 ;
        RECT 26.800 344.200 27.600 345.000 ;
        RECT 38.000 345.600 38.800 346.400 ;
        RECT 42.800 345.600 43.600 346.400 ;
        RECT 47.600 345.600 48.400 346.400 ;
        RECT 49.200 345.600 50.000 346.400 ;
        RECT 54.000 347.600 54.800 348.400 ;
        RECT 41.200 343.600 42.000 344.400 ;
        RECT 46.000 343.600 46.800 344.400 ;
        RECT 76.400 355.000 77.200 355.800 ;
        RECT 73.200 353.600 74.000 354.400 ;
        RECT 78.000 352.400 78.800 353.200 ;
        RECT 82.800 349.600 83.600 350.400 ;
        RECT 66.800 348.200 67.600 349.000 ;
        RECT 76.400 348.600 77.200 349.400 ;
        RECT 71.600 347.600 72.400 348.400 ;
        RECT 66.800 344.200 67.600 345.000 ;
        RECT 68.400 344.200 69.200 345.000 ;
        RECT 70.000 344.200 70.800 345.000 ;
        RECT 73.200 344.200 74.000 345.000 ;
        RECT 76.400 344.200 77.200 345.000 ;
        RECT 78.000 344.200 78.800 345.000 ;
        RECT 79.600 344.200 80.400 345.000 ;
        RECT 81.200 344.200 82.000 345.000 ;
        RECT 116.400 355.000 117.200 355.800 ;
        RECT 113.200 353.600 114.000 354.400 ;
        RECT 118.000 352.400 118.800 353.200 ;
        RECT 122.800 349.600 123.600 350.400 ;
        RECT 106.800 348.200 107.600 349.000 ;
        RECT 116.400 348.600 117.200 349.400 ;
        RECT 97.200 345.600 98.000 346.400 ;
        RECT 95.600 343.600 96.400 344.400 ;
        RECT 111.600 347.600 112.400 348.400 ;
        RECT 106.800 344.200 107.600 345.000 ;
        RECT 108.400 344.200 109.200 345.000 ;
        RECT 110.000 344.200 110.800 345.000 ;
        RECT 113.200 344.200 114.000 345.000 ;
        RECT 116.400 344.200 117.200 345.000 ;
        RECT 118.000 344.200 118.800 345.000 ;
        RECT 119.600 344.200 120.400 345.000 ;
        RECT 121.200 344.200 122.000 345.000 ;
        RECT 158.000 355.000 158.800 355.800 ;
        RECT 154.800 353.600 155.600 354.400 ;
        RECT 159.600 352.400 160.400 353.200 ;
        RECT 148.400 348.200 149.200 349.000 ;
        RECT 158.000 348.600 158.800 349.400 ;
        RECT 130.800 343.600 131.600 344.400 ;
        RECT 153.200 347.600 154.000 348.400 ;
        RECT 148.400 344.200 149.200 345.000 ;
        RECT 150.000 344.200 150.800 345.000 ;
        RECT 151.600 344.200 152.400 345.000 ;
        RECT 154.800 344.200 155.600 345.000 ;
        RECT 158.000 344.200 158.800 345.000 ;
        RECT 159.600 344.200 160.400 345.000 ;
        RECT 161.200 344.200 162.000 345.000 ;
        RECT 162.800 344.200 163.600 345.000 ;
        RECT 188.400 354.400 189.200 355.200 ;
        RECT 191.600 355.000 192.400 355.800 ;
        RECT 186.800 352.400 187.600 353.200 ;
        RECT 172.400 343.600 173.200 344.400 ;
        RECT 177.200 343.600 178.000 344.400 ;
        RECT 196.400 347.600 197.200 348.400 ;
        RECT 193.200 345.600 194.000 346.400 ;
        RECT 186.800 344.200 187.600 345.000 ;
        RECT 188.400 344.200 189.200 345.000 ;
        RECT 190.000 344.200 190.800 345.000 ;
        RECT 191.600 344.200 192.400 345.000 ;
        RECT 194.800 344.200 195.600 345.000 ;
        RECT 198.000 344.200 198.800 345.000 ;
        RECT 199.600 344.200 200.400 345.000 ;
        RECT 201.200 344.200 202.000 345.000 ;
        RECT 223.600 354.400 224.400 355.200 ;
        RECT 226.800 355.000 227.600 355.800 ;
        RECT 246.000 357.600 246.800 358.400 ;
        RECT 252.400 357.600 253.200 358.400 ;
        RECT 222.000 352.400 222.800 353.200 ;
        RECT 220.400 349.600 221.200 350.400 ;
        RECT 212.400 343.600 213.200 344.400 ;
        RECT 247.600 353.600 248.400 354.400 ;
        RECT 254.000 353.600 254.800 354.400 ;
        RECT 231.600 347.600 232.400 348.400 ;
        RECT 228.400 345.600 229.200 346.400 ;
        RECT 222.000 344.200 222.800 345.000 ;
        RECT 223.600 344.200 224.400 345.000 ;
        RECT 225.200 344.200 226.000 345.000 ;
        RECT 226.800 344.200 227.600 345.000 ;
        RECT 230.000 344.200 230.800 345.000 ;
        RECT 233.200 344.200 234.000 345.000 ;
        RECT 234.800 344.200 235.600 345.000 ;
        RECT 236.400 344.200 237.200 345.000 ;
        RECT 250.800 351.600 251.600 352.400 ;
        RECT 249.200 349.600 250.000 350.400 ;
        RECT 257.200 351.600 258.000 352.400 ;
        RECT 255.600 349.600 256.400 350.400 ;
        RECT 282.800 355.000 283.600 355.800 ;
        RECT 279.600 353.600 280.400 354.400 ;
        RECT 284.400 352.400 285.200 353.200 ;
        RECT 303.600 357.600 304.400 358.400 ;
        RECT 302.000 353.600 302.800 354.400 ;
        RECT 311.600 357.600 312.400 358.400 ;
        RECT 273.200 348.200 274.000 349.000 ;
        RECT 282.800 348.600 283.600 349.400 ;
        RECT 278.000 347.600 278.800 348.400 ;
        RECT 297.400 349.600 298.200 350.400 ;
        RECT 273.200 344.200 274.000 345.000 ;
        RECT 274.800 344.200 275.600 345.000 ;
        RECT 276.400 344.200 277.200 345.000 ;
        RECT 279.600 344.200 280.400 345.000 ;
        RECT 282.800 344.200 283.600 345.000 ;
        RECT 284.400 344.200 285.200 345.000 ;
        RECT 286.000 344.200 286.800 345.000 ;
        RECT 287.600 344.200 288.400 345.000 ;
        RECT 305.200 351.600 306.000 352.400 ;
        RECT 319.600 357.600 320.400 358.400 ;
        RECT 303.600 349.600 304.400 350.400 ;
        RECT 310.000 345.600 310.800 346.400 ;
        RECT 318.000 347.600 318.800 348.400 ;
        RECT 326.000 357.600 326.800 358.400 ;
        RECT 324.400 353.600 325.200 354.400 ;
        RECT 327.600 351.600 328.400 352.400 ;
        RECT 337.200 353.600 338.000 354.400 ;
        RECT 326.000 349.600 326.800 350.400 ;
        RECT 340.400 351.600 341.200 352.400 ;
        RECT 361.200 357.600 362.000 358.400 ;
        RECT 369.200 357.600 370.000 358.400 ;
        RECT 338.800 349.600 339.600 350.400 ;
        RECT 353.200 349.600 354.000 350.400 ;
        RECT 378.800 355.600 379.600 356.400 ;
        RECT 375.600 353.600 376.400 354.400 ;
        RECT 361.200 349.600 362.000 350.400 ;
        RECT 366.000 349.600 366.800 350.400 ;
        RECT 369.200 349.600 370.000 350.400 ;
        RECT 375.600 349.600 376.400 350.400 ;
        RECT 337.200 347.600 338.000 348.400 ;
        RECT 345.200 345.600 346.000 346.400 ;
        RECT 362.800 347.600 363.600 348.400 ;
        RECT 377.200 347.600 378.000 348.400 ;
        RECT 388.400 357.600 389.200 358.400 ;
        RECT 406.000 357.600 406.800 358.400 ;
        RECT 386.800 347.600 387.600 348.400 ;
        RECT 385.200 345.600 386.000 346.400 ;
        RECT 423.600 345.600 424.400 346.400 ;
        RECT 436.400 347.600 437.200 348.400 ;
        RECT 446.000 357.600 446.800 358.400 ;
        RECT 444.400 353.600 445.200 354.400 ;
        RECT 457.200 357.600 458.000 358.400 ;
        RECT 441.200 351.600 442.000 352.400 ;
        RECT 449.200 349.600 450.000 350.400 ;
        RECT 455.600 349.600 456.400 350.400 ;
        RECT 465.200 351.600 466.000 352.400 ;
        RECT 458.800 349.600 459.600 350.400 ;
        RECT 465.200 349.600 466.000 350.400 ;
        RECT 439.600 343.600 440.400 344.400 ;
        RECT 466.800 347.600 467.600 348.400 ;
        RECT 473.200 349.600 474.000 350.400 ;
        RECT 479.600 349.600 480.400 350.400 ;
        RECT 468.400 345.600 469.200 346.400 ;
        RECT 470.000 345.600 470.800 346.400 ;
        RECT 484.400 345.600 485.200 346.400 ;
        RECT 505.200 357.600 506.000 358.400 ;
        RECT 508.400 357.600 509.200 358.400 ;
        RECT 494.000 353.600 494.800 354.400 ;
        RECT 500.400 353.600 501.200 354.400 ;
        RECT 487.600 345.600 488.400 346.400 ;
        RECT 486.000 343.600 486.800 344.400 ;
        RECT 497.200 351.600 498.000 352.400 ;
        RECT 527.600 354.400 528.400 355.200 ;
        RECT 530.800 355.000 531.600 355.800 ;
        RECT 526.000 352.400 526.800 353.200 ;
        RECT 506.800 345.600 507.600 346.400 ;
        RECT 516.400 343.600 517.200 344.400 ;
        RECT 535.600 347.600 536.400 348.400 ;
        RECT 532.400 345.600 533.200 346.400 ;
        RECT 526.000 344.200 526.800 345.000 ;
        RECT 527.600 344.200 528.400 345.000 ;
        RECT 529.200 344.200 530.000 345.000 ;
        RECT 530.800 344.200 531.600 345.000 ;
        RECT 534.000 344.200 534.800 345.000 ;
        RECT 537.200 344.200 538.000 345.000 ;
        RECT 538.800 344.200 539.600 345.000 ;
        RECT 540.400 344.200 541.200 345.000 ;
        RECT 22.000 335.600 22.800 336.400 ;
        RECT 23.600 334.200 24.400 335.000 ;
        RECT 44.400 337.600 45.200 338.400 ;
        RECT 31.600 331.600 32.400 332.400 ;
        RECT 2.800 323.600 3.600 324.400 ;
        RECT 17.200 326.800 18.000 327.600 ;
        RECT 20.400 326.200 21.200 327.000 ;
        RECT 15.600 324.200 16.400 325.000 ;
        RECT 17.200 324.200 18.000 325.000 ;
        RECT 18.800 324.200 19.600 325.000 ;
        RECT 23.600 326.200 24.400 327.000 ;
        RECT 26.800 326.200 27.600 327.000 ;
        RECT 28.400 324.200 29.200 325.000 ;
        RECT 30.000 324.200 30.800 325.000 ;
        RECT 42.800 329.600 43.600 330.400 ;
        RECT 52.400 325.600 53.200 326.400 ;
        RECT 70.000 329.600 70.800 330.400 ;
        RECT 74.800 329.600 75.600 330.400 ;
        RECT 82.800 331.600 83.600 332.400 ;
        RECT 87.600 331.600 88.400 332.400 ;
        RECT 90.800 331.600 91.600 332.400 ;
        RECT 87.600 323.600 88.400 324.400 ;
        RECT 111.600 335.600 112.400 336.400 ;
        RECT 113.200 334.200 114.000 335.000 ;
        RECT 122.800 331.600 123.600 332.400 ;
        RECT 95.600 323.600 96.400 324.400 ;
        RECT 106.800 326.800 107.600 327.600 ;
        RECT 110.000 326.200 110.800 327.000 ;
        RECT 105.200 324.200 106.000 325.000 ;
        RECT 106.800 324.200 107.600 325.000 ;
        RECT 108.400 324.200 109.200 325.000 ;
        RECT 113.200 326.200 114.000 327.000 ;
        RECT 116.400 326.200 117.200 327.000 ;
        RECT 143.600 333.000 144.400 333.800 ;
        RECT 153.200 332.600 154.000 333.400 ;
        RECT 140.400 331.600 141.200 332.400 ;
        RECT 159.600 331.600 160.400 332.400 ;
        RECT 175.600 337.600 176.400 338.400 ;
        RECT 145.200 328.800 146.000 329.600 ;
        RECT 150.000 327.600 150.800 328.400 ;
        RECT 118.000 324.200 118.800 325.000 ;
        RECT 119.600 324.200 120.400 325.000 ;
        RECT 146.800 326.200 147.600 327.000 ;
        RECT 143.600 324.200 144.400 325.000 ;
        RECT 145.200 324.200 146.000 325.000 ;
        RECT 150.000 326.200 150.800 327.000 ;
        RECT 153.200 326.200 154.000 327.000 ;
        RECT 154.800 324.200 155.600 325.000 ;
        RECT 156.400 324.200 157.200 325.000 ;
        RECT 158.000 324.200 158.800 325.000 ;
        RECT 199.600 337.600 200.400 338.400 ;
        RECT 167.600 323.600 168.400 324.400 ;
        RECT 193.200 333.600 194.000 334.400 ;
        RECT 186.800 323.600 187.600 324.400 ;
        RECT 199.600 329.600 200.400 330.400 ;
        RECT 209.200 337.600 210.000 338.400 ;
        RECT 204.400 329.600 205.200 330.400 ;
        RECT 202.800 323.600 203.600 324.400 ;
        RECT 236.400 335.600 237.200 336.400 ;
        RECT 238.000 334.200 238.800 335.000 ;
        RECT 265.200 337.600 266.000 338.400 ;
        RECT 228.400 331.600 229.200 332.400 ;
        RECT 210.800 323.600 211.600 324.400 ;
        RECT 220.400 323.600 221.200 324.400 ;
        RECT 231.600 326.800 232.400 327.600 ;
        RECT 234.800 326.200 235.600 327.000 ;
        RECT 230.000 324.200 230.800 325.000 ;
        RECT 231.600 324.200 232.400 325.000 ;
        RECT 233.200 324.200 234.000 325.000 ;
        RECT 238.000 326.200 238.800 327.000 ;
        RECT 241.200 326.200 242.000 327.000 ;
        RECT 282.800 333.000 283.600 333.800 ;
        RECT 242.800 324.200 243.600 325.000 ;
        RECT 244.400 324.200 245.200 325.000 ;
        RECT 292.400 332.600 293.200 333.400 ;
        RECT 281.200 331.600 282.000 332.400 ;
        RECT 284.400 328.800 285.200 329.600 ;
        RECT 289.200 327.600 290.000 328.400 ;
        RECT 286.000 326.200 286.800 327.000 ;
        RECT 282.800 324.200 283.600 325.000 ;
        RECT 284.400 324.200 285.200 325.000 ;
        RECT 289.200 326.200 290.000 327.000 ;
        RECT 292.400 326.200 293.200 327.000 ;
        RECT 294.000 324.200 294.800 325.000 ;
        RECT 295.600 324.200 296.400 325.000 ;
        RECT 297.200 324.200 298.000 325.000 ;
        RECT 318.000 333.000 318.800 333.800 ;
        RECT 327.600 332.600 328.400 333.400 ;
        RECT 311.600 331.600 312.400 332.400 ;
        RECT 314.800 331.600 315.600 332.400 ;
        RECT 319.600 328.800 320.400 329.600 ;
        RECT 324.400 327.600 325.200 328.400 ;
        RECT 306.800 323.600 307.600 324.400 ;
        RECT 321.200 326.200 322.000 327.000 ;
        RECT 318.000 324.200 318.800 325.000 ;
        RECT 319.600 324.200 320.400 325.000 ;
        RECT 324.400 326.200 325.200 327.000 ;
        RECT 327.600 326.200 328.400 327.000 ;
        RECT 329.200 324.200 330.000 325.000 ;
        RECT 330.800 324.200 331.600 325.000 ;
        RECT 332.400 324.200 333.200 325.000 ;
        RECT 351.600 337.600 352.400 338.400 ;
        RECT 346.800 323.600 347.600 324.400 ;
        RECT 354.800 333.600 355.600 334.400 ;
        RECT 351.600 329.600 352.400 330.400 ;
        RECT 369.200 323.600 370.000 324.400 ;
        RECT 375.600 329.600 376.400 330.400 ;
        RECT 383.600 329.600 384.400 330.400 ;
        RECT 388.400 337.600 389.200 338.400 ;
        RECT 386.800 323.600 387.600 324.400 ;
        RECT 394.800 329.600 395.600 330.400 ;
        RECT 401.200 325.600 402.000 326.400 ;
        RECT 407.600 325.600 408.400 326.400 ;
        RECT 450.800 337.600 451.600 338.400 ;
        RECT 439.600 323.600 440.400 324.400 ;
        RECT 466.800 333.000 467.600 333.800 ;
        RECT 476.400 332.600 477.200 333.400 ;
        RECT 463.600 331.600 464.400 332.400 ;
        RECT 465.200 331.600 466.000 332.400 ;
        RECT 468.400 328.800 469.200 329.600 ;
        RECT 473.200 327.600 474.000 328.400 ;
        RECT 470.000 326.200 470.800 327.000 ;
        RECT 466.800 324.200 467.600 325.000 ;
        RECT 468.400 324.200 469.200 325.000 ;
        RECT 473.200 326.200 474.000 327.000 ;
        RECT 476.400 326.200 477.200 327.000 ;
        RECT 478.000 324.200 478.800 325.000 ;
        RECT 479.600 324.200 480.400 325.000 ;
        RECT 481.200 324.200 482.000 325.000 ;
        RECT 494.000 329.600 494.800 330.400 ;
        RECT 490.800 323.600 491.600 324.400 ;
        RECT 534.000 337.600 534.800 338.400 ;
        RECT 518.000 331.600 518.800 332.400 ;
        RECT 521.200 331.600 522.000 332.400 ;
        RECT 505.200 323.600 506.000 324.400 ;
        RECT 513.200 329.600 514.000 330.400 ;
        RECT 519.600 329.600 520.400 330.400 ;
        RECT 534.000 329.600 534.800 330.400 ;
        RECT 540.400 327.600 541.200 328.400 ;
        RECT 9.200 313.600 10.000 314.400 ;
        RECT 12.400 313.600 13.200 314.400 ;
        RECT 6.000 311.600 6.800 312.400 ;
        RECT 4.400 305.600 5.200 306.400 ;
        RECT 10.800 303.600 11.600 304.400 ;
        RECT 30.000 317.600 30.800 318.400 ;
        RECT 17.200 313.600 18.000 314.400 ;
        RECT 23.600 313.600 24.400 314.400 ;
        RECT 18.800 309.600 19.600 310.400 ;
        RECT 14.000 305.600 14.800 306.400 ;
        RECT 22.000 307.600 22.800 308.400 ;
        RECT 41.200 313.600 42.000 314.400 ;
        RECT 52.400 315.600 53.200 316.400 ;
        RECT 57.200 317.600 58.000 318.400 ;
        RECT 30.000 309.600 30.800 310.400 ;
        RECT 44.400 309.600 45.200 310.400 ;
        RECT 47.600 309.600 48.400 310.400 ;
        RECT 31.600 307.600 32.400 308.400 ;
        RECT 33.200 305.600 34.000 306.400 ;
        RECT 38.000 305.600 38.800 306.400 ;
        RECT 50.800 307.600 51.600 308.400 ;
        RECT 63.600 317.600 64.400 318.400 ;
        RECT 55.600 311.600 56.400 312.400 ;
        RECT 62.000 307.600 62.800 308.400 ;
        RECT 71.600 309.600 72.400 310.400 ;
        RECT 74.800 305.600 75.600 306.400 ;
        RECT 76.400 305.600 77.200 306.400 ;
        RECT 105.200 313.600 106.000 314.400 ;
        RECT 102.000 307.600 102.800 308.400 ;
        RECT 103.600 307.600 104.400 308.400 ;
        RECT 110.000 311.600 110.800 312.400 ;
        RECT 108.400 305.600 109.200 306.400 ;
        RECT 111.600 305.600 112.400 306.400 ;
        RECT 134.000 313.600 134.800 314.400 ;
        RECT 137.200 311.600 138.000 312.400 ;
        RECT 135.600 309.600 136.400 310.400 ;
        RECT 140.400 309.600 141.200 310.400 ;
        RECT 156.400 317.600 157.200 318.400 ;
        RECT 169.200 309.600 170.000 310.400 ;
        RECT 175.600 309.600 176.400 310.400 ;
        RECT 170.800 307.600 171.600 308.400 ;
        RECT 178.800 305.600 179.600 306.400 ;
        RECT 194.800 317.600 195.600 318.400 ;
        RECT 194.800 309.600 195.600 310.400 ;
        RECT 186.800 305.600 187.600 306.400 ;
        RECT 196.400 307.600 197.200 308.400 ;
        RECT 199.600 305.600 200.400 306.400 ;
        RECT 209.200 309.600 210.000 310.400 ;
        RECT 214.000 309.600 214.800 310.400 ;
        RECT 210.800 307.600 211.600 308.400 ;
        RECT 226.800 307.600 227.600 308.400 ;
        RECT 236.400 309.600 237.200 310.400 ;
        RECT 238.000 307.600 238.800 308.400 ;
        RECT 244.400 309.600 245.200 310.400 ;
        RECT 262.000 314.400 262.800 315.200 ;
        RECT 265.200 315.000 266.000 315.800 ;
        RECT 260.400 312.400 261.200 313.200 ;
        RECT 217.200 303.600 218.000 304.400 ;
        RECT 250.800 303.600 251.600 304.400 ;
        RECT 270.000 307.600 270.800 308.400 ;
        RECT 266.800 305.600 267.600 306.400 ;
        RECT 260.400 304.200 261.200 305.000 ;
        RECT 262.000 304.200 262.800 305.000 ;
        RECT 263.600 304.200 264.400 305.000 ;
        RECT 265.200 304.200 266.000 305.000 ;
        RECT 268.400 304.200 269.200 305.000 ;
        RECT 271.600 304.200 272.400 305.000 ;
        RECT 273.200 304.200 274.000 305.000 ;
        RECT 274.800 304.200 275.600 305.000 ;
        RECT 303.600 314.400 304.400 315.200 ;
        RECT 306.800 315.000 307.600 315.800 ;
        RECT 302.000 312.400 302.800 313.200 ;
        RECT 318.000 311.200 318.800 312.000 ;
        RECT 292.400 303.600 293.200 304.400 ;
        RECT 330.800 317.600 331.600 318.400 ;
        RECT 335.600 313.600 336.400 314.400 ;
        RECT 311.600 307.600 312.400 308.400 ;
        RECT 308.400 305.600 309.200 306.400 ;
        RECT 302.000 304.200 302.800 305.000 ;
        RECT 303.600 304.200 304.400 305.000 ;
        RECT 305.200 304.200 306.000 305.000 ;
        RECT 306.800 304.200 307.600 305.000 ;
        RECT 310.000 304.200 310.800 305.000 ;
        RECT 313.200 304.200 314.000 305.000 ;
        RECT 314.800 304.200 315.600 305.000 ;
        RECT 316.400 304.200 317.200 305.000 ;
        RECT 335.600 309.600 336.400 310.400 ;
        RECT 337.200 307.600 338.000 308.400 ;
        RECT 345.200 309.600 346.000 310.400 ;
        RECT 348.400 309.600 349.200 310.400 ;
        RECT 359.600 317.600 360.400 318.400 ;
        RECT 361.200 313.600 362.000 314.400 ;
        RECT 358.000 311.600 358.800 312.400 ;
        RECT 340.400 305.600 341.200 306.400 ;
        RECT 356.400 307.600 357.200 308.400 ;
        RECT 369.200 317.600 370.000 318.400 ;
        RECT 364.400 305.600 365.200 306.400 ;
        RECT 378.800 307.600 379.600 308.400 ;
        RECT 399.600 317.600 400.400 318.400 ;
        RECT 401.200 313.600 402.000 314.400 ;
        RECT 407.600 317.600 408.400 318.400 ;
        RECT 406.000 313.600 406.800 314.400 ;
        RECT 398.000 311.600 398.800 312.400 ;
        RECT 394.800 309.600 395.600 310.400 ;
        RECT 390.000 305.600 390.800 306.400 ;
        RECT 396.400 307.600 397.200 308.400 ;
        RECT 409.200 311.600 410.000 312.400 ;
        RECT 407.600 309.600 408.400 310.400 ;
        RECT 433.200 309.600 434.000 310.400 ;
        RECT 417.200 305.600 418.000 306.400 ;
        RECT 428.400 305.600 429.200 306.400 ;
        RECT 458.800 315.000 459.600 315.800 ;
        RECT 455.600 313.600 456.400 314.400 ;
        RECT 473.200 317.600 474.000 318.400 ;
        RECT 460.400 312.400 461.200 313.200 ;
        RECT 478.000 317.600 478.800 318.400 ;
        RECT 465.200 309.600 466.000 310.400 ;
        RECT 449.200 308.200 450.000 309.000 ;
        RECT 458.800 308.600 459.600 309.400 ;
        RECT 439.600 305.600 440.400 306.400 ;
        RECT 454.000 307.600 454.800 308.400 ;
        RECT 449.200 304.200 450.000 305.000 ;
        RECT 450.800 304.200 451.600 305.000 ;
        RECT 452.400 304.200 453.200 305.000 ;
        RECT 455.600 304.200 456.400 305.000 ;
        RECT 458.800 304.200 459.600 305.000 ;
        RECT 460.400 304.200 461.200 305.000 ;
        RECT 462.000 304.200 462.800 305.000 ;
        RECT 463.600 304.200 464.400 305.000 ;
        RECT 495.600 317.600 496.400 318.400 ;
        RECT 481.200 303.600 482.000 304.400 ;
        RECT 494.000 305.600 494.800 306.400 ;
        RECT 498.800 317.600 499.600 318.400 ;
        RECT 503.600 309.600 504.400 310.400 ;
        RECT 511.600 309.600 512.400 310.400 ;
        RECT 524.400 317.600 525.200 318.400 ;
        RECT 506.800 305.600 507.600 306.400 ;
        RECT 516.400 305.600 517.200 306.400 ;
        RECT 514.800 303.600 515.600 304.400 ;
        RECT 530.800 309.600 531.600 310.400 ;
        RECT 537.200 309.600 538.000 310.400 ;
        RECT 526.000 305.600 526.800 306.400 ;
        RECT 534.000 303.600 534.800 304.400 ;
        RECT 543.600 303.600 544.400 304.400 ;
        RECT 4.400 291.600 5.200 292.400 ;
        RECT 14.000 291.600 14.800 292.400 ;
        RECT 4.400 283.600 5.200 284.400 ;
        RECT 20.400 295.600 21.200 296.400 ;
        RECT 28.400 289.600 29.200 290.400 ;
        RECT 23.600 283.600 24.400 284.400 ;
        RECT 39.600 297.600 40.400 298.400 ;
        RECT 36.400 291.600 37.200 292.400 ;
        RECT 55.600 295.600 56.400 296.400 ;
        RECT 57.200 294.200 58.000 295.000 ;
        RECT 47.600 291.600 48.400 292.400 ;
        RECT 68.400 291.600 69.200 292.400 ;
        RECT 36.400 283.600 37.200 284.400 ;
        RECT 39.600 283.600 40.400 284.400 ;
        RECT 50.800 286.800 51.600 287.600 ;
        RECT 54.000 286.200 54.800 287.000 ;
        RECT 49.200 284.200 50.000 285.000 ;
        RECT 50.800 284.200 51.600 285.000 ;
        RECT 52.400 284.200 53.200 285.000 ;
        RECT 57.200 286.200 58.000 287.000 ;
        RECT 60.400 286.200 61.200 287.000 ;
        RECT 90.800 295.600 91.600 296.400 ;
        RECT 92.400 294.200 93.200 295.000 ;
        RECT 82.800 291.600 83.600 292.400 ;
        RECT 103.600 291.600 104.400 292.400 ;
        RECT 62.000 284.200 62.800 285.000 ;
        RECT 63.600 284.200 64.400 285.000 ;
        RECT 74.800 283.600 75.600 284.400 ;
        RECT 86.000 286.800 86.800 287.600 ;
        RECT 89.200 286.200 90.000 287.000 ;
        RECT 84.400 284.200 85.200 285.000 ;
        RECT 86.000 284.200 86.800 285.000 ;
        RECT 87.600 284.200 88.400 285.000 ;
        RECT 92.400 286.200 93.200 287.000 ;
        RECT 95.600 286.200 96.400 287.000 ;
        RECT 108.400 289.600 109.200 290.400 ;
        RECT 97.200 284.200 98.000 285.000 ;
        RECT 98.800 284.200 99.600 285.000 ;
        RECT 122.800 291.600 123.600 292.400 ;
        RECT 135.600 289.600 136.400 290.400 ;
        RECT 143.600 293.600 144.400 294.400 ;
        RECT 162.800 297.600 163.600 298.400 ;
        RECT 150.000 291.600 150.800 292.400 ;
        RECT 153.200 291.600 154.000 292.400 ;
        RECT 145.200 289.600 146.000 290.400 ;
        RECT 150.000 283.600 150.800 284.400 ;
        RECT 162.800 289.600 163.600 290.400 ;
        RECT 177.200 297.600 178.000 298.400 ;
        RECT 175.600 293.600 176.400 294.400 ;
        RECT 167.600 289.600 168.400 290.400 ;
        RECT 172.400 291.600 173.200 292.400 ;
        RECT 182.000 289.600 182.800 290.400 ;
        RECT 196.400 293.600 197.200 294.400 ;
        RECT 204.400 293.600 205.200 294.400 ;
        RECT 230.000 297.600 230.800 298.400 ;
        RECT 238.000 297.600 238.800 298.400 ;
        RECT 199.600 291.600 200.400 292.400 ;
        RECT 206.000 291.600 206.800 292.400 ;
        RECT 223.600 293.600 224.400 294.400 ;
        RECT 231.600 293.600 232.400 294.400 ;
        RECT 239.600 293.600 240.400 294.400 ;
        RECT 242.800 293.600 243.600 294.400 ;
        RECT 214.000 289.600 214.800 290.400 ;
        RECT 225.200 291.600 226.000 292.400 ;
        RECT 226.800 291.600 227.600 292.400 ;
        RECT 233.200 291.600 234.000 292.400 ;
        RECT 234.800 291.600 235.600 292.400 ;
        RECT 241.200 291.600 242.000 292.400 ;
        RECT 255.600 297.600 256.400 298.400 ;
        RECT 254.000 293.600 254.800 294.400 ;
        RECT 250.800 283.600 251.600 284.400 ;
        RECT 292.400 295.600 293.200 296.400 ;
        RECT 294.000 294.200 294.800 295.000 ;
        RECT 305.200 291.600 306.000 292.400 ;
        RECT 266.800 289.600 267.600 290.400 ;
        RECT 276.400 283.600 277.200 284.400 ;
        RECT 287.600 286.800 288.400 287.600 ;
        RECT 290.800 286.200 291.600 287.000 ;
        RECT 286.000 284.200 286.800 285.000 ;
        RECT 287.600 284.200 288.400 285.000 ;
        RECT 289.200 284.200 290.000 285.000 ;
        RECT 294.000 286.200 294.800 287.000 ;
        RECT 297.200 286.200 298.000 287.000 ;
        RECT 354.800 295.600 355.600 296.400 ;
        RECT 298.800 284.200 299.600 285.000 ;
        RECT 300.400 284.200 301.200 285.000 ;
        RECT 327.600 291.600 328.400 292.400 ;
        RECT 337.200 293.600 338.000 294.400 ;
        RECT 346.800 291.600 347.600 292.400 ;
        RECT 370.800 297.600 371.600 298.400 ;
        RECT 367.600 293.600 368.400 294.400 ;
        RECT 369.200 291.600 370.000 292.400 ;
        RECT 374.000 297.600 374.800 298.400 ;
        RECT 410.800 297.600 411.600 298.400 ;
        RECT 388.400 289.600 389.200 290.400 ;
        RECT 396.400 291.600 397.200 292.400 ;
        RECT 398.000 289.600 398.800 290.400 ;
        RECT 399.600 289.600 400.400 290.400 ;
        RECT 407.600 289.600 408.400 290.400 ;
        RECT 414.000 291.600 414.800 292.400 ;
        RECT 430.000 297.600 430.800 298.400 ;
        RECT 438.000 297.600 438.800 298.400 ;
        RECT 422.000 291.600 422.800 292.400 ;
        RECT 436.400 293.600 437.200 294.400 ;
        RECT 441.200 291.600 442.000 292.400 ;
        RECT 442.800 289.600 443.600 290.400 ;
        RECT 449.200 293.600 450.000 294.400 ;
        RECT 468.400 295.600 469.200 296.400 ;
        RECT 470.000 294.200 470.800 295.000 ;
        RECT 487.600 297.600 488.400 298.400 ;
        RECT 500.400 297.600 501.200 298.400 ;
        RECT 460.400 291.600 461.200 292.400 ;
        RECT 479.600 291.600 480.400 292.400 ;
        RECT 452.400 283.600 453.200 284.400 ;
        RECT 463.600 286.800 464.400 287.600 ;
        RECT 466.800 286.200 467.600 287.000 ;
        RECT 462.000 284.200 462.800 285.000 ;
        RECT 463.600 284.200 464.400 285.000 ;
        RECT 465.200 284.200 466.000 285.000 ;
        RECT 470.000 286.200 470.800 287.000 ;
        RECT 473.200 286.200 474.000 287.000 ;
        RECT 489.200 293.600 490.000 294.400 ;
        RECT 492.400 293.600 493.200 294.400 ;
        RECT 490.800 291.600 491.600 292.400 ;
        RECT 474.800 284.200 475.600 285.000 ;
        RECT 476.400 284.200 477.200 285.000 ;
        RECT 510.000 297.600 510.800 298.400 ;
        RECT 506.800 291.600 507.600 292.400 ;
        RECT 508.400 289.600 509.200 290.400 ;
        RECT 506.800 287.600 507.600 288.400 ;
        RECT 530.800 295.600 531.600 296.400 ;
        RECT 532.400 294.200 533.200 295.000 ;
        RECT 522.800 291.600 523.600 292.400 ;
        RECT 526.000 286.800 526.800 287.600 ;
        RECT 529.200 286.200 530.000 287.000 ;
        RECT 524.400 284.200 525.200 285.000 ;
        RECT 526.000 284.200 526.800 285.000 ;
        RECT 527.600 284.200 528.400 285.000 ;
        RECT 532.400 286.200 533.200 287.000 ;
        RECT 535.600 286.200 536.400 287.000 ;
        RECT 537.200 284.200 538.000 285.000 ;
        RECT 538.800 284.200 539.600 285.000 ;
        RECT 2.800 277.600 3.600 278.400 ;
        RECT 14.000 274.400 14.800 275.200 ;
        RECT 17.200 275.000 18.000 275.800 ;
        RECT 12.400 272.400 13.200 273.200 ;
        RECT 22.000 267.600 22.800 268.400 ;
        RECT 18.800 265.600 19.600 266.400 ;
        RECT 38.000 269.600 38.800 270.400 ;
        RECT 41.200 269.600 42.000 270.400 ;
        RECT 12.400 264.200 13.200 265.000 ;
        RECT 14.000 264.200 14.800 265.000 ;
        RECT 15.600 264.200 16.400 265.000 ;
        RECT 17.200 264.200 18.000 265.000 ;
        RECT 20.400 264.200 21.200 265.000 ;
        RECT 23.600 264.200 24.400 265.000 ;
        RECT 25.200 264.200 26.000 265.000 ;
        RECT 26.800 264.200 27.600 265.000 ;
        RECT 47.600 267.600 48.400 268.400 ;
        RECT 46.000 263.600 46.800 264.400 ;
        RECT 52.400 265.600 53.200 266.400 ;
        RECT 66.800 277.600 67.600 278.400 ;
        RECT 63.600 267.600 64.400 268.400 ;
        RECT 73.200 269.600 74.000 270.400 ;
        RECT 68.400 267.600 69.200 268.400 ;
        RECT 74.800 267.600 75.600 268.400 ;
        RECT 62.000 263.600 62.800 264.400 ;
        RECT 70.000 263.600 70.800 264.400 ;
        RECT 76.400 265.600 77.200 266.400 ;
        RECT 87.600 265.600 88.400 266.400 ;
        RECT 89.200 263.600 90.000 264.400 ;
        RECT 108.400 275.000 109.200 275.800 ;
        RECT 105.200 273.600 106.000 274.400 ;
        RECT 110.000 272.400 110.800 273.200 ;
        RECT 134.000 277.600 134.800 278.400 ;
        RECT 114.800 269.600 115.600 270.400 ;
        RECT 98.800 268.200 99.600 269.000 ;
        RECT 108.400 268.600 109.200 269.400 ;
        RECT 103.600 267.600 104.400 268.400 ;
        RECT 142.000 269.600 142.800 270.400 ;
        RECT 98.800 264.200 99.600 265.000 ;
        RECT 100.400 264.200 101.200 265.000 ;
        RECT 102.000 264.200 102.800 265.000 ;
        RECT 105.200 264.200 106.000 265.000 ;
        RECT 108.400 264.200 109.200 265.000 ;
        RECT 110.000 264.200 110.800 265.000 ;
        RECT 111.600 264.200 112.400 265.000 ;
        RECT 113.200 264.200 114.000 265.000 ;
        RECT 148.400 269.600 149.200 270.400 ;
        RECT 158.000 265.600 158.800 266.400 ;
        RECT 174.000 277.600 174.800 278.400 ;
        RECT 167.600 267.600 168.400 268.400 ;
        RECT 175.600 273.600 176.400 274.400 ;
        RECT 172.400 271.600 173.200 272.400 ;
        RECT 166.000 263.600 166.800 264.400 ;
        RECT 186.800 273.600 187.600 274.400 ;
        RECT 198.000 277.600 198.800 278.400 ;
        RECT 199.600 273.600 200.400 274.400 ;
        RECT 196.400 271.600 197.200 272.400 ;
        RECT 193.200 269.600 194.000 270.400 ;
        RECT 182.000 267.600 182.800 268.400 ;
        RECT 188.400 267.600 189.200 268.400 ;
        RECT 191.600 267.600 192.400 268.400 ;
        RECT 194.800 267.600 195.600 268.400 ;
        RECT 202.800 269.600 203.600 270.400 ;
        RECT 204.400 265.600 205.200 266.400 ;
        RECT 206.000 265.600 206.800 266.400 ;
        RECT 214.000 265.600 214.800 266.400 ;
        RECT 231.600 269.600 232.400 270.400 ;
        RECT 238.000 273.600 238.800 274.400 ;
        RECT 226.800 265.600 227.600 266.400 ;
        RECT 257.200 277.600 258.000 278.400 ;
        RECT 249.200 269.600 250.000 270.400 ;
        RECT 255.600 269.600 256.400 270.400 ;
        RECT 281.200 274.400 282.000 275.200 ;
        RECT 284.400 275.000 285.200 275.800 ;
        RECT 279.600 272.400 280.400 273.200 ;
        RECT 258.800 269.600 259.600 270.400 ;
        RECT 295.600 271.200 296.400 272.000 ;
        RECT 234.800 263.600 235.600 264.400 ;
        RECT 244.400 265.600 245.200 266.400 ;
        RECT 260.400 267.600 261.200 268.400 ;
        RECT 269.800 267.600 270.600 268.400 ;
        RECT 252.400 263.600 253.200 264.400 ;
        RECT 289.200 267.600 290.000 268.400 ;
        RECT 286.000 265.600 286.800 266.400 ;
        RECT 279.600 264.200 280.400 265.000 ;
        RECT 281.200 264.200 282.000 265.000 ;
        RECT 282.800 264.200 283.600 265.000 ;
        RECT 284.400 264.200 285.200 265.000 ;
        RECT 287.600 264.200 288.400 265.000 ;
        RECT 290.800 264.200 291.600 265.000 ;
        RECT 292.400 264.200 293.200 265.000 ;
        RECT 294.000 264.200 294.800 265.000 ;
        RECT 321.200 275.000 322.000 275.800 ;
        RECT 318.000 273.600 318.800 274.400 ;
        RECT 322.800 272.400 323.600 273.200 ;
        RECT 306.800 271.600 307.600 272.400 ;
        RECT 335.600 273.600 336.400 274.400 ;
        RECT 311.600 268.200 312.400 269.000 ;
        RECT 321.200 268.600 322.000 269.400 ;
        RECT 316.400 267.600 317.200 268.400 ;
        RECT 311.600 264.200 312.400 265.000 ;
        RECT 313.200 264.200 314.000 265.000 ;
        RECT 314.800 264.200 315.600 265.000 ;
        RECT 318.000 264.200 318.800 265.000 ;
        RECT 321.200 264.200 322.000 265.000 ;
        RECT 322.800 264.200 323.600 265.000 ;
        RECT 324.400 264.200 325.200 265.000 ;
        RECT 326.000 264.200 326.800 265.000 ;
        RECT 340.400 263.600 341.200 264.400 ;
        RECT 366.000 275.000 366.800 275.800 ;
        RECT 362.800 273.600 363.600 274.400 ;
        RECT 367.600 272.400 368.400 273.200 ;
        RECT 354.800 271.200 355.600 272.000 ;
        RECT 356.400 268.200 357.200 269.000 ;
        RECT 366.000 268.600 366.800 269.400 ;
        RECT 346.800 263.600 347.600 264.400 ;
        RECT 361.200 267.600 362.000 268.400 ;
        RECT 356.400 264.200 357.200 265.000 ;
        RECT 358.000 264.200 358.800 265.000 ;
        RECT 359.600 264.200 360.400 265.000 ;
        RECT 362.800 264.200 363.600 265.000 ;
        RECT 366.000 264.200 366.800 265.000 ;
        RECT 367.600 264.200 368.400 265.000 ;
        RECT 369.200 264.200 370.000 265.000 ;
        RECT 370.800 264.200 371.600 265.000 ;
        RECT 401.200 275.000 402.000 275.800 ;
        RECT 398.000 273.600 398.800 274.400 ;
        RECT 402.800 272.400 403.600 273.200 ;
        RECT 391.600 268.200 392.400 269.000 ;
        RECT 401.200 268.600 402.000 269.400 ;
        RECT 380.400 263.600 381.200 264.400 ;
        RECT 396.400 267.600 397.200 268.400 ;
        RECT 391.600 264.200 392.400 265.000 ;
        RECT 393.200 264.200 394.000 265.000 ;
        RECT 394.800 264.200 395.600 265.000 ;
        RECT 398.000 264.200 398.800 265.000 ;
        RECT 401.200 264.200 402.000 265.000 ;
        RECT 402.800 264.200 403.600 265.000 ;
        RECT 404.400 264.200 405.200 265.000 ;
        RECT 406.000 264.200 406.800 265.000 ;
        RECT 434.800 269.600 435.600 270.400 ;
        RECT 441.200 269.600 442.000 270.400 ;
        RECT 442.800 269.600 443.600 270.400 ;
        RECT 422.000 265.600 422.800 266.400 ;
        RECT 430.000 265.600 430.800 266.400 ;
        RECT 420.400 263.600 421.200 264.400 ;
        RECT 436.400 267.600 437.200 268.400 ;
        RECT 446.000 265.600 446.800 266.400 ;
        RECT 447.600 263.600 448.400 264.400 ;
        RECT 454.000 277.600 454.800 278.400 ;
        RECT 449.200 267.600 450.000 268.400 ;
        RECT 465.200 274.400 466.000 275.200 ;
        RECT 468.400 275.000 469.200 275.800 ;
        RECT 489.200 277.600 490.000 278.400 ;
        RECT 463.600 272.400 464.400 273.200 ;
        RECT 462.000 269.600 462.800 270.400 ;
        RECT 473.200 267.600 474.000 268.400 ;
        RECT 470.000 265.600 470.800 266.400 ;
        RECT 463.600 264.200 464.400 265.000 ;
        RECT 465.200 264.200 466.000 265.000 ;
        RECT 466.800 264.200 467.600 265.000 ;
        RECT 468.400 264.200 469.200 265.000 ;
        RECT 471.600 264.200 472.400 265.000 ;
        RECT 474.800 264.200 475.600 265.000 ;
        RECT 476.400 264.200 477.200 265.000 ;
        RECT 478.000 264.200 478.800 265.000 ;
        RECT 500.400 274.400 501.200 275.200 ;
        RECT 503.600 275.000 504.400 275.800 ;
        RECT 498.800 272.400 499.600 273.200 ;
        RECT 497.200 269.600 498.000 270.400 ;
        RECT 508.400 267.600 509.200 268.400 ;
        RECT 505.200 265.600 506.000 266.400 ;
        RECT 498.800 264.200 499.600 265.000 ;
        RECT 500.400 264.200 501.200 265.000 ;
        RECT 502.000 264.200 502.800 265.000 ;
        RECT 503.600 264.200 504.400 265.000 ;
        RECT 506.800 264.200 507.600 265.000 ;
        RECT 510.000 264.200 510.800 265.000 ;
        RECT 511.600 264.200 512.400 265.000 ;
        RECT 513.200 264.200 514.000 265.000 ;
        RECT 527.600 267.600 528.400 268.400 ;
        RECT 524.400 265.600 525.200 266.400 ;
        RECT 526.000 266.200 526.800 267.000 ;
        RECT 522.800 263.600 523.600 264.400 ;
        RECT 7.600 251.600 8.400 252.400 ;
        RECT 14.000 253.600 14.800 254.400 ;
        RECT 30.000 257.600 30.800 258.400 ;
        RECT 25.200 253.600 26.000 254.400 ;
        RECT 12.400 249.600 13.200 250.400 ;
        RECT 10.800 247.600 11.600 248.400 ;
        RECT 7.600 243.600 8.400 244.400 ;
        RECT 20.400 251.600 21.200 252.400 ;
        RECT 44.400 255.600 45.200 256.400 ;
        RECT 34.800 251.600 35.600 252.400 ;
        RECT 38.000 251.600 38.800 252.400 ;
        RECT 18.800 243.600 19.600 244.400 ;
        RECT 30.000 243.600 30.800 244.400 ;
        RECT 36.400 249.600 37.200 250.400 ;
        RECT 39.600 243.600 40.400 244.400 ;
        RECT 57.200 257.600 58.000 258.400 ;
        RECT 46.000 249.600 46.800 250.400 ;
        RECT 52.400 243.600 53.200 244.400 ;
        RECT 57.200 249.600 58.000 250.400 ;
        RECT 58.800 249.600 59.600 250.400 ;
        RECT 81.200 255.600 82.000 256.400 ;
        RECT 97.200 255.600 98.000 256.400 ;
        RECT 98.800 254.200 99.600 255.000 ;
        RECT 110.000 251.600 110.800 252.400 ;
        RECT 92.400 246.800 93.200 247.600 ;
        RECT 95.600 246.200 96.400 247.000 ;
        RECT 90.800 244.200 91.600 245.000 ;
        RECT 92.400 244.200 93.200 245.000 ;
        RECT 94.000 244.200 94.800 245.000 ;
        RECT 98.800 246.200 99.600 247.000 ;
        RECT 102.000 246.200 102.800 247.000 ;
        RECT 122.800 257.600 123.600 258.400 ;
        RECT 137.200 257.600 138.000 258.400 ;
        RECT 142.000 257.600 142.800 258.400 ;
        RECT 122.800 253.600 123.600 254.400 ;
        RECT 138.800 253.600 139.600 254.400 ;
        RECT 121.200 251.600 122.000 252.400 ;
        RECT 140.400 251.600 141.200 252.400 ;
        RECT 103.600 244.200 104.400 245.000 ;
        RECT 105.200 244.200 106.000 245.000 ;
        RECT 153.200 253.000 154.000 253.800 ;
        RECT 162.800 252.600 163.600 253.400 ;
        RECT 177.200 257.600 178.000 258.400 ;
        RECT 182.000 257.600 182.800 258.400 ;
        RECT 158.000 251.600 158.800 252.400 ;
        RECT 154.800 248.800 155.600 249.600 ;
        RECT 159.600 247.600 160.400 248.400 ;
        RECT 156.400 246.200 157.200 247.000 ;
        RECT 153.200 244.200 154.000 245.000 ;
        RECT 154.800 244.200 155.600 245.000 ;
        RECT 159.600 246.200 160.400 247.000 ;
        RECT 162.800 246.200 163.600 247.000 ;
        RECT 164.400 244.200 165.200 245.000 ;
        RECT 166.000 244.200 166.800 245.000 ;
        RECT 167.600 244.200 168.400 245.000 ;
        RECT 188.400 257.600 189.200 258.400 ;
        RECT 190.000 257.600 190.800 258.400 ;
        RECT 188.400 249.600 189.200 250.400 ;
        RECT 207.600 257.600 208.400 258.400 ;
        RECT 223.600 255.600 224.400 256.400 ;
        RECT 225.200 254.200 226.000 255.000 ;
        RECT 242.800 257.600 243.600 258.400 ;
        RECT 233.200 251.600 234.000 252.400 ;
        RECT 218.800 246.800 219.600 247.600 ;
        RECT 222.000 246.200 222.800 247.000 ;
        RECT 217.200 244.200 218.000 245.000 ;
        RECT 218.800 244.200 219.600 245.000 ;
        RECT 220.400 244.200 221.200 245.000 ;
        RECT 225.200 246.200 226.000 247.000 ;
        RECT 228.400 246.200 229.200 247.000 ;
        RECT 241.200 249.600 242.000 250.400 ;
        RECT 230.000 244.200 230.800 245.000 ;
        RECT 231.600 244.200 232.400 245.000 ;
        RECT 263.600 255.600 264.400 256.400 ;
        RECT 265.200 254.200 266.000 255.000 ;
        RECT 289.200 257.600 290.000 258.400 ;
        RECT 247.600 243.600 248.400 244.400 ;
        RECT 258.800 246.800 259.600 247.600 ;
        RECT 262.000 246.200 262.800 247.000 ;
        RECT 257.200 244.200 258.000 245.000 ;
        RECT 258.800 244.200 259.600 245.000 ;
        RECT 260.400 244.200 261.200 245.000 ;
        RECT 265.200 246.200 266.000 247.000 ;
        RECT 268.400 246.200 269.200 247.000 ;
        RECT 305.200 255.600 306.000 256.400 ;
        RECT 306.800 254.200 307.600 255.000 ;
        RECT 322.800 257.600 323.600 258.400 ;
        RECT 337.200 257.600 338.000 258.400 ;
        RECT 270.000 244.200 270.800 245.000 ;
        RECT 271.600 244.200 272.400 245.000 ;
        RECT 300.400 246.800 301.200 247.600 ;
        RECT 303.600 246.200 304.400 247.000 ;
        RECT 298.800 244.200 299.600 245.000 ;
        RECT 300.400 244.200 301.200 245.000 ;
        RECT 302.000 244.200 302.800 245.000 ;
        RECT 306.800 246.200 307.600 247.000 ;
        RECT 310.000 246.200 310.800 247.000 ;
        RECT 311.600 244.200 312.400 245.000 ;
        RECT 313.200 244.200 314.000 245.000 ;
        RECT 348.400 257.600 349.200 258.400 ;
        RECT 358.000 253.000 358.800 253.800 ;
        RECT 348.400 249.600 349.200 250.400 ;
        RECT 367.600 252.600 368.400 253.400 ;
        RECT 354.800 251.600 355.600 252.400 ;
        RECT 362.800 251.600 363.600 252.400 ;
        RECT 359.600 248.800 360.400 249.600 ;
        RECT 364.400 247.600 365.200 248.400 ;
        RECT 361.200 246.200 362.000 247.000 ;
        RECT 358.000 244.200 358.800 245.000 ;
        RECT 359.600 244.200 360.400 245.000 ;
        RECT 364.400 246.200 365.200 247.000 ;
        RECT 367.600 246.200 368.400 247.000 ;
        RECT 369.200 244.200 370.000 245.000 ;
        RECT 370.800 244.200 371.600 245.000 ;
        RECT 372.400 244.200 373.200 245.000 ;
        RECT 406.000 255.600 406.800 256.400 ;
        RECT 407.600 254.200 408.400 255.000 ;
        RECT 418.800 251.600 419.600 252.400 ;
        RECT 385.200 243.600 386.000 244.400 ;
        RECT 401.200 246.800 402.000 247.600 ;
        RECT 404.400 246.200 405.200 247.000 ;
        RECT 399.600 244.200 400.400 245.000 ;
        RECT 401.200 244.200 402.000 245.000 ;
        RECT 402.800 244.200 403.600 245.000 ;
        RECT 407.600 246.200 408.400 247.000 ;
        RECT 410.800 246.200 411.600 247.000 ;
        RECT 412.400 244.200 413.200 245.000 ;
        RECT 414.000 244.200 414.800 245.000 ;
        RECT 434.600 253.600 435.400 254.400 ;
        RECT 450.800 255.600 451.600 256.400 ;
        RECT 452.400 254.200 453.200 255.000 ;
        RECT 442.800 251.600 443.600 252.400 ;
        RECT 462.000 251.600 462.800 252.400 ;
        RECT 431.600 245.600 432.400 246.400 ;
        RECT 446.000 246.800 446.800 247.600 ;
        RECT 449.200 246.200 450.000 247.000 ;
        RECT 444.400 244.200 445.200 245.000 ;
        RECT 446.000 244.200 446.800 245.000 ;
        RECT 447.600 244.200 448.400 245.000 ;
        RECT 452.400 246.200 453.200 247.000 ;
        RECT 455.600 246.200 456.400 247.000 ;
        RECT 471.600 253.600 472.400 254.400 ;
        RECT 470.000 251.600 470.800 252.400 ;
        RECT 473.200 251.600 474.000 252.400 ;
        RECT 474.800 251.600 475.600 252.400 ;
        RECT 487.600 253.000 488.400 253.800 ;
        RECT 457.200 244.200 458.000 245.000 ;
        RECT 458.800 244.200 459.600 245.000 ;
        RECT 497.200 252.600 498.000 253.400 ;
        RECT 482.800 251.600 483.600 252.400 ;
        RECT 511.800 251.600 512.600 252.400 ;
        RECT 527.600 253.600 528.400 254.400 ;
        RECT 489.200 248.800 490.000 249.600 ;
        RECT 494.000 247.600 494.800 248.400 ;
        RECT 490.800 246.200 491.600 247.000 ;
        RECT 487.600 244.200 488.400 245.000 ;
        RECT 489.200 244.200 490.000 245.000 ;
        RECT 494.000 246.200 494.800 247.000 ;
        RECT 497.200 246.200 498.000 247.000 ;
        RECT 498.800 244.200 499.600 245.000 ;
        RECT 500.400 244.200 501.200 245.000 ;
        RECT 502.000 244.200 502.800 245.000 ;
        RECT 534.000 252.200 534.800 253.000 ;
        RECT 542.000 251.800 542.800 252.600 ;
        RECT 546.800 250.200 547.600 251.000 ;
        RECT 14.000 234.400 14.800 235.200 ;
        RECT 17.200 235.000 18.000 235.800 ;
        RECT 41.200 237.600 42.000 238.400 ;
        RECT 12.400 232.400 13.200 233.200 ;
        RECT 2.800 223.600 3.600 224.400 ;
        RECT 39.600 233.600 40.400 234.400 ;
        RECT 36.400 231.600 37.200 232.400 ;
        RECT 22.000 227.600 22.800 228.400 ;
        RECT 18.800 225.600 19.600 226.400 ;
        RECT 44.400 229.600 45.200 230.400 ;
        RECT 47.600 229.600 48.400 230.400 ;
        RECT 12.400 224.200 13.200 225.000 ;
        RECT 14.000 224.200 14.800 225.000 ;
        RECT 15.600 224.200 16.400 225.000 ;
        RECT 17.200 224.200 18.000 225.000 ;
        RECT 20.400 224.200 21.200 225.000 ;
        RECT 23.600 224.200 24.400 225.000 ;
        RECT 25.200 224.200 26.000 225.000 ;
        RECT 26.800 224.200 27.600 225.000 ;
        RECT 54.000 225.600 54.800 226.400 ;
        RECT 68.400 233.600 69.200 234.400 ;
        RECT 71.600 231.600 72.400 232.400 ;
        RECT 78.000 233.600 78.800 234.400 ;
        RECT 70.000 229.600 70.800 230.400 ;
        RECT 65.200 227.600 66.000 228.400 ;
        RECT 116.400 234.400 117.200 235.200 ;
        RECT 119.600 235.000 120.400 235.800 ;
        RECT 146.800 237.600 147.600 238.400 ;
        RECT 114.800 232.400 115.600 233.200 ;
        RECT 86.000 225.600 86.800 226.400 ;
        RECT 81.200 223.600 82.000 224.400 ;
        RECT 105.000 229.600 105.800 230.400 ;
        RECT 95.600 223.600 96.400 224.400 ;
        RECT 98.800 223.600 99.600 224.400 ;
        RECT 124.400 227.600 125.200 228.400 ;
        RECT 121.200 225.600 122.000 226.400 ;
        RECT 114.800 224.200 115.600 225.000 ;
        RECT 116.400 224.200 117.200 225.000 ;
        RECT 118.000 224.200 118.800 225.000 ;
        RECT 119.600 224.200 120.400 225.000 ;
        RECT 122.800 224.200 123.600 225.000 ;
        RECT 126.000 224.200 126.800 225.000 ;
        RECT 127.600 224.200 128.400 225.000 ;
        RECT 129.200 224.200 130.000 225.000 ;
        RECT 145.200 227.600 146.000 228.400 ;
        RECT 146.800 223.600 147.600 224.400 ;
        RECT 150.000 233.600 150.800 234.400 ;
        RECT 156.400 231.600 157.200 232.400 ;
        RECT 161.200 229.600 162.000 230.400 ;
        RECT 162.800 229.600 163.600 230.400 ;
        RECT 151.600 225.600 152.400 226.400 ;
        RECT 158.000 227.600 158.800 228.400 ;
        RECT 175.600 237.600 176.400 238.400 ;
        RECT 169.200 227.600 170.000 228.400 ;
        RECT 182.000 237.600 182.800 238.400 ;
        RECT 178.800 231.600 179.600 232.400 ;
        RECT 177.200 227.600 178.000 228.400 ;
        RECT 194.800 237.600 195.600 238.400 ;
        RECT 186.800 227.600 187.600 228.400 ;
        RECT 194.800 229.600 195.600 230.400 ;
        RECT 199.600 229.600 200.400 230.400 ;
        RECT 217.200 234.400 218.000 235.200 ;
        RECT 220.400 235.000 221.200 235.800 ;
        RECT 215.600 232.400 216.400 233.200 ;
        RECT 196.400 227.600 197.200 228.400 ;
        RECT 206.000 223.600 206.800 224.400 ;
        RECT 225.200 227.600 226.000 228.400 ;
        RECT 222.000 225.600 222.800 226.400 ;
        RECT 215.600 224.200 216.400 225.000 ;
        RECT 217.200 224.200 218.000 225.000 ;
        RECT 218.800 224.200 219.600 225.000 ;
        RECT 220.400 224.200 221.200 225.000 ;
        RECT 223.600 224.200 224.400 225.000 ;
        RECT 226.800 224.200 227.600 225.000 ;
        RECT 228.400 224.200 229.200 225.000 ;
        RECT 230.000 224.200 230.800 225.000 ;
        RECT 252.400 234.400 253.200 235.200 ;
        RECT 255.600 235.000 256.400 235.800 ;
        RECT 250.800 232.400 251.600 233.200 ;
        RECT 249.200 229.600 250.000 230.400 ;
        RECT 260.400 227.600 261.200 228.400 ;
        RECT 257.200 225.600 258.000 226.400 ;
        RECT 250.800 224.200 251.600 225.000 ;
        RECT 252.400 224.200 253.200 225.000 ;
        RECT 254.000 224.200 254.800 225.000 ;
        RECT 255.600 224.200 256.400 225.000 ;
        RECT 258.800 224.200 259.600 225.000 ;
        RECT 262.000 224.200 262.800 225.000 ;
        RECT 263.600 224.200 264.400 225.000 ;
        RECT 265.200 224.200 266.000 225.000 ;
        RECT 282.800 227.600 283.600 228.400 ;
        RECT 297.200 234.400 298.000 235.200 ;
        RECT 300.400 235.000 301.200 235.800 ;
        RECT 295.600 232.400 296.400 233.200 ;
        RECT 311.600 231.200 312.400 232.000 ;
        RECT 286.000 223.600 286.800 224.400 ;
        RECT 305.200 227.600 306.000 228.400 ;
        RECT 302.000 225.600 302.800 226.400 ;
        RECT 321.200 229.600 322.000 230.400 ;
        RECT 327.600 229.600 328.400 230.400 ;
        RECT 361.200 237.600 362.000 238.400 ;
        RECT 295.600 224.200 296.400 225.000 ;
        RECT 297.200 224.200 298.000 225.000 ;
        RECT 298.800 224.200 299.600 225.000 ;
        RECT 300.400 224.200 301.200 225.000 ;
        RECT 303.600 224.200 304.400 225.000 ;
        RECT 306.800 224.200 307.600 225.000 ;
        RECT 308.400 224.200 309.200 225.000 ;
        RECT 310.000 224.200 310.800 225.000 ;
        RECT 329.200 227.600 330.000 228.400 ;
        RECT 337.200 227.600 338.000 228.400 ;
        RECT 343.600 227.600 344.400 228.400 ;
        RECT 356.400 229.600 357.200 230.400 ;
        RECT 353.200 227.600 354.000 228.400 ;
        RECT 378.800 237.600 379.600 238.400 ;
        RECT 390.000 234.400 390.800 235.200 ;
        RECT 393.200 235.000 394.000 235.800 ;
        RECT 388.400 232.400 389.200 233.200 ;
        RECT 370.800 227.600 371.600 228.400 ;
        RECT 386.800 229.600 387.600 230.400 ;
        RECT 378.800 225.600 379.600 226.400 ;
        RECT 398.000 227.600 398.800 228.400 ;
        RECT 394.800 225.600 395.600 226.400 ;
        RECT 388.400 224.200 389.200 225.000 ;
        RECT 390.000 224.200 390.800 225.000 ;
        RECT 391.600 224.200 392.400 225.000 ;
        RECT 393.200 224.200 394.000 225.000 ;
        RECT 396.400 224.200 397.200 225.000 ;
        RECT 399.600 224.200 400.400 225.000 ;
        RECT 401.200 224.200 402.000 225.000 ;
        RECT 402.800 224.200 403.600 225.000 ;
        RECT 431.600 233.600 432.400 234.400 ;
        RECT 441.200 237.600 442.000 238.400 ;
        RECT 417.200 229.600 418.000 230.400 ;
        RECT 428.400 231.600 429.200 232.400 ;
        RECT 412.400 225.600 413.200 226.400 ;
        RECT 418.800 227.600 419.600 228.400 ;
        RECT 414.000 223.600 414.800 224.400 ;
        RECT 438.000 225.600 438.800 226.400 ;
        RECT 446.000 227.600 446.800 228.400 ;
        RECT 458.800 237.600 459.600 238.400 ;
        RECT 465.200 237.600 466.000 238.400 ;
        RECT 460.400 233.600 461.200 234.400 ;
        RECT 466.800 233.600 467.600 234.400 ;
        RECT 457.200 231.600 458.000 232.400 ;
        RECT 463.600 231.600 464.400 232.400 ;
        RECT 452.400 229.600 453.200 230.400 ;
        RECT 454.000 229.600 454.800 230.400 ;
        RECT 487.600 231.600 488.400 232.400 ;
        RECT 470.000 225.600 470.800 226.400 ;
        RECT 474.800 225.600 475.600 226.400 ;
        RECT 508.400 234.400 509.200 235.200 ;
        RECT 511.600 235.000 512.400 235.800 ;
        RECT 506.800 232.400 507.600 233.200 ;
        RECT 497.000 227.600 497.800 228.400 ;
        RECT 505.200 229.600 506.000 230.400 ;
        RECT 516.400 227.600 517.200 228.400 ;
        RECT 513.200 225.600 514.000 226.400 ;
        RECT 506.800 224.200 507.600 225.000 ;
        RECT 508.400 224.200 509.200 225.000 ;
        RECT 510.000 224.200 510.800 225.000 ;
        RECT 511.600 224.200 512.400 225.000 ;
        RECT 514.800 224.200 515.600 225.000 ;
        RECT 518.000 224.200 518.800 225.000 ;
        RECT 519.600 224.200 520.400 225.000 ;
        RECT 521.200 224.200 522.000 225.000 ;
        RECT 546.800 229.600 547.600 230.400 ;
        RECT 542.000 225.600 542.800 226.400 ;
        RECT 532.400 223.600 533.200 224.400 ;
        RECT 15.600 217.600 16.400 218.400 ;
        RECT 12.400 213.600 13.200 214.400 ;
        RECT 9.200 211.600 10.000 212.400 ;
        RECT 17.200 211.600 18.000 212.400 ;
        RECT 2.800 203.600 3.600 204.400 ;
        RECT 18.800 209.600 19.600 210.400 ;
        RECT 30.000 213.600 30.800 214.400 ;
        RECT 26.800 211.600 27.600 212.400 ;
        RECT 36.400 213.600 37.200 214.400 ;
        RECT 26.800 205.600 27.600 206.400 ;
        RECT 57.200 217.600 58.000 218.400 ;
        RECT 46.000 211.600 46.800 212.400 ;
        RECT 86.000 217.600 86.800 218.400 ;
        RECT 95.600 217.600 96.400 218.400 ;
        RECT 41.200 203.600 42.000 204.400 ;
        RECT 46.000 203.600 46.800 204.400 ;
        RECT 63.600 203.600 64.400 204.400 ;
        RECT 73.200 203.600 74.000 204.400 ;
        RECT 89.200 213.600 90.000 214.400 ;
        RECT 94.000 213.600 94.800 214.400 ;
        RECT 87.600 209.600 88.400 210.400 ;
        RECT 100.400 209.600 101.200 210.400 ;
        RECT 102.000 209.600 102.800 210.400 ;
        RECT 124.400 213.000 125.200 213.800 ;
        RECT 108.400 209.600 109.200 210.400 ;
        RECT 134.000 212.600 134.800 213.400 ;
        RECT 129.200 211.600 130.000 212.400 ;
        RECT 140.400 211.600 141.200 212.400 ;
        RECT 158.000 213.600 158.800 214.400 ;
        RECT 175.600 217.600 176.400 218.400 ;
        RECT 164.400 213.600 165.200 214.400 ;
        RECT 151.600 211.600 152.400 212.400 ;
        RECT 126.000 208.800 126.800 209.600 ;
        RECT 130.800 207.600 131.600 208.400 ;
        RECT 127.600 206.200 128.400 207.000 ;
        RECT 124.400 204.200 125.200 205.000 ;
        RECT 126.000 204.200 126.800 205.000 ;
        RECT 130.800 206.200 131.600 207.000 ;
        RECT 134.000 206.200 134.800 207.000 ;
        RECT 135.600 204.200 136.400 205.000 ;
        RECT 137.200 204.200 138.000 205.000 ;
        RECT 138.800 204.200 139.600 205.000 ;
        RECT 159.600 209.600 160.400 210.400 ;
        RECT 174.000 211.600 174.800 212.400 ;
        RECT 166.000 209.600 166.800 210.400 ;
        RECT 178.800 213.600 179.600 214.400 ;
        RECT 185.200 211.600 186.000 212.400 ;
        RECT 198.000 211.600 198.800 212.400 ;
        RECT 175.600 203.600 176.400 204.400 ;
        RECT 194.800 209.600 195.600 210.400 ;
        RECT 212.400 213.600 213.200 214.400 ;
        RECT 204.400 211.600 205.200 212.400 ;
        RECT 207.600 211.600 208.400 212.400 ;
        RECT 199.600 209.600 200.400 210.400 ;
        RECT 214.000 211.600 214.800 212.400 ;
        RECT 201.200 203.600 202.000 204.400 ;
        RECT 215.600 209.600 216.400 210.400 ;
        RECT 217.200 209.600 218.000 210.400 ;
        RECT 225.200 209.600 226.000 210.400 ;
        RECT 231.600 209.600 232.400 210.400 ;
        RECT 263.600 215.600 264.400 216.400 ;
        RECT 265.200 214.200 266.000 215.000 ;
        RECT 289.200 217.600 290.000 218.400 ;
        RECT 276.400 211.600 277.200 212.400 ;
        RECT 247.600 203.600 248.400 204.400 ;
        RECT 258.800 206.800 259.600 207.600 ;
        RECT 262.000 206.200 262.800 207.000 ;
        RECT 257.200 204.200 258.000 205.000 ;
        RECT 258.800 204.200 259.600 205.000 ;
        RECT 260.400 204.200 261.200 205.000 ;
        RECT 265.200 206.200 266.000 207.000 ;
        RECT 268.400 206.200 269.200 207.000 ;
        RECT 270.000 204.200 270.800 205.000 ;
        RECT 271.600 204.200 272.400 205.000 ;
        RECT 292.400 215.600 293.200 216.400 ;
        RECT 308.400 215.600 309.200 216.400 ;
        RECT 310.000 214.200 310.800 215.000 ;
        RECT 318.000 210.000 318.800 210.800 ;
        RECT 292.400 203.600 293.200 204.400 ;
        RECT 303.600 206.800 304.400 207.600 ;
        RECT 306.800 206.200 307.600 207.000 ;
        RECT 302.000 204.200 302.800 205.000 ;
        RECT 303.600 204.200 304.400 205.000 ;
        RECT 305.200 204.200 306.000 205.000 ;
        RECT 310.000 206.200 310.800 207.000 ;
        RECT 313.200 206.200 314.000 207.000 ;
        RECT 343.600 217.600 344.400 218.400 ;
        RECT 314.800 204.200 315.600 205.000 ;
        RECT 316.400 204.200 317.200 205.000 ;
        RECT 332.400 213.600 333.200 214.400 ;
        RECT 345.200 217.600 346.000 218.400 ;
        RECT 361.200 213.600 362.000 214.400 ;
        RECT 366.000 213.600 366.800 214.400 ;
        RECT 388.400 217.600 389.200 218.400 ;
        RECT 370.800 213.600 371.600 214.400 ;
        RECT 350.000 212.200 350.800 213.000 ;
        RECT 358.000 211.800 358.800 212.600 ;
        RECT 362.800 210.200 363.600 211.000 ;
        RECT 382.000 213.600 382.800 214.400 ;
        RECT 383.600 211.600 384.400 212.400 ;
        RECT 394.800 213.600 395.600 214.400 ;
        RECT 396.400 213.600 397.200 214.400 ;
        RECT 404.400 213.600 405.200 214.400 ;
        RECT 433.200 217.600 434.000 218.400 ;
        RECT 388.400 209.600 389.200 210.400 ;
        RECT 394.800 209.600 395.600 210.400 ;
        RECT 412.400 211.600 413.200 212.400 ;
        RECT 401.200 203.600 402.000 204.400 ;
        RECT 434.800 213.600 435.600 214.400 ;
        RECT 430.000 211.600 430.800 212.400 ;
        RECT 436.400 211.600 437.200 212.400 ;
        RECT 447.600 213.600 448.400 214.400 ;
        RECT 481.200 217.600 482.000 218.400 ;
        RECT 462.000 213.600 462.800 214.400 ;
        RECT 441.200 211.600 442.000 212.400 ;
        RECT 442.800 211.600 443.600 212.400 ;
        RECT 414.000 203.600 414.800 204.400 ;
        RECT 444.400 207.600 445.200 208.400 ;
        RECT 476.400 211.600 477.200 212.400 ;
        RECT 497.200 215.600 498.000 216.400 ;
        RECT 498.800 214.200 499.600 215.000 ;
        RECT 506.800 211.600 507.600 212.400 ;
        RECT 468.400 203.600 469.200 204.400 ;
        RECT 478.000 209.600 478.800 210.400 ;
        RECT 481.200 203.600 482.000 204.400 ;
        RECT 492.400 206.800 493.200 207.600 ;
        RECT 495.600 206.200 496.400 207.000 ;
        RECT 490.800 204.200 491.600 205.000 ;
        RECT 492.400 204.200 493.200 205.000 ;
        RECT 494.000 204.200 494.800 205.000 ;
        RECT 498.800 206.200 499.600 207.000 ;
        RECT 502.000 206.200 502.800 207.000 ;
        RECT 522.800 213.000 523.600 213.800 ;
        RECT 532.400 212.600 533.200 213.400 ;
        RECT 518.000 211.600 518.800 212.400 ;
        RECT 524.400 208.800 525.200 209.600 ;
        RECT 529.200 207.600 530.000 208.400 ;
        RECT 503.600 204.200 504.400 205.000 ;
        RECT 505.200 204.200 506.000 205.000 ;
        RECT 526.000 206.200 526.800 207.000 ;
        RECT 522.800 204.200 523.600 205.000 ;
        RECT 524.400 204.200 525.200 205.000 ;
        RECT 529.200 206.200 530.000 207.000 ;
        RECT 532.400 206.200 533.200 207.000 ;
        RECT 534.000 204.200 534.800 205.000 ;
        RECT 535.600 204.200 536.400 205.000 ;
        RECT 537.200 204.200 538.000 205.000 ;
        RECT 1.200 187.600 2.000 188.400 ;
        RECT 9.200 187.600 10.000 188.400 ;
        RECT 31.600 195.600 32.400 196.400 ;
        RECT 36.400 193.600 37.200 194.400 ;
        RECT 42.800 197.600 43.600 198.400 ;
        RECT 41.200 193.600 42.000 194.400 ;
        RECT 4.400 183.600 5.200 184.400 ;
        RECT 7.600 183.600 8.400 184.400 ;
        RECT 14.000 185.600 14.800 186.400 ;
        RECT 33.200 191.600 34.000 192.400 ;
        RECT 22.000 185.600 22.800 186.400 ;
        RECT 20.400 183.600 21.200 184.400 ;
        RECT 26.800 185.600 27.600 186.400 ;
        RECT 44.400 191.600 45.200 192.400 ;
        RECT 42.800 189.600 43.600 190.400 ;
        RECT 46.000 185.600 46.800 186.400 ;
        RECT 49.200 187.600 50.000 188.400 ;
        RECT 57.200 197.600 58.000 198.400 ;
        RECT 55.600 193.600 56.400 194.400 ;
        RECT 58.800 191.600 59.600 192.400 ;
        RECT 57.200 189.600 58.000 190.400 ;
        RECT 47.600 183.600 48.400 184.400 ;
        RECT 52.400 183.600 53.200 184.400 ;
        RECT 84.400 195.000 85.200 195.800 ;
        RECT 81.200 193.600 82.000 194.400 ;
        RECT 98.800 197.600 99.600 198.400 ;
        RECT 86.000 192.400 86.800 193.200 ;
        RECT 90.800 189.600 91.600 190.400 ;
        RECT 74.800 188.200 75.600 189.000 ;
        RECT 84.400 188.600 85.200 189.400 ;
        RECT 79.600 187.600 80.400 188.400 ;
        RECT 74.800 184.200 75.600 185.000 ;
        RECT 76.400 184.200 77.200 185.000 ;
        RECT 78.000 184.200 78.800 185.000 ;
        RECT 81.200 184.200 82.000 185.000 ;
        RECT 84.400 184.200 85.200 185.000 ;
        RECT 86.000 184.200 86.800 185.000 ;
        RECT 87.600 184.200 88.400 185.000 ;
        RECT 89.200 184.200 90.000 185.000 ;
        RECT 114.800 194.400 115.600 195.200 ;
        RECT 118.000 195.000 118.800 195.800 ;
        RECT 113.200 192.400 114.000 193.200 ;
        RECT 129.200 191.200 130.000 192.000 ;
        RECT 103.600 183.600 104.400 184.400 ;
        RECT 122.800 187.600 123.600 188.400 ;
        RECT 119.600 185.600 120.400 186.400 ;
        RECT 113.200 184.200 114.000 185.000 ;
        RECT 114.800 184.200 115.600 185.000 ;
        RECT 116.400 184.200 117.200 185.000 ;
        RECT 118.000 184.200 118.800 185.000 ;
        RECT 121.200 184.200 122.000 185.000 ;
        RECT 124.400 184.200 125.200 185.000 ;
        RECT 126.000 184.200 126.800 185.000 ;
        RECT 127.600 184.200 128.400 185.000 ;
        RECT 161.200 195.000 162.000 195.800 ;
        RECT 158.000 193.600 158.800 194.400 ;
        RECT 175.600 197.600 176.400 198.400 ;
        RECT 162.800 192.400 163.600 193.200 ;
        RECT 151.600 188.200 152.400 189.000 ;
        RECT 161.200 188.600 162.000 189.400 ;
        RECT 156.400 187.600 157.200 188.400 ;
        RECT 151.600 184.200 152.400 185.000 ;
        RECT 153.200 184.200 154.000 185.000 ;
        RECT 154.800 184.200 155.600 185.000 ;
        RECT 158.000 184.200 158.800 185.000 ;
        RECT 161.200 184.200 162.000 185.000 ;
        RECT 162.800 184.200 163.600 185.000 ;
        RECT 164.400 184.200 165.200 185.000 ;
        RECT 166.000 184.200 166.800 185.000 ;
        RECT 183.600 197.600 184.400 198.400 ;
        RECT 194.800 194.400 195.600 195.200 ;
        RECT 198.000 195.000 198.800 195.800 ;
        RECT 193.200 192.400 194.000 193.200 ;
        RECT 191.600 189.600 192.400 190.400 ;
        RECT 178.800 183.600 179.600 184.400 ;
        RECT 202.800 187.600 203.600 188.400 ;
        RECT 199.600 185.600 200.400 186.400 ;
        RECT 193.200 184.200 194.000 185.000 ;
        RECT 194.800 184.200 195.600 185.000 ;
        RECT 196.400 184.200 197.200 185.000 ;
        RECT 198.000 184.200 198.800 185.000 ;
        RECT 201.200 184.200 202.000 185.000 ;
        RECT 204.400 184.200 205.200 185.000 ;
        RECT 206.000 184.200 206.800 185.000 ;
        RECT 207.600 184.200 208.400 185.000 ;
        RECT 223.600 197.600 224.400 198.400 ;
        RECT 222.000 193.600 222.800 194.400 ;
        RECT 223.600 189.600 224.400 190.400 ;
        RECT 218.800 185.600 219.600 186.400 ;
        RECT 230.000 187.600 230.800 188.400 ;
        RECT 228.400 185.600 229.200 186.400 ;
        RECT 233.200 183.600 234.000 184.400 ;
        RECT 238.000 185.600 238.800 186.400 ;
        RECT 249.200 189.600 250.000 190.400 ;
        RECT 279.600 194.400 280.400 195.200 ;
        RECT 282.800 195.000 283.600 195.800 ;
        RECT 278.000 192.400 278.800 193.200 ;
        RECT 244.400 185.600 245.200 186.400 ;
        RECT 268.200 189.600 269.000 190.400 ;
        RECT 287.600 187.600 288.400 188.400 ;
        RECT 284.400 185.600 285.200 186.400 ;
        RECT 278.000 184.200 278.800 185.000 ;
        RECT 279.600 184.200 280.400 185.000 ;
        RECT 281.200 184.200 282.000 185.000 ;
        RECT 282.800 184.200 283.600 185.000 ;
        RECT 286.000 184.200 286.800 185.000 ;
        RECT 289.200 184.200 290.000 185.000 ;
        RECT 290.800 184.200 291.600 185.000 ;
        RECT 292.400 184.200 293.200 185.000 ;
        RECT 314.800 194.400 315.600 195.200 ;
        RECT 318.000 195.000 318.800 195.800 ;
        RECT 313.200 192.400 314.000 193.200 ;
        RECT 332.400 191.600 333.200 192.400 ;
        RECT 303.600 183.600 304.400 184.400 ;
        RECT 322.800 187.600 323.600 188.400 ;
        RECT 319.600 185.600 320.400 186.400 ;
        RECT 313.200 184.200 314.000 185.000 ;
        RECT 314.800 184.200 315.600 185.000 ;
        RECT 316.400 184.200 317.200 185.000 ;
        RECT 318.000 184.200 318.800 185.000 ;
        RECT 321.200 184.200 322.000 185.000 ;
        RECT 324.400 184.200 325.200 185.000 ;
        RECT 326.000 184.200 326.800 185.000 ;
        RECT 327.600 184.200 328.400 185.000 ;
        RECT 342.000 189.600 342.800 190.400 ;
        RECT 364.400 195.000 365.200 195.800 ;
        RECT 361.200 193.600 362.000 194.400 ;
        RECT 366.000 192.400 366.800 193.200 ;
        RECT 353.200 191.200 354.000 192.000 ;
        RECT 393.200 197.600 394.000 198.400 ;
        RECT 391.600 193.600 392.400 194.400 ;
        RECT 337.200 185.600 338.000 186.400 ;
        RECT 345.200 187.600 346.000 188.400 ;
        RECT 354.800 188.200 355.600 189.000 ;
        RECT 364.400 188.600 365.200 189.400 ;
        RECT 359.600 187.600 360.400 188.400 ;
        RECT 379.000 189.600 379.800 190.400 ;
        RECT 354.800 184.200 355.600 185.000 ;
        RECT 356.400 184.200 357.200 185.000 ;
        RECT 358.000 184.200 358.800 185.000 ;
        RECT 361.200 184.200 362.000 185.000 ;
        RECT 364.400 184.200 365.200 185.000 ;
        RECT 366.000 184.200 366.800 185.000 ;
        RECT 367.600 184.200 368.400 185.000 ;
        RECT 369.200 184.200 370.000 185.000 ;
        RECT 388.400 191.600 389.200 192.400 ;
        RECT 385.200 189.600 386.000 190.400 ;
        RECT 386.800 187.600 387.600 188.400 ;
        RECT 407.600 197.600 408.400 198.400 ;
        RECT 401.200 189.600 402.000 190.400 ;
        RECT 398.000 187.600 398.800 188.400 ;
        RECT 404.400 183.600 405.200 184.400 ;
        RECT 410.800 197.600 411.600 198.400 ;
        RECT 412.400 193.600 413.200 194.400 ;
        RECT 415.600 193.600 416.400 194.400 ;
        RECT 409.200 191.600 410.000 192.400 ;
        RECT 417.200 185.600 418.000 186.400 ;
        RECT 447.600 197.600 448.400 198.400 ;
        RECT 446.000 193.600 446.800 194.400 ;
        RECT 434.800 189.600 435.600 190.400 ;
        RECT 436.400 189.600 437.200 190.400 ;
        RECT 465.200 197.600 466.000 198.400 ;
        RECT 470.000 197.600 470.800 198.400 ;
        RECT 447.600 189.600 448.400 190.400 ;
        RECT 433.200 185.600 434.000 186.400 ;
        RECT 439.600 183.600 440.400 184.400 ;
        RECT 460.400 191.600 461.200 192.400 ;
        RECT 458.800 189.600 459.600 190.400 ;
        RECT 481.200 194.400 482.000 195.200 ;
        RECT 484.400 195.000 485.200 195.800 ;
        RECT 508.400 197.600 509.200 198.400 ;
        RECT 479.600 192.400 480.400 193.200 ;
        RECT 465.200 189.600 466.000 190.400 ;
        RECT 454.000 183.600 454.800 184.400 ;
        RECT 466.800 187.600 467.600 188.400 ;
        RECT 478.000 189.600 478.800 190.400 ;
        RECT 489.200 187.600 490.000 188.400 ;
        RECT 486.000 185.600 486.800 186.400 ;
        RECT 505.200 189.600 506.000 190.400 ;
        RECT 508.400 189.600 509.200 190.400 ;
        RECT 511.600 189.600 512.400 190.400 ;
        RECT 513.200 189.600 514.000 190.400 ;
        RECT 479.600 184.200 480.400 185.000 ;
        RECT 481.200 184.200 482.000 185.000 ;
        RECT 482.800 184.200 483.600 185.000 ;
        RECT 484.400 184.200 485.200 185.000 ;
        RECT 487.600 184.200 488.400 185.000 ;
        RECT 490.800 184.200 491.600 185.000 ;
        RECT 492.400 184.200 493.200 185.000 ;
        RECT 494.000 184.200 494.800 185.000 ;
        RECT 527.600 189.600 528.400 190.400 ;
        RECT 521.200 186.200 522.000 187.000 ;
        RECT 542.000 189.600 542.800 190.400 ;
        RECT 550.000 187.600 550.800 188.400 ;
        RECT 538.800 183.600 539.600 184.400 ;
        RECT 20.400 173.600 21.200 174.400 ;
        RECT 12.400 171.600 13.200 172.400 ;
        RECT 14.000 171.600 14.800 172.400 ;
        RECT 15.600 169.600 16.400 170.400 ;
        RECT 22.000 175.600 22.800 176.400 ;
        RECT 36.400 177.600 37.200 178.400 ;
        RECT 49.200 177.600 50.000 178.400 ;
        RECT 52.400 177.600 53.200 178.400 ;
        RECT 57.200 177.600 58.000 178.400 ;
        RECT 44.400 173.600 45.200 174.400 ;
        RECT 28.400 171.600 29.200 172.400 ;
        RECT 28.400 163.600 29.200 164.400 ;
        RECT 49.200 169.600 50.000 170.400 ;
        RECT 73.200 175.600 74.000 176.400 ;
        RECT 74.800 174.200 75.600 175.000 ;
        RECT 86.000 171.600 86.800 172.400 ;
        RECT 68.400 166.800 69.200 167.600 ;
        RECT 71.600 166.200 72.400 167.000 ;
        RECT 66.800 164.200 67.600 165.000 ;
        RECT 68.400 164.200 69.200 165.000 ;
        RECT 70.000 164.200 70.800 165.000 ;
        RECT 74.800 166.200 75.600 167.000 ;
        RECT 78.000 166.200 78.800 167.000 ;
        RECT 97.200 171.600 98.000 172.400 ;
        RECT 79.600 164.200 80.400 165.000 ;
        RECT 81.200 164.200 82.000 165.000 ;
        RECT 95.600 169.600 96.400 170.400 ;
        RECT 106.800 173.600 107.600 174.400 ;
        RECT 134.000 175.600 134.800 176.400 ;
        RECT 135.600 174.200 136.400 175.000 ;
        RECT 118.000 163.600 118.800 164.400 ;
        RECT 129.200 166.800 130.000 167.600 ;
        RECT 132.400 166.200 133.200 167.000 ;
        RECT 127.600 164.200 128.400 165.000 ;
        RECT 129.200 164.200 130.000 165.000 ;
        RECT 130.800 164.200 131.600 165.000 ;
        RECT 135.600 166.200 136.400 167.000 ;
        RECT 138.800 166.200 139.600 167.000 ;
        RECT 159.600 173.000 160.400 173.800 ;
        RECT 169.200 172.600 170.000 173.400 ;
        RECT 153.200 171.600 154.000 172.400 ;
        RECT 175.600 171.600 176.400 172.400 ;
        RECT 161.200 168.800 162.000 169.600 ;
        RECT 166.000 167.600 166.800 168.400 ;
        RECT 140.400 164.200 141.200 165.000 ;
        RECT 142.000 164.200 142.800 165.000 ;
        RECT 162.800 166.200 163.600 167.000 ;
        RECT 159.600 164.200 160.400 165.000 ;
        RECT 161.200 164.200 162.000 165.000 ;
        RECT 166.000 166.200 166.800 167.000 ;
        RECT 169.200 166.200 170.000 167.000 ;
        RECT 170.800 164.200 171.600 165.000 ;
        RECT 172.400 164.200 173.200 165.000 ;
        RECT 174.000 164.200 174.800 165.000 ;
        RECT 183.600 163.600 184.400 164.400 ;
        RECT 190.000 169.600 190.800 170.400 ;
        RECT 196.400 171.600 197.200 172.400 ;
        RECT 218.800 175.600 219.600 176.400 ;
        RECT 220.400 174.200 221.200 175.000 ;
        RECT 210.800 171.600 211.600 172.400 ;
        RECT 222.000 171.600 222.800 172.400 ;
        RECT 202.800 163.600 203.600 164.400 ;
        RECT 214.000 166.800 214.800 167.600 ;
        RECT 217.200 166.200 218.000 167.000 ;
        RECT 212.400 164.200 213.200 165.000 ;
        RECT 214.000 164.200 214.800 165.000 ;
        RECT 215.600 164.200 216.400 165.000 ;
        RECT 220.400 166.200 221.200 167.000 ;
        RECT 223.600 166.200 224.400 167.000 ;
        RECT 254.000 177.600 254.800 178.400 ;
        RECT 258.800 177.600 259.600 178.400 ;
        RECT 241.200 171.600 242.000 172.400 ;
        RECT 225.200 164.200 226.000 165.000 ;
        RECT 226.800 164.200 227.600 165.000 ;
        RECT 252.400 169.600 253.200 170.400 ;
        RECT 271.600 177.600 272.400 178.400 ;
        RECT 260.400 173.600 261.200 174.400 ;
        RECT 265.200 173.600 266.000 174.400 ;
        RECT 262.000 171.600 262.800 172.400 ;
        RECT 266.800 171.600 267.600 172.400 ;
        RECT 273.200 173.600 274.000 174.400 ;
        RECT 286.000 173.600 286.800 174.400 ;
        RECT 287.600 169.600 288.400 170.400 ;
        RECT 292.400 171.600 293.200 172.400 ;
        RECT 311.600 175.600 312.400 176.400 ;
        RECT 313.200 174.200 314.000 175.000 ;
        RECT 321.200 171.600 322.000 172.400 ;
        RECT 324.400 171.600 325.200 172.400 ;
        RECT 306.800 166.800 307.600 167.600 ;
        RECT 310.000 166.200 310.800 167.000 ;
        RECT 305.200 164.200 306.000 165.000 ;
        RECT 306.800 164.200 307.600 165.000 ;
        RECT 308.400 164.200 309.200 165.000 ;
        RECT 313.200 166.200 314.000 167.000 ;
        RECT 316.400 166.200 317.200 167.000 ;
        RECT 329.200 169.600 330.000 170.400 ;
        RECT 318.000 164.200 318.800 165.000 ;
        RECT 319.600 164.200 320.400 165.000 ;
        RECT 342.000 177.600 342.800 178.400 ;
        RECT 353.200 175.600 354.000 176.400 ;
        RECT 330.800 163.600 331.600 164.400 ;
        RECT 353.200 163.600 354.000 164.400 ;
        RECT 362.800 177.600 363.600 178.400 ;
        RECT 372.400 173.000 373.200 173.800 ;
        RECT 362.800 169.600 363.600 170.400 ;
        RECT 382.000 172.600 382.800 173.400 ;
        RECT 388.400 171.600 389.200 172.400 ;
        RECT 374.000 168.800 374.800 169.600 ;
        RECT 378.800 167.600 379.600 168.400 ;
        RECT 375.600 166.200 376.400 167.000 ;
        RECT 372.400 164.200 373.200 165.000 ;
        RECT 374.000 164.200 374.800 165.000 ;
        RECT 378.800 166.200 379.600 167.000 ;
        RECT 382.000 166.200 382.800 167.000 ;
        RECT 383.600 164.200 384.400 165.000 ;
        RECT 385.200 164.200 386.000 165.000 ;
        RECT 386.800 164.200 387.600 165.000 ;
        RECT 402.800 171.600 403.600 172.400 ;
        RECT 406.000 171.600 406.800 172.400 ;
        RECT 434.800 175.600 435.600 176.400 ;
        RECT 436.400 174.200 437.200 175.000 ;
        RECT 447.600 171.600 448.400 172.400 ;
        RECT 396.400 163.600 397.200 164.400 ;
        RECT 402.800 163.600 403.600 164.400 ;
        RECT 407.600 163.600 408.400 164.400 ;
        RECT 430.000 166.800 430.800 167.600 ;
        RECT 433.200 166.200 434.000 167.000 ;
        RECT 428.400 164.200 429.200 165.000 ;
        RECT 430.000 164.200 430.800 165.000 ;
        RECT 431.600 164.200 432.400 165.000 ;
        RECT 436.400 166.200 437.200 167.000 ;
        RECT 439.600 166.200 440.400 167.000 ;
        RECT 452.400 171.600 453.200 172.400 ;
        RECT 474.800 177.600 475.600 178.400 ;
        RECT 441.200 164.200 442.000 165.000 ;
        RECT 442.800 164.200 443.600 165.000 ;
        RECT 454.000 163.600 454.800 164.400 ;
        RECT 470.000 171.600 470.800 172.400 ;
        RECT 487.600 177.600 488.400 178.400 ;
        RECT 479.600 167.600 480.400 168.400 ;
        RECT 466.800 165.600 467.600 166.400 ;
        RECT 511.600 177.600 512.400 178.400 ;
        RECT 514.800 177.600 515.600 178.400 ;
        RECT 489.200 167.600 490.000 168.400 ;
        RECT 487.600 163.600 488.400 164.400 ;
        RECT 495.600 163.600 496.400 164.400 ;
        RECT 505.200 173.600 506.000 174.400 ;
        RECT 506.800 171.600 507.600 172.400 ;
        RECT 502.000 163.600 502.800 164.400 ;
        RECT 530.800 175.600 531.600 176.400 ;
        RECT 532.400 174.200 533.200 175.000 ;
        RECT 511.600 169.600 512.400 170.400 ;
        RECT 526.000 166.800 526.800 167.600 ;
        RECT 529.200 166.200 530.000 167.000 ;
        RECT 524.400 164.200 525.200 165.000 ;
        RECT 526.000 164.200 526.800 165.000 ;
        RECT 527.600 164.200 528.400 165.000 ;
        RECT 532.400 166.200 533.200 167.000 ;
        RECT 535.600 166.200 536.400 167.000 ;
        RECT 537.200 164.200 538.000 165.000 ;
        RECT 538.800 164.200 539.600 165.000 ;
        RECT 6.000 151.600 6.800 152.400 ;
        RECT 4.400 149.600 5.200 150.400 ;
        RECT 18.800 149.600 19.600 150.400 ;
        RECT 20.400 147.600 21.200 148.400 ;
        RECT 36.400 153.600 37.200 154.400 ;
        RECT 25.200 145.600 26.000 146.400 ;
        RECT 20.400 143.600 21.200 144.400 ;
        RECT 28.400 145.600 29.200 146.400 ;
        RECT 33.200 145.600 34.000 146.400 ;
        RECT 42.800 157.600 43.600 158.400 ;
        RECT 41.200 147.600 42.000 148.400 ;
        RECT 39.600 145.600 40.400 146.400 ;
        RECT 49.200 145.600 50.000 146.400 ;
        RECT 82.800 154.400 83.600 155.200 ;
        RECT 86.000 155.000 86.800 155.800 ;
        RECT 81.200 152.400 82.000 153.200 ;
        RECT 79.600 149.600 80.400 150.400 ;
        RECT 71.600 143.600 72.400 144.400 ;
        RECT 90.800 147.600 91.600 148.400 ;
        RECT 87.600 145.600 88.400 146.400 ;
        RECT 81.200 144.200 82.000 145.000 ;
        RECT 82.800 144.200 83.600 145.000 ;
        RECT 84.400 144.200 85.200 145.000 ;
        RECT 86.000 144.200 86.800 145.000 ;
        RECT 89.200 144.200 90.000 145.000 ;
        RECT 92.400 144.200 93.200 145.000 ;
        RECT 94.000 144.200 94.800 145.000 ;
        RECT 95.600 144.200 96.400 145.000 ;
        RECT 121.200 155.600 122.000 156.400 ;
        RECT 114.800 149.600 115.600 150.400 ;
        RECT 116.400 147.600 117.200 148.400 ;
        RECT 111.600 143.600 112.400 144.400 ;
        RECT 119.600 145.600 120.400 146.400 ;
        RECT 135.600 149.600 136.400 150.400 ;
        RECT 129.200 146.200 130.000 147.000 ;
        RECT 146.800 143.600 147.600 144.400 ;
        RECT 166.000 155.000 166.800 155.800 ;
        RECT 162.800 153.600 163.600 154.400 ;
        RECT 167.600 152.400 168.400 153.200 ;
        RECT 172.400 149.600 173.200 150.400 ;
        RECT 156.400 148.200 157.200 149.000 ;
        RECT 166.000 148.600 166.800 149.400 ;
        RECT 161.200 147.600 162.000 148.400 ;
        RECT 185.200 149.600 186.000 150.400 ;
        RECT 156.400 144.200 157.200 145.000 ;
        RECT 158.000 144.200 158.800 145.000 ;
        RECT 159.600 144.200 160.400 145.000 ;
        RECT 162.800 144.200 163.600 145.000 ;
        RECT 166.000 144.200 166.800 145.000 ;
        RECT 167.600 144.200 168.400 145.000 ;
        RECT 169.200 144.200 170.000 145.000 ;
        RECT 170.800 144.200 171.600 145.000 ;
        RECT 180.400 143.600 181.200 144.400 ;
        RECT 201.200 145.600 202.000 146.400 ;
        RECT 207.600 145.600 208.400 146.400 ;
        RECT 218.800 149.600 219.600 150.400 ;
        RECT 239.600 155.000 240.400 155.800 ;
        RECT 236.400 153.600 237.200 154.400 ;
        RECT 241.200 152.400 242.000 153.200 ;
        RECT 258.800 157.600 259.600 158.400 ;
        RECT 230.000 148.200 230.800 149.000 ;
        RECT 239.600 148.600 240.400 149.400 ;
        RECT 234.800 147.600 235.600 148.400 ;
        RECT 230.000 144.200 230.800 145.000 ;
        RECT 231.600 144.200 232.400 145.000 ;
        RECT 233.200 144.200 234.000 145.000 ;
        RECT 236.400 144.200 237.200 145.000 ;
        RECT 239.600 144.200 240.400 145.000 ;
        RECT 241.200 144.200 242.000 145.000 ;
        RECT 242.800 144.200 243.600 145.000 ;
        RECT 244.400 144.200 245.200 145.000 ;
        RECT 270.000 157.600 270.800 158.400 ;
        RECT 271.600 153.600 272.400 154.400 ;
        RECT 268.400 151.600 269.200 152.400 ;
        RECT 286.000 157.600 286.800 158.400 ;
        RECT 260.400 147.600 261.200 148.400 ;
        RECT 254.000 143.600 254.800 144.400 ;
        RECT 306.800 154.400 307.600 155.200 ;
        RECT 310.000 155.000 310.800 155.800 ;
        RECT 305.200 152.400 306.000 153.200 ;
        RECT 321.200 151.200 322.000 152.000 ;
        RECT 290.800 149.600 291.600 150.400 ;
        RECT 295.400 149.600 296.200 150.400 ;
        RECT 314.800 147.600 315.600 148.400 ;
        RECT 311.600 145.600 312.400 146.400 ;
        RECT 332.400 149.600 333.200 150.400 ;
        RECT 305.200 144.200 306.000 145.000 ;
        RECT 306.800 144.200 307.600 145.000 ;
        RECT 308.400 144.200 309.200 145.000 ;
        RECT 310.000 144.200 310.800 145.000 ;
        RECT 313.200 144.200 314.000 145.000 ;
        RECT 316.400 144.200 317.200 145.000 ;
        RECT 318.000 144.200 318.800 145.000 ;
        RECT 319.600 144.200 320.400 145.000 ;
        RECT 354.800 157.600 355.600 158.400 ;
        RECT 361.200 149.600 362.000 150.400 ;
        RECT 337.200 145.600 338.000 146.400 ;
        RECT 343.600 147.600 344.400 148.400 ;
        RECT 350.000 147.600 350.800 148.400 ;
        RECT 356.400 147.600 357.200 148.400 ;
        RECT 383.600 149.600 384.400 150.400 ;
        RECT 385.200 149.600 386.000 150.400 ;
        RECT 386.800 149.600 387.600 150.400 ;
        RECT 372.400 143.600 373.200 144.400 ;
        RECT 398.000 153.600 398.800 154.400 ;
        RECT 404.400 153.600 405.200 154.400 ;
        RECT 388.400 145.600 389.200 146.400 ;
        RECT 401.200 151.600 402.000 152.400 ;
        RECT 399.600 149.600 400.400 150.400 ;
        RECT 407.600 151.600 408.400 152.400 ;
        RECT 406.000 149.600 406.800 150.400 ;
        RECT 412.400 149.600 413.200 150.400 ;
        RECT 418.800 149.600 419.600 150.400 ;
        RECT 420.400 149.600 421.200 150.400 ;
        RECT 462.000 157.600 462.800 158.400 ;
        RECT 455.600 153.600 456.400 154.400 ;
        RECT 463.600 153.600 464.400 154.400 ;
        RECT 404.400 143.600 405.200 144.400 ;
        RECT 415.600 145.600 416.400 146.400 ;
        RECT 417.200 143.600 418.000 144.400 ;
        RECT 436.400 147.600 437.200 148.400 ;
        RECT 434.800 146.200 435.600 147.000 ;
        RECT 452.400 147.600 453.200 148.400 ;
        RECT 457.200 149.600 458.000 150.400 ;
        RECT 486.000 149.600 486.800 150.400 ;
        RECT 487.600 149.600 488.400 150.400 ;
        RECT 497.200 157.600 498.000 158.400 ;
        RECT 494.000 149.600 494.800 150.400 ;
        RECT 497.200 149.600 498.000 150.400 ;
        RECT 510.000 157.600 510.800 158.400 ;
        RECT 489.200 145.600 490.000 146.400 ;
        RECT 490.800 145.600 491.600 146.400 ;
        RECT 498.800 147.600 499.600 148.400 ;
        RECT 506.800 149.600 507.600 150.400 ;
        RECT 508.400 149.600 509.200 150.400 ;
        RECT 511.600 145.600 512.400 146.400 ;
        RECT 521.200 157.600 522.000 158.400 ;
        RECT 516.400 149.600 517.200 150.400 ;
        RECT 518.000 149.600 518.800 150.400 ;
        RECT 543.600 157.600 544.400 158.400 ;
        RECT 514.800 145.600 515.600 146.400 ;
        RECT 526.000 146.200 526.800 147.000 ;
        RECT 545.200 149.600 546.000 150.400 ;
        RECT 6.000 133.600 6.800 134.400 ;
        RECT 1.200 123.600 2.000 124.400 ;
        RECT 20.400 133.600 21.200 134.400 ;
        RECT 41.200 133.600 42.000 134.400 ;
        RECT 50.800 137.600 51.600 138.400 ;
        RECT 9.200 131.600 10.000 132.400 ;
        RECT 7.600 129.600 8.400 130.400 ;
        RECT 15.600 131.600 16.400 132.400 ;
        RECT 26.800 131.600 27.600 132.400 ;
        RECT 22.000 129.600 22.800 130.400 ;
        RECT 33.200 131.600 34.000 132.400 ;
        RECT 46.000 131.600 46.800 132.400 ;
        RECT 26.800 123.600 27.600 124.400 ;
        RECT 33.200 125.600 34.000 126.400 ;
        RECT 41.200 129.600 42.000 130.400 ;
        RECT 66.800 135.600 67.600 136.400 ;
        RECT 68.400 134.200 69.200 135.000 ;
        RECT 70.000 131.600 70.800 132.400 ;
        RECT 79.600 131.600 80.400 132.400 ;
        RECT 46.000 123.600 46.800 124.400 ;
        RECT 62.000 126.800 62.800 127.600 ;
        RECT 65.200 126.200 66.000 127.000 ;
        RECT 60.400 124.200 61.200 125.000 ;
        RECT 62.000 124.200 62.800 125.000 ;
        RECT 63.600 124.200 64.400 125.000 ;
        RECT 68.400 126.200 69.200 127.000 ;
        RECT 71.600 126.200 72.400 127.000 ;
        RECT 89.200 137.600 90.000 138.400 ;
        RECT 94.000 133.600 94.800 134.400 ;
        RECT 86.000 129.600 86.800 130.400 ;
        RECT 73.200 124.200 74.000 125.000 ;
        RECT 74.800 124.200 75.600 125.000 ;
        RECT 106.800 133.000 107.600 133.800 ;
        RECT 97.200 131.600 98.000 132.400 ;
        RECT 116.400 132.600 117.200 133.400 ;
        RECT 100.400 131.600 101.200 132.400 ;
        RECT 122.800 131.600 123.600 132.400 ;
        RECT 108.400 128.800 109.200 129.600 ;
        RECT 113.200 127.600 114.000 128.400 ;
        RECT 110.000 126.200 110.800 127.000 ;
        RECT 106.800 124.200 107.600 125.000 ;
        RECT 108.400 124.200 109.200 125.000 ;
        RECT 113.200 126.200 114.000 127.000 ;
        RECT 116.400 126.200 117.200 127.000 ;
        RECT 118.000 124.200 118.800 125.000 ;
        RECT 119.600 124.200 120.400 125.000 ;
        RECT 121.200 124.200 122.000 125.000 ;
        RECT 130.800 123.600 131.600 124.400 ;
        RECT 154.800 137.600 155.600 138.400 ;
        RECT 172.400 137.600 173.200 138.400 ;
        RECT 175.600 137.600 176.400 138.400 ;
        RECT 161.200 133.600 162.000 134.400 ;
        RECT 162.800 131.600 163.600 132.400 ;
        RECT 156.400 129.600 157.200 130.400 ;
        RECT 172.400 129.600 173.200 130.400 ;
        RECT 183.400 131.600 184.200 132.400 ;
        RECT 199.600 135.600 200.400 136.400 ;
        RECT 201.200 134.200 202.000 135.000 ;
        RECT 210.800 131.600 211.600 132.400 ;
        RECT 194.800 126.800 195.600 127.600 ;
        RECT 198.000 126.200 198.800 127.000 ;
        RECT 193.200 124.200 194.000 125.000 ;
        RECT 194.800 124.200 195.600 125.000 ;
        RECT 196.400 124.200 197.200 125.000 ;
        RECT 201.200 126.200 202.000 127.000 ;
        RECT 204.400 126.200 205.200 127.000 ;
        RECT 231.600 131.600 232.400 132.400 ;
        RECT 238.000 131.600 238.800 132.400 ;
        RECT 206.000 124.200 206.800 125.000 ;
        RECT 207.600 124.200 208.400 125.000 ;
        RECT 233.200 129.600 234.000 130.400 ;
        RECT 246.000 135.600 246.800 136.400 ;
        RECT 273.200 135.600 274.000 136.400 ;
        RECT 249.200 131.600 250.000 132.400 ;
        RECT 257.200 131.600 258.000 132.400 ;
        RECT 289.200 135.600 290.000 136.400 ;
        RECT 290.800 134.200 291.600 135.000 ;
        RECT 246.000 123.600 246.800 124.400 ;
        RECT 250.800 123.600 251.600 124.400 ;
        RECT 263.600 129.600 264.400 130.400 ;
        RECT 284.400 126.800 285.200 127.600 ;
        RECT 287.600 126.200 288.400 127.000 ;
        RECT 282.800 124.200 283.600 125.000 ;
        RECT 284.400 124.200 285.200 125.000 ;
        RECT 286.000 124.200 286.800 125.000 ;
        RECT 290.800 126.200 291.600 127.000 ;
        RECT 294.000 126.200 294.800 127.000 ;
        RECT 295.600 124.200 296.400 125.000 ;
        RECT 297.200 124.200 298.000 125.000 ;
        RECT 330.800 133.000 331.600 133.800 ;
        RECT 340.400 132.600 341.200 133.400 ;
        RECT 326.000 131.600 326.800 132.400 ;
        RECT 332.400 128.800 333.200 129.600 ;
        RECT 337.200 127.600 338.000 128.400 ;
        RECT 334.000 126.200 334.800 127.000 ;
        RECT 330.800 124.200 331.600 125.000 ;
        RECT 332.400 124.200 333.200 125.000 ;
        RECT 337.200 126.200 338.000 127.000 ;
        RECT 340.400 126.200 341.200 127.000 ;
        RECT 342.000 124.200 342.800 125.000 ;
        RECT 343.600 124.200 344.400 125.000 ;
        RECT 345.200 124.200 346.000 125.000 ;
        RECT 362.800 135.600 363.600 136.400 ;
        RECT 364.400 133.600 365.200 134.400 ;
        RECT 374.000 133.600 374.800 134.400 ;
        RECT 385.200 133.600 386.000 134.400 ;
        RECT 396.400 137.600 397.200 138.400 ;
        RECT 382.000 131.600 382.800 132.400 ;
        RECT 390.000 131.600 390.800 132.400 ;
        RECT 377.200 123.600 378.000 124.400 ;
        RECT 388.400 127.600 389.200 128.400 ;
        RECT 412.400 135.600 413.200 136.400 ;
        RECT 414.000 134.200 414.800 135.000 ;
        RECT 425.200 131.600 426.000 132.400 ;
        RECT 391.600 123.600 392.400 124.400 ;
        RECT 407.600 126.800 408.400 127.600 ;
        RECT 410.800 126.200 411.600 127.000 ;
        RECT 406.000 124.200 406.800 125.000 ;
        RECT 407.600 124.200 408.400 125.000 ;
        RECT 409.200 124.200 410.000 125.000 ;
        RECT 414.000 126.200 414.800 127.000 ;
        RECT 417.200 126.200 418.000 127.000 ;
        RECT 442.800 133.600 443.600 134.400 ;
        RECT 439.600 131.600 440.400 132.400 ;
        RECT 418.800 124.200 419.600 125.000 ;
        RECT 420.400 124.200 421.200 125.000 ;
        RECT 457.200 123.600 458.000 124.400 ;
        RECT 473.200 133.000 474.000 133.800 ;
        RECT 482.800 132.600 483.600 133.400 ;
        RECT 497.200 137.600 498.000 138.400 ;
        RECT 470.000 131.600 470.800 132.400 ;
        RECT 474.800 128.800 475.600 129.600 ;
        RECT 479.600 127.600 480.400 128.400 ;
        RECT 476.400 126.200 477.200 127.000 ;
        RECT 473.200 124.200 474.000 125.000 ;
        RECT 474.800 124.200 475.600 125.000 ;
        RECT 479.600 126.200 480.400 127.000 ;
        RECT 482.800 126.200 483.600 127.000 ;
        RECT 484.400 124.200 485.200 125.000 ;
        RECT 486.000 124.200 486.800 125.000 ;
        RECT 487.600 124.200 488.400 125.000 ;
        RECT 506.800 131.600 507.600 132.400 ;
        RECT 532.400 135.600 533.200 136.400 ;
        RECT 534.000 134.200 534.800 135.000 ;
        RECT 543.600 131.600 544.400 132.400 ;
        RECT 513.200 129.600 514.000 130.400 ;
        RECT 505.200 123.600 506.000 124.400 ;
        RECT 527.600 126.800 528.400 127.600 ;
        RECT 530.800 126.200 531.600 127.000 ;
        RECT 526.000 124.200 526.800 125.000 ;
        RECT 527.600 124.200 528.400 125.000 ;
        RECT 529.200 124.200 530.000 125.000 ;
        RECT 534.000 126.200 534.800 127.000 ;
        RECT 537.200 126.200 538.000 127.000 ;
        RECT 538.800 124.200 539.600 125.000 ;
        RECT 540.400 124.200 541.200 125.000 ;
        RECT 4.400 117.600 5.200 118.400 ;
        RECT 9.200 117.600 10.000 118.400 ;
        RECT 4.400 109.600 5.200 110.400 ;
        RECT 7.600 107.600 8.400 108.400 ;
        RECT 22.000 117.600 22.800 118.400 ;
        RECT 30.000 117.600 30.800 118.400 ;
        RECT 14.000 113.600 14.800 114.400 ;
        RECT 20.400 113.600 21.200 114.400 ;
        RECT 28.400 113.600 29.200 114.400 ;
        RECT 17.200 111.600 18.000 112.400 ;
        RECT 15.600 109.600 16.400 110.400 ;
        RECT 23.600 111.600 24.400 112.400 ;
        RECT 25.200 111.600 26.000 112.400 ;
        RECT 22.000 109.600 22.800 110.400 ;
        RECT 33.200 107.600 34.000 108.400 ;
        RECT 36.400 107.600 37.200 108.400 ;
        RECT 55.600 114.400 56.400 115.200 ;
        RECT 58.800 115.000 59.600 115.800 ;
        RECT 54.000 112.400 54.800 113.200 ;
        RECT 41.200 107.600 42.000 108.400 ;
        RECT 39.600 103.600 40.400 104.400 ;
        RECT 44.400 103.600 45.200 104.400 ;
        RECT 63.600 107.600 64.400 108.400 ;
        RECT 60.400 105.600 61.200 106.400 ;
        RECT 79.600 109.600 80.400 110.400 ;
        RECT 102.000 115.000 102.800 115.800 ;
        RECT 98.800 113.600 99.600 114.400 ;
        RECT 116.400 117.600 117.200 118.400 ;
        RECT 103.600 112.400 104.400 113.200 ;
        RECT 119.600 117.600 120.400 118.400 ;
        RECT 108.400 109.600 109.200 110.400 ;
        RECT 54.000 104.200 54.800 105.000 ;
        RECT 55.600 104.200 56.400 105.000 ;
        RECT 57.200 104.200 58.000 105.000 ;
        RECT 58.800 104.200 59.600 105.000 ;
        RECT 62.000 104.200 62.800 105.000 ;
        RECT 65.200 104.200 66.000 105.000 ;
        RECT 66.800 104.200 67.600 105.000 ;
        RECT 68.400 104.200 69.200 105.000 ;
        RECT 92.400 108.200 93.200 109.000 ;
        RECT 102.000 108.600 102.800 109.400 ;
        RECT 82.800 103.600 83.600 104.400 ;
        RECT 97.200 107.600 98.000 108.400 ;
        RECT 92.400 104.200 93.200 105.000 ;
        RECT 94.000 104.200 94.800 105.000 ;
        RECT 95.600 104.200 96.400 105.000 ;
        RECT 98.800 104.200 99.600 105.000 ;
        RECT 102.000 104.200 102.800 105.000 ;
        RECT 103.600 104.200 104.400 105.000 ;
        RECT 105.200 104.200 106.000 105.000 ;
        RECT 106.800 104.200 107.600 105.000 ;
        RECT 132.400 105.600 133.200 106.400 ;
        RECT 140.400 105.600 141.200 106.400 ;
        RECT 150.000 109.600 150.800 110.400 ;
        RECT 159.600 117.600 160.400 118.400 ;
        RECT 135.600 103.600 136.400 104.400 ;
        RECT 151.600 107.600 152.400 108.400 ;
        RECT 146.800 105.600 147.600 106.400 ;
        RECT 167.600 109.600 168.400 110.400 ;
        RECT 161.200 105.600 162.000 106.400 ;
        RECT 175.600 107.600 176.400 108.400 ;
        RECT 174.000 105.600 174.800 106.400 ;
        RECT 198.000 115.000 198.800 115.800 ;
        RECT 194.800 113.600 195.600 114.400 ;
        RECT 199.600 112.400 200.400 113.200 ;
        RECT 212.400 113.600 213.200 114.400 ;
        RECT 188.400 108.200 189.200 109.000 ;
        RECT 198.000 108.600 198.800 109.400 ;
        RECT 193.200 107.600 194.000 108.400 ;
        RECT 188.400 104.200 189.200 105.000 ;
        RECT 190.000 104.200 190.800 105.000 ;
        RECT 191.600 104.200 192.400 105.000 ;
        RECT 194.800 104.200 195.600 105.000 ;
        RECT 198.000 104.200 198.800 105.000 ;
        RECT 199.600 104.200 200.400 105.000 ;
        RECT 201.200 104.200 202.000 105.000 ;
        RECT 202.800 104.200 203.600 105.000 ;
        RECT 225.200 107.600 226.000 108.400 ;
        RECT 233.200 105.600 234.000 106.400 ;
        RECT 250.800 109.600 251.600 110.400 ;
        RECT 286.000 114.400 286.800 115.200 ;
        RECT 289.200 115.000 290.000 115.800 ;
        RECT 284.400 112.400 285.200 113.200 ;
        RECT 300.400 111.200 301.200 112.000 ;
        RECT 303.600 111.600 304.400 112.400 ;
        RECT 239.600 105.600 240.400 106.400 ;
        RECT 241.200 105.600 242.000 106.400 ;
        RECT 252.400 107.600 253.200 108.400 ;
        RECT 274.600 109.600 275.400 110.400 ;
        RECT 247.600 103.600 248.400 104.400 ;
        RECT 263.600 103.600 264.400 104.400 ;
        RECT 294.000 107.600 294.800 108.400 ;
        RECT 290.800 105.600 291.600 106.400 ;
        RECT 318.000 109.600 318.800 110.400 ;
        RECT 284.400 104.200 285.200 105.000 ;
        RECT 286.000 104.200 286.800 105.000 ;
        RECT 287.600 104.200 288.400 105.000 ;
        RECT 289.200 104.200 290.000 105.000 ;
        RECT 292.400 104.200 293.200 105.000 ;
        RECT 295.600 104.200 296.400 105.000 ;
        RECT 297.200 104.200 298.000 105.000 ;
        RECT 298.800 104.200 299.600 105.000 ;
        RECT 316.400 107.600 317.200 108.400 ;
        RECT 321.200 105.600 322.000 106.400 ;
        RECT 356.400 115.000 357.200 115.800 ;
        RECT 353.200 113.600 354.000 114.400 ;
        RECT 358.000 112.400 358.800 113.200 ;
        RECT 382.000 117.600 382.800 118.400 ;
        RECT 346.800 108.200 347.600 109.000 ;
        RECT 356.400 108.600 357.200 109.400 ;
        RECT 351.600 107.600 352.400 108.400 ;
        RECT 346.800 104.200 347.600 105.000 ;
        RECT 348.400 104.200 349.200 105.000 ;
        RECT 350.000 104.200 350.800 105.000 ;
        RECT 353.200 104.200 354.000 105.000 ;
        RECT 356.400 104.200 357.200 105.000 ;
        RECT 358.000 104.200 358.800 105.000 ;
        RECT 359.600 104.200 360.400 105.000 ;
        RECT 361.200 104.200 362.000 105.000 ;
        RECT 375.600 109.600 376.400 110.400 ;
        RECT 378.800 109.600 379.600 110.400 ;
        RECT 377.200 107.600 378.000 108.400 ;
        RECT 390.000 117.600 390.800 118.400 ;
        RECT 370.800 103.600 371.600 104.400 ;
        RECT 383.600 105.600 384.400 106.400 ;
        RECT 399.600 107.600 400.400 108.400 ;
        RECT 396.400 105.600 397.200 106.400 ;
        RECT 407.600 109.600 408.400 110.400 ;
        RECT 417.200 111.600 418.000 112.400 ;
        RECT 444.400 117.600 445.200 118.400 ;
        RECT 442.800 113.600 443.600 114.400 ;
        RECT 417.200 109.600 418.000 110.400 ;
        RECT 433.200 109.600 434.000 110.400 ;
        RECT 439.600 111.600 440.400 112.400 ;
        RECT 404.400 105.600 405.200 106.400 ;
        RECT 412.400 107.600 413.200 108.400 ;
        RECT 418.800 107.600 419.600 108.400 ;
        RECT 402.800 103.600 403.600 104.400 ;
        RECT 407.600 103.600 408.400 104.400 ;
        RECT 438.000 107.600 438.800 108.400 ;
        RECT 423.600 105.600 424.400 106.400 ;
        RECT 422.000 103.600 422.800 104.400 ;
        RECT 433.200 105.600 434.000 106.400 ;
        RECT 458.800 109.600 459.600 110.400 ;
        RECT 455.600 107.600 456.400 108.400 ;
        RECT 463.600 105.600 464.400 106.400 ;
        RECT 481.200 117.600 482.000 118.400 ;
        RECT 473.200 107.600 474.000 108.400 ;
        RECT 465.200 103.600 466.000 104.400 ;
        RECT 484.400 109.600 485.200 110.400 ;
        RECT 486.000 109.600 486.800 110.400 ;
        RECT 490.800 107.600 491.600 108.400 ;
        RECT 500.400 109.600 501.200 110.400 ;
        RECT 518.000 117.600 518.800 118.400 ;
        RECT 529.200 114.400 530.000 115.200 ;
        RECT 532.400 115.000 533.200 115.800 ;
        RECT 527.600 112.400 528.400 113.200 ;
        RECT 513.200 109.600 514.000 110.400 ;
        RECT 508.400 107.600 509.200 108.400 ;
        RECT 511.600 107.600 512.400 108.400 ;
        RECT 514.800 107.600 515.600 108.400 ;
        RECT 497.200 103.600 498.000 104.400 ;
        RECT 503.600 103.600 504.400 104.400 ;
        RECT 537.200 107.600 538.000 108.400 ;
        RECT 534.000 105.600 534.800 106.400 ;
        RECT 527.600 104.200 528.400 105.000 ;
        RECT 529.200 104.200 530.000 105.000 ;
        RECT 530.800 104.200 531.600 105.000 ;
        RECT 532.400 104.200 533.200 105.000 ;
        RECT 535.600 104.200 536.400 105.000 ;
        RECT 538.800 104.200 539.600 105.000 ;
        RECT 540.400 104.200 541.200 105.000 ;
        RECT 542.000 104.200 542.800 105.000 ;
        RECT 38.000 97.600 38.800 98.400 ;
        RECT 4.400 89.600 5.200 90.400 ;
        RECT 14.000 91.600 14.800 92.400 ;
        RECT 20.400 91.600 21.200 92.400 ;
        RECT 7.600 83.600 8.400 84.400 ;
        RECT 10.800 83.600 11.600 84.400 ;
        RECT 20.400 83.600 21.200 84.400 ;
        RECT 28.400 89.600 29.200 90.400 ;
        RECT 33.200 89.600 34.000 90.400 ;
        RECT 42.800 93.600 43.600 94.400 ;
        RECT 38.000 89.600 38.800 90.400 ;
        RECT 54.000 93.000 54.800 93.800 ;
        RECT 44.400 89.600 45.200 90.400 ;
        RECT 63.600 92.600 64.400 93.400 ;
        RECT 81.200 97.600 82.000 98.400 ;
        RECT 55.600 88.800 56.400 89.600 ;
        RECT 60.400 87.600 61.200 88.400 ;
        RECT 57.200 86.200 58.000 87.000 ;
        RECT 54.000 84.200 54.800 85.000 ;
        RECT 55.600 84.200 56.400 85.000 ;
        RECT 60.400 86.200 61.200 87.000 ;
        RECT 63.600 86.200 64.400 87.000 ;
        RECT 65.200 84.200 66.000 85.000 ;
        RECT 66.800 84.200 67.600 85.000 ;
        RECT 68.400 84.200 69.200 85.000 ;
        RECT 90.800 91.600 91.600 92.400 ;
        RECT 95.600 93.600 96.400 94.400 ;
        RECT 106.800 93.000 107.600 93.800 ;
        RECT 97.200 91.600 98.000 92.400 ;
        RECT 116.400 92.600 117.200 93.400 ;
        RECT 140.400 97.600 141.200 98.400 ;
        RECT 103.600 91.600 104.400 92.400 ;
        RECT 108.400 88.800 109.200 89.600 ;
        RECT 113.200 87.600 114.000 88.400 ;
        RECT 110.000 86.200 110.800 87.000 ;
        RECT 106.800 84.200 107.600 85.000 ;
        RECT 108.400 84.200 109.200 85.000 ;
        RECT 113.200 86.200 114.000 87.000 ;
        RECT 116.400 86.200 117.200 87.000 ;
        RECT 118.000 84.200 118.800 85.000 ;
        RECT 119.600 84.200 120.400 85.000 ;
        RECT 121.200 84.200 122.000 85.000 ;
        RECT 174.000 97.600 174.800 98.400 ;
        RECT 164.400 93.600 165.200 94.400 ;
        RECT 161.200 91.800 162.000 92.600 ;
        RECT 153.200 89.600 154.000 90.400 ;
        RECT 156.400 90.200 157.200 91.000 ;
        RECT 183.600 97.600 184.400 98.400 ;
        RECT 178.800 83.600 179.600 84.400 ;
        RECT 196.400 95.600 197.200 96.400 ;
        RECT 193.200 83.600 194.000 84.400 ;
        RECT 199.600 89.600 200.400 90.400 ;
        RECT 226.800 95.600 227.600 96.400 ;
        RECT 222.000 91.600 222.800 92.400 ;
        RECT 226.800 89.600 227.600 90.400 ;
        RECT 234.800 93.600 235.600 94.400 ;
        RECT 236.400 91.600 237.200 92.400 ;
        RECT 257.200 91.600 258.000 92.400 ;
        RECT 231.600 83.600 232.400 84.400 ;
        RECT 242.800 89.600 243.600 90.400 ;
        RECT 286.000 95.600 286.800 96.400 ;
        RECT 287.600 94.200 288.400 95.000 ;
        RECT 278.000 91.600 278.800 92.400 ;
        RECT 300.400 91.600 301.200 92.400 ;
        RECT 281.200 86.800 282.000 87.600 ;
        RECT 284.400 86.200 285.200 87.000 ;
        RECT 279.600 84.200 280.400 85.000 ;
        RECT 281.200 84.200 282.000 85.000 ;
        RECT 282.800 84.200 283.600 85.000 ;
        RECT 287.600 86.200 288.400 87.000 ;
        RECT 290.800 86.200 291.600 87.000 ;
        RECT 292.400 84.200 293.200 85.000 ;
        RECT 294.000 84.200 294.800 85.000 ;
        RECT 324.400 95.600 325.200 96.400 ;
        RECT 326.000 94.200 326.800 95.000 ;
        RECT 345.200 93.600 346.000 94.400 ;
        RECT 305.200 83.600 306.000 84.400 ;
        RECT 319.600 86.800 320.400 87.600 ;
        RECT 322.800 86.200 323.600 87.000 ;
        RECT 318.000 84.200 318.800 85.000 ;
        RECT 319.600 84.200 320.400 85.000 ;
        RECT 321.200 84.200 322.000 85.000 ;
        RECT 326.000 86.200 326.800 87.000 ;
        RECT 329.200 86.200 330.000 87.000 ;
        RECT 362.800 93.000 363.600 93.800 ;
        RECT 330.800 84.200 331.600 85.000 ;
        RECT 332.400 84.200 333.200 85.000 ;
        RECT 372.400 92.600 373.200 93.400 ;
        RECT 367.600 91.600 368.400 92.400 ;
        RECT 378.800 91.600 379.600 92.400 ;
        RECT 364.400 88.800 365.200 89.600 ;
        RECT 369.200 87.600 370.000 88.400 ;
        RECT 366.000 86.200 366.800 87.000 ;
        RECT 362.800 84.200 363.600 85.000 ;
        RECT 364.400 84.200 365.200 85.000 ;
        RECT 369.200 86.200 370.000 87.000 ;
        RECT 372.400 86.200 373.200 87.000 ;
        RECT 374.000 84.200 374.800 85.000 ;
        RECT 375.600 84.200 376.400 85.000 ;
        RECT 377.200 84.200 378.000 85.000 ;
        RECT 390.000 89.600 390.800 90.400 ;
        RECT 391.600 83.600 392.400 84.400 ;
        RECT 409.200 97.600 410.000 98.400 ;
        RECT 417.200 97.600 418.000 98.400 ;
        RECT 396.400 83.600 397.200 84.400 ;
        RECT 402.800 89.600 403.600 90.400 ;
        RECT 401.200 83.600 402.000 84.400 ;
        RECT 407.600 89.600 408.400 90.400 ;
        RECT 431.600 97.600 432.400 98.400 ;
        RECT 418.800 83.600 419.600 84.400 ;
        RECT 436.400 93.600 437.200 94.400 ;
        RECT 438.000 91.600 438.800 92.400 ;
        RECT 433.200 83.600 434.000 84.400 ;
        RECT 444.400 83.600 445.200 84.400 ;
        RECT 454.000 97.600 454.800 98.400 ;
        RECT 468.400 97.600 469.200 98.400 ;
        RECT 482.800 97.600 483.600 98.400 ;
        RECT 449.200 89.600 450.000 90.400 ;
        RECT 447.600 83.600 448.400 84.400 ;
        RECT 466.800 93.600 467.600 94.400 ;
        RECT 471.600 91.600 472.400 92.400 ;
        RECT 473.200 91.600 474.000 92.400 ;
        RECT 479.600 91.600 480.400 92.400 ;
        RECT 498.800 95.600 499.600 96.400 ;
        RECT 500.400 94.200 501.200 95.000 ;
        RECT 518.000 97.600 518.800 98.400 ;
        RECT 511.600 91.600 512.400 92.400 ;
        RECT 454.000 83.600 454.800 84.400 ;
        RECT 460.400 83.600 461.200 84.400 ;
        RECT 494.000 86.800 494.800 87.600 ;
        RECT 497.200 86.200 498.000 87.000 ;
        RECT 492.400 84.200 493.200 85.000 ;
        RECT 494.000 84.200 494.800 85.000 ;
        RECT 495.600 84.200 496.400 85.000 ;
        RECT 500.400 86.200 501.200 87.000 ;
        RECT 503.600 86.200 504.400 87.000 ;
        RECT 534.000 95.600 534.800 96.400 ;
        RECT 535.600 94.200 536.400 95.000 ;
        RECT 526.000 91.600 526.800 92.400 ;
        RECT 545.200 91.600 546.000 92.400 ;
        RECT 505.200 84.200 506.000 85.000 ;
        RECT 506.800 84.200 507.600 85.000 ;
        RECT 529.200 86.800 530.000 87.600 ;
        RECT 532.400 86.200 533.200 87.000 ;
        RECT 527.600 84.200 528.400 85.000 ;
        RECT 529.200 84.200 530.000 85.000 ;
        RECT 530.800 84.200 531.600 85.000 ;
        RECT 535.600 86.200 536.400 87.000 ;
        RECT 538.800 86.200 539.600 87.000 ;
        RECT 540.400 84.200 541.200 85.000 ;
        RECT 542.000 84.200 542.800 85.000 ;
        RECT 15.600 77.600 16.400 78.400 ;
        RECT 1.200 65.600 2.000 66.400 ;
        RECT 6.000 65.600 6.800 66.400 ;
        RECT 23.600 77.600 24.400 78.400 ;
        RECT 9.200 65.600 10.000 66.400 ;
        RECT 17.200 65.600 18.000 66.400 ;
        RECT 18.800 65.600 19.600 66.400 ;
        RECT 25.200 65.600 26.000 66.400 ;
        RECT 30.000 65.600 30.800 66.400 ;
        RECT 34.800 65.600 35.600 66.400 ;
        RECT 39.600 67.600 40.400 68.400 ;
        RECT 46.000 69.600 46.800 70.400 ;
        RECT 49.200 69.600 50.000 70.400 ;
        RECT 54.000 69.600 54.800 70.400 ;
        RECT 65.200 77.600 66.000 78.400 ;
        RECT 82.800 77.600 83.600 78.400 ;
        RECT 81.200 73.600 82.000 74.400 ;
        RECT 87.600 77.600 88.400 78.400 ;
        RECT 86.000 73.600 86.800 74.400 ;
        RECT 42.800 65.600 43.600 66.400 ;
        RECT 55.600 67.600 56.400 68.400 ;
        RECT 62.000 67.600 62.800 68.400 ;
        RECT 87.600 69.600 88.400 70.400 ;
        RECT 103.600 74.400 104.400 75.200 ;
        RECT 106.800 75.000 107.600 75.800 ;
        RECT 134.000 77.600 134.800 78.400 ;
        RECT 102.000 72.400 102.800 73.200 ;
        RECT 49.200 63.600 50.000 64.400 ;
        RECT 92.400 63.600 93.200 64.400 ;
        RECT 111.600 67.600 112.400 68.400 ;
        RECT 108.400 65.600 109.200 66.400 ;
        RECT 102.000 64.200 102.800 65.000 ;
        RECT 103.600 64.200 104.400 65.000 ;
        RECT 105.200 64.200 106.000 65.000 ;
        RECT 106.800 64.200 107.600 65.000 ;
        RECT 110.000 64.200 110.800 65.000 ;
        RECT 113.200 64.200 114.000 65.000 ;
        RECT 114.800 64.200 115.600 65.000 ;
        RECT 116.400 64.200 117.200 65.000 ;
        RECT 145.200 74.400 146.000 75.200 ;
        RECT 148.400 75.000 149.200 75.800 ;
        RECT 143.600 72.400 144.400 73.200 ;
        RECT 162.800 71.600 163.600 72.400 ;
        RECT 153.200 67.600 154.000 68.400 ;
        RECT 150.000 65.600 150.800 66.400 ;
        RECT 143.600 64.200 144.400 65.000 ;
        RECT 145.200 64.200 146.000 65.000 ;
        RECT 146.800 64.200 147.600 65.000 ;
        RECT 148.400 64.200 149.200 65.000 ;
        RECT 151.600 64.200 152.400 65.000 ;
        RECT 154.800 64.200 155.600 65.000 ;
        RECT 156.400 64.200 157.200 65.000 ;
        RECT 158.000 64.200 158.800 65.000 ;
        RECT 167.600 73.600 168.400 74.400 ;
        RECT 190.000 75.000 190.800 75.800 ;
        RECT 186.800 73.600 187.600 74.400 ;
        RECT 204.400 77.600 205.200 78.400 ;
        RECT 191.600 72.400 192.400 73.200 ;
        RECT 209.200 77.600 210.000 78.400 ;
        RECT 196.400 69.600 197.200 70.400 ;
        RECT 180.400 68.200 181.200 69.000 ;
        RECT 190.000 68.600 190.800 69.400 ;
        RECT 185.200 67.600 186.000 68.400 ;
        RECT 180.400 64.200 181.200 65.000 ;
        RECT 182.000 64.200 182.800 65.000 ;
        RECT 183.600 64.200 184.400 65.000 ;
        RECT 186.800 64.200 187.600 65.000 ;
        RECT 190.000 64.200 190.800 65.000 ;
        RECT 191.600 64.200 192.400 65.000 ;
        RECT 193.200 64.200 194.000 65.000 ;
        RECT 194.800 64.200 195.600 65.000 ;
        RECT 220.400 74.400 221.200 75.200 ;
        RECT 223.600 75.000 224.400 75.800 ;
        RECT 218.800 72.400 219.600 73.200 ;
        RECT 217.200 69.600 218.000 70.400 ;
        RECT 228.400 67.600 229.200 68.400 ;
        RECT 225.200 65.600 226.000 66.400 ;
        RECT 218.800 64.200 219.600 65.000 ;
        RECT 220.400 64.200 221.200 65.000 ;
        RECT 222.000 64.200 222.800 65.000 ;
        RECT 223.600 64.200 224.400 65.000 ;
        RECT 226.800 64.200 227.600 65.000 ;
        RECT 230.000 64.200 230.800 65.000 ;
        RECT 231.600 64.200 232.400 65.000 ;
        RECT 233.200 64.200 234.000 65.000 ;
        RECT 252.400 69.600 253.200 70.400 ;
        RECT 286.000 74.400 286.800 75.200 ;
        RECT 289.200 75.000 290.000 75.800 ;
        RECT 284.400 72.400 285.200 73.200 ;
        RECT 242.800 65.600 243.600 66.400 ;
        RECT 247.600 65.600 248.400 66.400 ;
        RECT 262.000 67.600 262.800 68.400 ;
        RECT 255.600 63.600 256.400 64.400 ;
        RECT 263.600 65.600 264.400 66.400 ;
        RECT 303.600 71.600 304.400 72.400 ;
        RECT 294.000 67.600 294.800 68.400 ;
        RECT 290.800 65.600 291.600 66.400 ;
        RECT 310.000 69.600 310.800 70.400 ;
        RECT 334.000 75.600 334.800 76.400 ;
        RECT 284.400 64.200 285.200 65.000 ;
        RECT 286.000 64.200 286.800 65.000 ;
        RECT 287.600 64.200 288.400 65.000 ;
        RECT 289.200 64.200 290.000 65.000 ;
        RECT 292.400 64.200 293.200 65.000 ;
        RECT 295.600 64.200 296.400 65.000 ;
        RECT 297.200 64.200 298.000 65.000 ;
        RECT 298.800 64.200 299.600 65.000 ;
        RECT 311.600 67.600 312.400 68.400 ;
        RECT 319.600 67.600 320.400 68.400 ;
        RECT 327.600 69.600 328.400 70.400 ;
        RECT 330.800 69.600 331.600 70.400 ;
        RECT 324.400 65.600 325.200 66.400 ;
        RECT 327.600 63.600 328.400 64.400 ;
        RECT 350.000 74.400 350.800 75.200 ;
        RECT 353.200 75.000 354.000 75.800 ;
        RECT 348.400 72.400 349.200 73.200 ;
        RECT 358.000 67.600 358.800 68.400 ;
        RECT 354.800 65.600 355.600 66.400 ;
        RECT 374.000 69.600 374.800 70.400 ;
        RECT 375.600 69.600 376.400 70.400 ;
        RECT 380.400 69.600 381.200 70.400 ;
        RECT 388.400 69.600 389.200 70.400 ;
        RECT 348.400 64.200 349.200 65.000 ;
        RECT 350.000 64.200 350.800 65.000 ;
        RECT 351.600 64.200 352.400 65.000 ;
        RECT 353.200 64.200 354.000 65.000 ;
        RECT 356.400 64.200 357.200 65.000 ;
        RECT 359.600 64.200 360.400 65.000 ;
        RECT 361.200 64.200 362.000 65.000 ;
        RECT 362.800 64.200 363.600 65.000 ;
        RECT 393.200 67.600 394.000 68.400 ;
        RECT 380.400 63.600 381.200 64.400 ;
        RECT 391.600 63.600 392.400 64.400 ;
        RECT 399.600 67.600 400.400 68.400 ;
        RECT 394.800 65.600 395.600 66.400 ;
        RECT 398.000 65.600 398.800 66.400 ;
        RECT 404.400 65.600 405.200 66.400 ;
        RECT 406.000 65.600 406.800 66.400 ;
        RECT 402.800 63.600 403.600 64.400 ;
        RECT 417.200 77.600 418.000 78.400 ;
        RECT 428.400 74.400 429.200 75.200 ;
        RECT 431.600 75.000 432.400 75.800 ;
        RECT 426.800 72.400 427.600 73.200 ;
        RECT 457.200 77.600 458.000 78.400 ;
        RECT 436.400 67.600 437.200 68.400 ;
        RECT 433.200 65.600 434.000 66.400 ;
        RECT 426.800 64.200 427.600 65.000 ;
        RECT 428.400 64.200 429.200 65.000 ;
        RECT 430.000 64.200 430.800 65.000 ;
        RECT 431.600 64.200 432.400 65.000 ;
        RECT 434.800 64.200 435.600 65.000 ;
        RECT 438.000 64.200 438.800 65.000 ;
        RECT 439.600 64.200 440.400 65.000 ;
        RECT 441.200 64.200 442.000 65.000 ;
        RECT 450.800 63.600 451.600 64.400 ;
        RECT 458.800 65.600 459.600 66.400 ;
        RECT 468.400 65.600 469.200 66.400 ;
        RECT 484.400 69.600 485.200 70.400 ;
        RECT 502.000 77.600 502.800 78.400 ;
        RECT 482.800 65.600 483.600 66.400 ;
        RECT 487.600 67.600 488.400 68.400 ;
        RECT 494.000 69.600 494.800 70.400 ;
        RECT 502.000 69.600 502.800 70.400 ;
        RECT 503.600 67.600 504.400 68.400 ;
        RECT 527.600 74.400 528.400 75.200 ;
        RECT 530.800 75.000 531.600 75.800 ;
        RECT 526.000 72.400 526.800 73.200 ;
        RECT 516.200 67.600 517.000 68.400 ;
        RECT 497.200 63.600 498.000 64.400 ;
        RECT 511.600 63.600 512.400 64.400 ;
        RECT 535.600 67.600 536.400 68.400 ;
        RECT 532.400 65.600 533.200 66.400 ;
        RECT 526.000 64.200 526.800 65.000 ;
        RECT 527.600 64.200 528.400 65.000 ;
        RECT 529.200 64.200 530.000 65.000 ;
        RECT 530.800 64.200 531.600 65.000 ;
        RECT 534.000 64.200 534.800 65.000 ;
        RECT 537.200 64.200 538.000 65.000 ;
        RECT 538.800 64.200 539.600 65.000 ;
        RECT 540.400 64.200 541.200 65.000 ;
        RECT 7.600 57.600 8.400 58.400 ;
        RECT 15.600 57.600 16.400 58.400 ;
        RECT 38.000 57.600 38.800 58.400 ;
        RECT 10.800 53.600 11.600 54.400 ;
        RECT 23.600 53.600 24.400 54.400 ;
        RECT 31.600 53.600 32.400 54.400 ;
        RECT 15.600 49.600 16.400 50.400 ;
        RECT 20.400 43.600 21.200 44.400 ;
        RECT 49.200 53.000 50.000 53.800 ;
        RECT 58.800 52.600 59.600 53.400 ;
        RECT 46.000 51.600 46.800 52.400 ;
        RECT 87.600 57.600 88.400 58.400 ;
        RECT 50.800 48.800 51.600 49.600 ;
        RECT 55.600 47.600 56.400 48.400 ;
        RECT 52.400 46.200 53.200 47.000 ;
        RECT 49.200 44.200 50.000 45.000 ;
        RECT 50.800 44.200 51.600 45.000 ;
        RECT 55.600 46.200 56.400 47.000 ;
        RECT 58.800 46.200 59.600 47.000 ;
        RECT 60.400 44.200 61.200 45.000 ;
        RECT 62.000 44.200 62.800 45.000 ;
        RECT 63.600 44.200 64.400 45.000 ;
        RECT 98.800 53.000 99.600 53.800 ;
        RECT 108.400 52.600 109.200 53.400 ;
        RECT 123.000 51.600 123.800 52.400 ;
        RECT 100.400 48.800 101.200 49.600 ;
        RECT 105.200 47.600 106.000 48.400 ;
        RECT 102.000 46.200 102.800 47.000 ;
        RECT 98.800 44.200 99.600 45.000 ;
        RECT 100.400 44.200 101.200 45.000 ;
        RECT 105.200 46.200 106.000 47.000 ;
        RECT 108.400 46.200 109.200 47.000 ;
        RECT 110.000 44.200 110.800 45.000 ;
        RECT 111.600 44.200 112.400 45.000 ;
        RECT 113.200 44.200 114.000 45.000 ;
        RECT 135.600 51.600 136.400 52.400 ;
        RECT 145.200 49.600 146.000 50.400 ;
        RECT 142.000 43.600 142.800 44.400 ;
        RECT 158.000 51.600 158.800 52.400 ;
        RECT 159.600 49.600 160.400 50.400 ;
        RECT 174.000 53.600 174.800 54.400 ;
        RECT 185.200 53.000 186.000 53.800 ;
        RECT 194.800 52.600 195.600 53.400 ;
        RECT 215.600 51.600 216.400 52.400 ;
        RECT 186.800 48.800 187.600 49.600 ;
        RECT 191.600 47.600 192.400 48.400 ;
        RECT 188.400 46.200 189.200 47.000 ;
        RECT 185.200 44.200 186.000 45.000 ;
        RECT 186.800 44.200 187.600 45.000 ;
        RECT 191.600 46.200 192.400 47.000 ;
        RECT 194.800 46.200 195.600 47.000 ;
        RECT 196.400 44.200 197.200 45.000 ;
        RECT 198.000 44.200 198.800 45.000 ;
        RECT 199.600 44.200 200.400 45.000 ;
        RECT 236.200 51.600 237.000 52.400 ;
        RECT 252.400 55.600 253.200 56.400 ;
        RECT 254.000 54.200 254.800 55.000 ;
        RECT 233.200 49.600 234.000 50.400 ;
        RECT 262.000 50.000 262.800 50.800 ;
        RECT 247.600 46.800 248.400 47.600 ;
        RECT 250.800 46.200 251.600 47.000 ;
        RECT 246.000 44.200 246.800 45.000 ;
        RECT 247.600 44.200 248.400 45.000 ;
        RECT 249.200 44.200 250.000 45.000 ;
        RECT 254.000 46.200 254.800 47.000 ;
        RECT 257.200 46.200 258.000 47.000 ;
        RECT 258.800 44.200 259.600 45.000 ;
        RECT 260.400 44.200 261.200 45.000 ;
        RECT 289.200 53.000 290.000 53.800 ;
        RECT 298.800 52.600 299.600 53.400 ;
        RECT 313.200 57.600 314.000 58.400 ;
        RECT 290.800 48.800 291.600 49.600 ;
        RECT 295.600 47.600 296.400 48.400 ;
        RECT 292.400 46.200 293.200 47.000 ;
        RECT 289.200 44.200 290.000 45.000 ;
        RECT 290.800 44.200 291.600 45.000 ;
        RECT 295.600 46.200 296.400 47.000 ;
        RECT 298.800 46.200 299.600 47.000 ;
        RECT 300.400 44.200 301.200 45.000 ;
        RECT 302.000 44.200 302.800 45.000 ;
        RECT 303.600 44.200 304.400 45.000 ;
        RECT 318.000 53.600 318.800 54.400 ;
        RECT 327.600 53.000 328.400 53.800 ;
        RECT 337.200 52.600 338.000 53.400 ;
        RECT 321.200 51.600 322.000 52.400 ;
        RECT 343.600 51.600 344.400 52.400 ;
        RECT 329.200 48.800 330.000 49.600 ;
        RECT 334.000 47.600 334.800 48.400 ;
        RECT 330.800 46.200 331.600 47.000 ;
        RECT 327.600 44.200 328.400 45.000 ;
        RECT 329.200 44.200 330.000 45.000 ;
        RECT 334.000 46.200 334.800 47.000 ;
        RECT 337.200 46.200 338.000 47.000 ;
        RECT 338.800 44.200 339.600 45.000 ;
        RECT 340.400 44.200 341.200 45.000 ;
        RECT 342.000 44.200 342.800 45.000 ;
        RECT 367.600 57.600 368.400 58.400 ;
        RECT 358.000 51.600 358.800 52.400 ;
        RECT 369.200 49.600 370.000 50.400 ;
        RECT 382.000 53.000 382.800 53.800 ;
        RECT 391.600 52.600 392.400 53.400 ;
        RECT 406.000 57.600 406.800 58.400 ;
        RECT 377.200 51.600 378.000 52.400 ;
        RECT 410.800 51.600 411.600 52.400 ;
        RECT 383.600 48.800 384.400 49.600 ;
        RECT 388.400 47.600 389.200 48.400 ;
        RECT 385.200 46.200 386.000 47.000 ;
        RECT 382.000 44.200 382.800 45.000 ;
        RECT 383.600 44.200 384.400 45.000 ;
        RECT 388.400 46.200 389.200 47.000 ;
        RECT 391.600 46.200 392.400 47.000 ;
        RECT 393.200 44.200 394.000 45.000 ;
        RECT 394.800 44.200 395.600 45.000 ;
        RECT 396.400 44.200 397.200 45.000 ;
        RECT 442.800 57.600 443.600 58.400 ;
        RECT 438.000 53.600 438.800 54.400 ;
        RECT 418.800 47.600 419.600 48.400 ;
        RECT 458.800 55.600 459.600 56.400 ;
        RECT 460.400 54.200 461.200 55.000 ;
        RECT 450.800 51.600 451.600 52.400 ;
        RECT 473.200 51.600 474.000 52.400 ;
        RECT 454.000 46.800 454.800 47.600 ;
        RECT 457.200 46.200 458.000 47.000 ;
        RECT 452.400 44.200 453.200 45.000 ;
        RECT 454.000 44.200 454.800 45.000 ;
        RECT 455.600 44.200 456.400 45.000 ;
        RECT 460.400 46.200 461.200 47.000 ;
        RECT 463.600 46.200 464.400 47.000 ;
        RECT 465.200 44.200 466.000 45.000 ;
        RECT 466.800 44.200 467.600 45.000 ;
        RECT 514.800 57.600 515.600 58.400 ;
        RECT 482.800 51.600 483.600 52.400 ;
        RECT 484.400 51.600 485.200 52.400 ;
        RECT 479.600 49.600 480.400 50.400 ;
        RECT 478.000 43.600 478.800 44.400 ;
        RECT 497.200 51.600 498.000 52.400 ;
        RECT 503.600 53.600 504.400 54.400 ;
        RECT 511.600 53.600 512.400 54.400 ;
        RECT 505.200 49.600 506.000 50.400 ;
        RECT 530.800 55.600 531.600 56.400 ;
        RECT 532.400 54.200 533.200 55.000 ;
        RECT 534.000 51.600 534.800 52.400 ;
        RECT 542.000 51.600 542.800 52.400 ;
        RECT 526.000 46.800 526.800 47.600 ;
        RECT 529.200 46.200 530.000 47.000 ;
        RECT 524.400 44.200 525.200 45.000 ;
        RECT 526.000 44.200 526.800 45.000 ;
        RECT 527.600 44.200 528.400 45.000 ;
        RECT 532.400 46.200 533.200 47.000 ;
        RECT 535.600 46.200 536.400 47.000 ;
        RECT 537.200 44.200 538.000 45.000 ;
        RECT 538.800 44.200 539.600 45.000 ;
        RECT 2.800 37.600 3.600 38.400 ;
        RECT 14.000 34.400 14.800 35.200 ;
        RECT 17.200 35.000 18.000 35.800 ;
        RECT 38.000 37.600 38.800 38.400 ;
        RECT 12.400 32.400 13.200 33.200 ;
        RECT 22.000 27.600 22.800 28.400 ;
        RECT 18.800 25.600 19.600 26.400 ;
        RECT 12.400 24.200 13.200 25.000 ;
        RECT 14.000 24.200 14.800 25.000 ;
        RECT 15.600 24.200 16.400 25.000 ;
        RECT 17.200 24.200 18.000 25.000 ;
        RECT 20.400 24.200 21.200 25.000 ;
        RECT 23.600 24.200 24.400 25.000 ;
        RECT 25.200 24.200 26.000 25.000 ;
        RECT 26.800 24.200 27.600 25.000 ;
        RECT 49.200 34.400 50.000 35.200 ;
        RECT 52.400 35.000 53.200 35.800 ;
        RECT 47.600 32.400 48.400 33.200 ;
        RECT 46.000 29.600 46.800 30.400 ;
        RECT 57.200 27.600 58.000 28.400 ;
        RECT 54.000 25.600 54.800 26.400 ;
        RECT 47.600 24.200 48.400 25.000 ;
        RECT 49.200 24.200 50.000 25.000 ;
        RECT 50.800 24.200 51.600 25.000 ;
        RECT 52.400 24.200 53.200 25.000 ;
        RECT 55.600 24.200 56.400 25.000 ;
        RECT 58.800 24.200 59.600 25.000 ;
        RECT 60.400 24.200 61.200 25.000 ;
        RECT 62.000 24.200 62.800 25.000 ;
        RECT 74.800 29.600 75.600 30.400 ;
        RECT 108.400 35.000 109.200 35.800 ;
        RECT 105.200 33.600 106.000 34.400 ;
        RECT 110.000 32.400 110.800 33.200 ;
        RECT 134.000 37.600 134.800 38.400 ;
        RECT 114.800 29.600 115.600 30.400 ;
        RECT 98.800 28.200 99.600 29.000 ;
        RECT 108.400 28.600 109.200 29.400 ;
        RECT 87.600 23.600 88.400 24.400 ;
        RECT 103.600 27.600 104.400 28.400 ;
        RECT 98.800 24.200 99.600 25.000 ;
        RECT 100.400 24.200 101.200 25.000 ;
        RECT 102.000 24.200 102.800 25.000 ;
        RECT 105.200 24.200 106.000 25.000 ;
        RECT 108.400 24.200 109.200 25.000 ;
        RECT 110.000 24.200 110.800 25.000 ;
        RECT 111.600 24.200 112.400 25.000 ;
        RECT 113.200 24.200 114.000 25.000 ;
        RECT 145.200 34.400 146.000 35.200 ;
        RECT 148.400 35.000 149.200 35.800 ;
        RECT 169.200 37.600 170.000 38.400 ;
        RECT 143.600 32.400 144.400 33.200 ;
        RECT 162.800 31.600 163.600 32.400 ;
        RECT 122.800 23.600 123.600 24.400 ;
        RECT 153.200 27.600 154.000 28.400 ;
        RECT 150.000 25.600 150.800 26.400 ;
        RECT 143.600 24.200 144.400 25.000 ;
        RECT 145.200 24.200 146.000 25.000 ;
        RECT 146.800 24.200 147.600 25.000 ;
        RECT 148.400 24.200 149.200 25.000 ;
        RECT 151.600 24.200 152.400 25.000 ;
        RECT 154.800 24.200 155.600 25.000 ;
        RECT 156.400 24.200 157.200 25.000 ;
        RECT 158.000 24.200 158.800 25.000 ;
        RECT 180.400 34.400 181.200 35.200 ;
        RECT 183.600 35.000 184.400 35.800 ;
        RECT 178.800 32.400 179.600 33.200 ;
        RECT 194.800 31.200 195.600 32.000 ;
        RECT 188.400 27.600 189.200 28.400 ;
        RECT 185.200 25.600 186.000 26.400 ;
        RECT 210.800 29.600 211.600 30.400 ;
        RECT 178.800 24.200 179.600 25.000 ;
        RECT 180.400 24.200 181.200 25.000 ;
        RECT 182.000 24.200 182.800 25.000 ;
        RECT 183.600 24.200 184.400 25.000 ;
        RECT 186.800 24.200 187.600 25.000 ;
        RECT 190.000 24.200 190.800 25.000 ;
        RECT 191.600 24.200 192.400 25.000 ;
        RECT 193.200 24.200 194.000 25.000 ;
        RECT 202.800 27.600 203.600 28.400 ;
        RECT 204.400 27.600 205.200 28.400 ;
        RECT 212.400 27.600 213.200 28.400 ;
        RECT 214.000 25.600 214.800 26.400 ;
        RECT 242.800 34.400 243.600 35.200 ;
        RECT 246.000 35.000 246.800 35.800 ;
        RECT 241.200 32.400 242.000 33.200 ;
        RECT 231.600 23.600 232.400 24.400 ;
        RECT 250.800 27.600 251.600 28.400 ;
        RECT 247.600 25.600 248.400 26.400 ;
        RECT 241.200 24.200 242.000 25.000 ;
        RECT 242.800 24.200 243.600 25.000 ;
        RECT 244.400 24.200 245.200 25.000 ;
        RECT 246.000 24.200 246.800 25.000 ;
        RECT 249.200 24.200 250.000 25.000 ;
        RECT 252.400 24.200 253.200 25.000 ;
        RECT 254.000 24.200 254.800 25.000 ;
        RECT 255.600 24.200 256.400 25.000 ;
        RECT 270.000 29.600 270.800 30.400 ;
        RECT 300.400 34.400 301.200 35.200 ;
        RECT 303.600 35.000 304.400 35.800 ;
        RECT 298.800 32.400 299.600 33.200 ;
        RECT 265.200 25.600 266.000 26.400 ;
        RECT 271.600 27.600 272.400 28.400 ;
        RECT 286.000 27.600 286.800 28.400 ;
        RECT 314.800 31.200 315.600 32.000 ;
        RECT 266.800 23.600 267.600 24.400 ;
        RECT 289.200 23.600 290.000 24.400 ;
        RECT 308.400 27.600 309.200 28.400 ;
        RECT 305.200 25.600 306.000 26.400 ;
        RECT 298.800 24.200 299.600 25.000 ;
        RECT 300.400 24.200 301.200 25.000 ;
        RECT 302.000 24.200 302.800 25.000 ;
        RECT 303.600 24.200 304.400 25.000 ;
        RECT 306.800 24.200 307.600 25.000 ;
        RECT 310.000 24.200 310.800 25.000 ;
        RECT 311.600 24.200 312.400 25.000 ;
        RECT 313.200 24.200 314.000 25.000 ;
        RECT 335.600 34.400 336.400 35.200 ;
        RECT 338.800 35.000 339.600 35.800 ;
        RECT 334.000 32.400 334.800 33.200 ;
        RECT 324.200 29.600 325.000 30.400 ;
        RECT 343.600 27.600 344.400 28.400 ;
        RECT 340.400 25.600 341.200 26.400 ;
        RECT 334.000 24.200 334.800 25.000 ;
        RECT 335.600 24.200 336.400 25.000 ;
        RECT 337.200 24.200 338.000 25.000 ;
        RECT 338.800 24.200 339.600 25.000 ;
        RECT 342.000 24.200 342.800 25.000 ;
        RECT 345.200 24.200 346.000 25.000 ;
        RECT 346.800 24.200 347.600 25.000 ;
        RECT 348.400 24.200 349.200 25.000 ;
        RECT 390.000 35.000 390.800 35.800 ;
        RECT 386.800 33.600 387.600 34.400 ;
        RECT 404.400 37.600 405.200 38.400 ;
        RECT 391.600 32.400 392.400 33.200 ;
        RECT 396.400 29.600 397.200 30.400 ;
        RECT 380.400 28.200 381.200 29.000 ;
        RECT 390.000 28.600 390.800 29.400 ;
        RECT 359.600 23.600 360.400 24.400 ;
        RECT 385.200 27.600 386.000 28.400 ;
        RECT 380.400 24.200 381.200 25.000 ;
        RECT 382.000 24.200 382.800 25.000 ;
        RECT 383.600 24.200 384.400 25.000 ;
        RECT 386.800 24.200 387.600 25.000 ;
        RECT 390.000 24.200 390.800 25.000 ;
        RECT 391.600 24.200 392.400 25.000 ;
        RECT 393.200 24.200 394.000 25.000 ;
        RECT 394.800 24.200 395.600 25.000 ;
        RECT 407.600 25.600 408.400 26.400 ;
        RECT 434.800 35.000 435.600 35.800 ;
        RECT 431.600 33.600 432.400 34.400 ;
        RECT 449.200 37.600 450.000 38.400 ;
        RECT 436.400 32.400 437.200 33.200 ;
        RECT 425.200 28.200 426.000 29.000 ;
        RECT 434.800 28.600 435.600 29.400 ;
        RECT 430.000 27.600 430.800 28.400 ;
        RECT 425.200 24.200 426.000 25.000 ;
        RECT 426.800 24.200 427.600 25.000 ;
        RECT 428.400 24.200 429.200 25.000 ;
        RECT 431.600 24.200 432.400 25.000 ;
        RECT 434.800 24.200 435.600 25.000 ;
        RECT 436.400 24.200 437.200 25.000 ;
        RECT 438.000 24.200 438.800 25.000 ;
        RECT 439.600 24.200 440.400 25.000 ;
        RECT 466.800 32.400 467.600 33.200 ;
        RECT 470.000 31.000 470.800 31.800 ;
        RECT 482.800 37.600 483.600 38.400 ;
        RECT 476.400 29.600 477.200 30.400 ;
        RECT 494.000 34.400 494.800 35.200 ;
        RECT 497.200 35.000 498.000 35.800 ;
        RECT 492.400 32.400 493.200 33.200 ;
        RECT 470.000 26.200 470.800 27.000 ;
        RECT 471.600 25.600 472.400 26.400 ;
        RECT 490.800 29.600 491.600 30.400 ;
        RECT 479.600 23.600 480.400 24.400 ;
        RECT 502.000 27.600 502.800 28.400 ;
        RECT 498.800 25.600 499.600 26.400 ;
        RECT 530.800 37.600 531.600 38.400 ;
        RECT 492.400 24.200 493.200 25.000 ;
        RECT 494.000 24.200 494.800 25.000 ;
        RECT 495.600 24.200 496.400 25.000 ;
        RECT 497.200 24.200 498.000 25.000 ;
        RECT 500.400 24.200 501.200 25.000 ;
        RECT 503.600 24.200 504.400 25.000 ;
        RECT 505.200 24.200 506.000 25.000 ;
        RECT 506.800 24.200 507.600 25.000 ;
        RECT 522.800 29.600 523.600 30.400 ;
        RECT 524.400 29.600 525.200 30.400 ;
        RECT 527.600 29.600 528.400 30.400 ;
        RECT 546.800 37.600 547.600 38.400 ;
        RECT 2.800 17.600 3.600 18.400 ;
        RECT 18.800 15.600 19.600 16.400 ;
        RECT 20.400 14.200 21.200 15.000 ;
        RECT 31.600 11.600 32.400 12.400 ;
        RECT 14.000 6.800 14.800 7.600 ;
        RECT 17.200 6.200 18.000 7.000 ;
        RECT 12.400 4.200 13.200 5.000 ;
        RECT 14.000 4.200 14.800 5.000 ;
        RECT 15.600 4.200 16.400 5.000 ;
        RECT 20.400 6.200 21.200 7.000 ;
        RECT 23.600 6.200 24.400 7.000 ;
        RECT 44.400 13.000 45.200 13.800 ;
        RECT 54.000 12.600 54.800 13.400 ;
        RECT 60.400 11.600 61.200 12.400 ;
        RECT 68.600 11.600 69.400 12.400 ;
        RECT 46.000 8.800 46.800 9.600 ;
        RECT 50.800 7.600 51.600 8.400 ;
        RECT 25.200 4.200 26.000 5.000 ;
        RECT 26.800 4.200 27.600 5.000 ;
        RECT 47.600 6.200 48.400 7.000 ;
        RECT 44.400 4.200 45.200 5.000 ;
        RECT 46.000 4.200 46.800 5.000 ;
        RECT 50.800 6.200 51.600 7.000 ;
        RECT 54.000 6.200 54.800 7.000 ;
        RECT 55.600 4.200 56.400 5.000 ;
        RECT 57.200 4.200 58.000 5.000 ;
        RECT 58.800 4.200 59.600 5.000 ;
        RECT 78.000 13.600 78.800 14.400 ;
        RECT 92.400 13.000 93.200 13.800 ;
        RECT 102.000 12.600 102.800 13.400 ;
        RECT 90.800 11.600 91.600 12.400 ;
        RECT 116.600 11.600 117.400 12.400 ;
        RECT 94.000 8.800 94.800 9.600 ;
        RECT 98.800 7.600 99.600 8.400 ;
        RECT 95.600 6.200 96.400 7.000 ;
        RECT 92.400 4.200 93.200 5.000 ;
        RECT 94.000 4.200 94.800 5.000 ;
        RECT 98.800 6.200 99.600 7.000 ;
        RECT 102.000 6.200 102.800 7.000 ;
        RECT 103.600 4.200 104.400 5.000 ;
        RECT 105.200 4.200 106.000 5.000 ;
        RECT 106.800 4.200 107.600 5.000 ;
        RECT 154.800 15.600 155.600 16.400 ;
        RECT 156.400 14.200 157.200 15.000 ;
        RECT 166.000 11.600 166.800 12.400 ;
        RECT 150.000 6.800 150.800 7.600 ;
        RECT 153.200 6.200 154.000 7.000 ;
        RECT 148.400 4.200 149.200 5.000 ;
        RECT 150.000 4.200 150.800 5.000 ;
        RECT 151.600 4.200 152.400 5.000 ;
        RECT 156.400 6.200 157.200 7.000 ;
        RECT 159.600 6.200 160.400 7.000 ;
        RECT 190.000 13.000 190.800 13.800 ;
        RECT 161.200 4.200 162.000 5.000 ;
        RECT 162.800 4.200 163.600 5.000 ;
        RECT 199.600 12.600 200.400 13.400 ;
        RECT 214.000 17.600 214.800 18.400 ;
        RECT 191.600 8.800 192.400 9.600 ;
        RECT 196.400 7.600 197.200 8.400 ;
        RECT 193.200 6.200 194.000 7.000 ;
        RECT 190.000 4.200 190.800 5.000 ;
        RECT 191.600 4.200 192.400 5.000 ;
        RECT 196.400 6.200 197.200 7.000 ;
        RECT 199.600 6.200 200.400 7.000 ;
        RECT 201.200 4.200 202.000 5.000 ;
        RECT 202.800 4.200 203.600 5.000 ;
        RECT 204.400 4.200 205.200 5.000 ;
        RECT 223.600 13.600 224.400 14.400 ;
        RECT 225.200 9.600 226.000 10.400 ;
        RECT 231.600 9.600 232.400 10.400 ;
        RECT 263.600 13.600 264.400 14.400 ;
        RECT 236.400 9.600 237.200 10.400 ;
        RECT 242.800 9.600 243.600 10.400 ;
        RECT 249.200 9.600 250.000 10.400 ;
        RECT 254.000 7.600 254.800 8.400 ;
        RECT 287.600 17.600 288.400 18.400 ;
        RECT 268.400 13.600 269.200 14.400 ;
        RECT 274.800 9.600 275.600 10.400 ;
        RECT 290.600 11.600 291.400 12.400 ;
        RECT 306.800 15.600 307.600 16.400 ;
        RECT 308.400 14.200 309.200 15.000 ;
        RECT 335.600 17.600 336.400 18.400 ;
        RECT 287.600 9.600 288.400 10.400 ;
        RECT 302.000 6.800 302.800 7.600 ;
        RECT 305.200 6.200 306.000 7.000 ;
        RECT 300.400 4.200 301.200 5.000 ;
        RECT 302.000 4.200 302.800 5.000 ;
        RECT 303.600 4.200 304.400 5.000 ;
        RECT 308.400 6.200 309.200 7.000 ;
        RECT 311.600 6.200 312.400 7.000 ;
        RECT 324.400 13.600 325.200 14.400 ;
        RECT 330.800 13.600 331.600 14.400 ;
        RECT 313.200 4.200 314.000 5.000 ;
        RECT 314.800 4.200 315.600 5.000 ;
        RECT 354.800 15.600 355.600 16.400 ;
        RECT 356.400 14.200 357.200 15.000 ;
        RECT 367.600 11.600 368.400 12.400 ;
        RECT 338.800 9.600 339.600 10.400 ;
        RECT 350.000 6.800 350.800 7.600 ;
        RECT 353.200 6.200 354.000 7.000 ;
        RECT 348.400 4.200 349.200 5.000 ;
        RECT 350.000 4.200 350.800 5.000 ;
        RECT 351.600 4.200 352.400 5.000 ;
        RECT 356.400 6.200 357.200 7.000 ;
        RECT 359.600 6.200 360.400 7.000 ;
        RECT 386.800 13.600 387.600 14.400 ;
        RECT 382.000 12.200 382.800 13.000 ;
        RECT 361.200 4.200 362.000 5.000 ;
        RECT 362.800 4.200 363.600 5.000 ;
        RECT 404.400 13.000 405.200 13.800 ;
        RECT 390.000 11.800 390.800 12.600 ;
        RECT 394.800 10.200 395.600 11.000 ;
        RECT 414.000 12.600 414.800 13.400 ;
        RECT 428.400 17.600 429.200 18.400 ;
        RECT 399.600 11.600 400.400 12.400 ;
        RECT 420.400 11.600 421.200 12.400 ;
        RECT 442.800 11.800 443.600 12.600 ;
        RECT 406.000 8.800 406.800 9.600 ;
        RECT 410.800 7.600 411.600 8.400 ;
        RECT 407.600 6.200 408.400 7.000 ;
        RECT 404.400 4.200 405.200 5.000 ;
        RECT 406.000 4.200 406.800 5.000 ;
        RECT 410.800 6.200 411.600 7.000 ;
        RECT 414.000 6.200 414.800 7.000 ;
        RECT 415.600 4.200 416.400 5.000 ;
        RECT 417.200 4.200 418.000 5.000 ;
        RECT 418.800 4.200 419.600 5.000 ;
        RECT 438.000 10.200 438.800 11.000 ;
        RECT 474.800 13.000 475.600 13.800 ;
        RECT 484.400 12.600 485.200 13.400 ;
        RECT 498.800 17.600 499.600 18.400 ;
        RECT 503.600 17.600 504.400 18.400 ;
        RECT 473.200 11.600 474.000 12.400 ;
        RECT 490.800 11.600 491.600 12.400 ;
        RECT 476.400 8.800 477.200 9.600 ;
        RECT 481.200 7.600 482.000 8.400 ;
        RECT 478.000 6.200 478.800 7.000 ;
        RECT 474.800 4.200 475.600 5.000 ;
        RECT 476.400 4.200 477.200 5.000 ;
        RECT 481.200 6.200 482.000 7.000 ;
        RECT 484.400 6.200 485.200 7.000 ;
        RECT 486.000 4.200 486.800 5.000 ;
        RECT 487.600 4.200 488.400 5.000 ;
        RECT 489.200 4.200 490.000 5.000 ;
        RECT 513.200 13.000 514.000 13.800 ;
        RECT 522.800 12.600 523.600 13.400 ;
        RECT 510.000 11.600 510.800 12.400 ;
        RECT 514.800 8.800 515.600 9.600 ;
        RECT 519.600 7.600 520.400 8.400 ;
        RECT 516.400 6.200 517.200 7.000 ;
        RECT 513.200 4.200 514.000 5.000 ;
        RECT 514.800 4.200 515.600 5.000 ;
        RECT 519.600 6.200 520.400 7.000 ;
        RECT 522.800 6.200 523.600 7.000 ;
        RECT 524.400 4.200 525.200 5.000 ;
        RECT 526.000 4.200 526.800 5.000 ;
        RECT 527.600 4.200 528.400 5.000 ;
      LAYER metal2 ;
        RECT 1.200 367.600 2.000 368.400 ;
        RECT 1.300 336.400 1.900 367.600 ;
        RECT 12.400 364.200 13.200 377.800 ;
        RECT 14.000 364.200 14.800 377.800 ;
        RECT 15.600 364.200 16.400 377.800 ;
        RECT 17.200 366.200 18.000 377.800 ;
        RECT 18.800 375.600 19.600 376.400 ;
        RECT 2.800 343.600 3.600 344.400 ;
        RECT 12.400 344.200 13.200 357.800 ;
        RECT 14.000 344.200 14.800 357.800 ;
        RECT 15.600 344.200 16.400 357.800 ;
        RECT 17.200 344.200 18.000 355.800 ;
        RECT 18.900 346.400 19.500 375.600 ;
        RECT 20.400 366.200 21.200 377.800 ;
        RECT 22.000 373.600 22.800 374.400 ;
        RECT 23.600 366.200 24.400 377.800 ;
        RECT 25.200 364.200 26.000 377.800 ;
        RECT 26.800 364.200 27.600 377.800 ;
        RECT 28.400 371.600 29.200 372.400 ;
        RECT 31.600 371.600 32.400 372.400 ;
        RECT 38.000 371.600 38.800 372.400 ;
        RECT 18.800 345.600 19.600 346.400 ;
        RECT 18.900 340.400 19.500 345.600 ;
        RECT 20.400 344.200 21.200 355.800 ;
        RECT 22.000 347.600 22.800 348.400 ;
        RECT 23.600 344.200 24.400 355.800 ;
        RECT 25.200 344.200 26.000 357.800 ;
        RECT 26.800 344.200 27.600 357.800 ;
        RECT 28.500 350.400 29.100 371.600 ;
        RECT 44.400 364.200 45.200 377.800 ;
        RECT 46.000 364.200 46.800 377.800 ;
        RECT 47.600 366.200 48.400 377.800 ;
        RECT 49.200 373.600 50.000 374.400 ;
        RECT 49.300 364.300 49.900 373.600 ;
        RECT 50.800 366.200 51.600 377.800 ;
        RECT 52.400 375.600 53.200 376.400 ;
        RECT 54.000 366.200 54.800 377.800 ;
        RECT 49.300 363.700 51.500 364.300 ;
        RECT 55.600 364.200 56.400 377.800 ;
        RECT 57.200 364.200 58.000 377.800 ;
        RECT 58.800 364.200 59.600 377.800 ;
        RECT 60.400 371.600 61.200 372.400 ;
        RECT 38.000 357.600 38.800 358.400 ;
        RECT 44.400 357.600 45.200 358.400 ;
        RECT 49.200 357.600 50.000 358.400 ;
        RECT 28.400 349.600 29.200 350.400 ;
        RECT 31.600 349.600 32.400 350.400 ;
        RECT 18.800 339.600 19.600 340.400 ;
        RECT 22.000 339.600 22.800 340.400 ;
        RECT 1.200 335.600 2.000 336.400 ;
        RECT 1.300 312.400 1.900 335.600 ;
        RECT 4.400 327.600 5.200 328.400 ;
        RECT 2.800 323.600 3.600 324.400 ;
        RECT 2.900 318.400 3.500 323.600 ;
        RECT 2.800 317.600 3.600 318.400 ;
        RECT 1.200 311.600 2.000 312.400 ;
        RECT 1.300 310.400 1.900 311.600 ;
        RECT 1.200 309.600 2.000 310.400 ;
        RECT 4.500 306.400 5.100 327.600 ;
        RECT 15.600 324.200 16.400 337.800 ;
        RECT 17.200 324.200 18.000 337.800 ;
        RECT 18.800 324.200 19.600 337.800 ;
        RECT 20.400 326.200 21.200 337.800 ;
        RECT 22.100 336.400 22.700 339.600 ;
        RECT 22.000 335.600 22.800 336.400 ;
        RECT 23.600 326.200 24.400 337.800 ;
        RECT 25.200 333.600 26.000 334.400 ;
        RECT 25.300 330.400 25.900 333.600 ;
        RECT 25.200 329.600 26.000 330.400 ;
        RECT 26.800 326.200 27.600 337.800 ;
        RECT 28.400 324.200 29.200 337.800 ;
        RECT 30.000 324.200 30.800 337.800 ;
        RECT 31.700 332.400 32.300 349.600 ;
        RECT 38.100 346.400 38.700 357.600 ;
        RECT 42.800 351.600 43.600 352.400 ;
        RECT 42.900 346.400 43.500 351.600 ;
        RECT 44.500 350.400 45.100 357.600 ;
        RECT 47.600 351.600 48.400 352.400 ;
        RECT 44.400 349.600 45.200 350.400 ;
        RECT 44.400 347.600 45.200 348.400 ;
        RECT 38.000 345.600 38.800 346.400 ;
        RECT 42.800 345.600 43.600 346.400 ;
        RECT 39.600 343.600 40.400 344.400 ;
        RECT 41.200 343.600 42.000 344.400 ;
        RECT 39.700 334.400 40.300 343.600 ;
        RECT 39.600 333.600 40.400 334.400 ;
        RECT 31.600 331.600 32.400 332.400 ;
        RECT 30.000 321.600 30.800 322.400 ;
        RECT 30.100 318.400 30.700 321.600 ;
        RECT 17.200 317.600 18.000 318.400 ;
        RECT 25.200 317.600 26.000 318.400 ;
        RECT 30.000 317.600 30.800 318.400 ;
        RECT 31.600 317.600 32.400 318.400 ;
        RECT 17.300 314.400 17.900 317.600 ;
        RECT 9.200 313.600 10.000 314.400 ;
        RECT 12.400 313.600 13.200 314.400 ;
        RECT 17.200 313.600 18.000 314.400 ;
        RECT 23.600 313.600 24.400 314.400 ;
        RECT 25.300 312.400 25.900 317.600 ;
        RECT 6.000 311.600 6.800 312.400 ;
        RECT 22.000 311.600 22.800 312.400 ;
        RECT 25.200 311.600 26.000 312.400 ;
        RECT 26.800 312.300 27.600 312.400 ;
        RECT 26.800 311.700 29.100 312.300 ;
        RECT 26.800 311.600 27.600 311.700 ;
        RECT 7.600 309.600 8.400 310.400 ;
        RECT 18.800 309.600 19.600 310.400 ;
        RECT 1.200 305.600 2.000 306.400 ;
        RECT 4.400 305.600 5.200 306.400 ;
        RECT 1.300 256.400 1.900 305.600 ;
        RECT 4.400 291.600 5.200 292.400 ;
        RECT 2.800 289.600 3.600 290.400 ;
        RECT 2.900 278.400 3.500 289.600 ;
        RECT 4.500 288.300 5.100 291.600 ;
        RECT 6.000 289.600 6.800 290.400 ;
        RECT 7.700 288.300 8.300 309.600 ;
        RECT 22.100 308.400 22.700 311.600 ;
        RECT 23.600 309.600 24.400 310.400 ;
        RECT 22.000 307.600 22.800 308.400 ;
        RECT 22.100 306.400 22.700 307.600 ;
        RECT 14.000 305.600 14.800 306.400 ;
        RECT 22.000 305.600 22.800 306.400 ;
        RECT 10.800 303.600 11.600 304.400 ;
        RECT 18.800 303.600 19.600 304.400 ;
        RECT 18.900 298.400 19.500 303.600 ;
        RECT 18.800 297.600 19.600 298.400 ;
        RECT 10.800 295.600 11.600 296.400 ;
        RECT 12.400 295.600 13.200 296.400 ;
        RECT 14.000 295.600 14.800 296.400 ;
        RECT 18.800 295.600 19.600 296.400 ;
        RECT 20.400 295.600 21.200 296.400 ;
        RECT 10.900 292.400 11.500 295.600 ;
        RECT 14.100 292.400 14.700 295.600 ;
        RECT 23.700 292.400 24.300 309.600 ;
        RECT 28.500 298.400 29.100 311.700 ;
        RECT 30.000 309.600 30.800 310.400 ;
        RECT 30.100 308.400 30.700 309.600 ;
        RECT 31.700 308.400 32.300 317.600 ;
        RECT 38.000 313.600 38.800 314.400 ;
        RECT 36.400 309.600 37.200 310.400 ;
        RECT 30.000 307.600 30.800 308.400 ;
        RECT 31.600 307.600 32.400 308.400 ;
        RECT 33.200 305.600 34.000 306.400 ;
        RECT 34.800 305.600 35.600 306.400 ;
        RECT 33.300 304.400 33.900 305.600 ;
        RECT 33.200 303.600 34.000 304.400 ;
        RECT 28.400 297.600 29.200 298.400 ;
        RECT 33.200 297.600 34.000 298.400 ;
        RECT 33.300 296.400 33.900 297.600 ;
        RECT 36.500 296.400 37.100 309.600 ;
        RECT 38.100 306.400 38.700 313.600 ;
        RECT 38.000 305.600 38.800 306.400 ;
        RECT 39.700 304.300 40.300 333.600 ;
        RECT 41.300 332.400 41.900 343.600 ;
        RECT 44.500 338.400 45.100 347.600 ;
        RECT 47.700 346.400 48.300 351.600 ;
        RECT 49.300 346.400 49.900 357.600 ;
        RECT 47.600 345.600 48.400 346.400 ;
        RECT 49.200 345.600 50.000 346.400 ;
        RECT 46.000 343.600 46.800 344.400 ;
        RECT 44.400 337.600 45.200 338.400 ;
        RECT 46.100 334.400 46.700 343.600 ;
        RECT 50.900 342.400 51.500 363.700 ;
        RECT 54.000 351.600 54.800 352.400 ;
        RECT 57.200 351.600 58.000 352.400 ;
        RECT 54.100 348.400 54.700 351.600 ;
        RECT 54.000 347.600 54.800 348.400 ;
        RECT 52.400 345.600 53.200 346.400 ;
        RECT 50.800 341.600 51.600 342.400 ;
        RECT 52.500 340.400 53.100 345.600 ;
        RECT 52.400 339.600 53.200 340.400 ;
        RECT 57.300 338.400 57.900 351.600 ;
        RECT 60.500 350.400 61.100 371.600 ;
        RECT 73.200 367.600 74.000 368.400 ;
        RECT 68.400 363.600 69.200 364.400 ;
        RECT 73.300 358.400 73.900 367.600 ;
        RECT 82.800 364.200 83.600 377.800 ;
        RECT 84.400 364.200 85.200 377.800 ;
        RECT 86.000 364.200 86.800 377.800 ;
        RECT 87.600 366.200 88.400 377.800 ;
        RECT 89.200 375.600 90.000 376.400 ;
        RECT 60.400 349.600 61.200 350.400 ;
        RECT 66.800 344.200 67.600 357.800 ;
        RECT 68.400 344.200 69.200 357.800 ;
        RECT 73.200 357.600 74.000 358.400 ;
        RECT 70.000 344.200 70.800 355.800 ;
        RECT 71.600 347.600 72.400 348.400 ;
        RECT 68.400 341.600 69.200 342.400 ;
        RECT 57.200 337.600 58.000 338.400 ;
        RECT 49.200 335.600 50.000 336.400 ;
        RECT 49.300 334.400 49.900 335.600 ;
        RECT 46.000 333.600 46.800 334.400 ;
        RECT 49.200 333.600 50.000 334.400 ;
        RECT 52.400 333.600 53.200 334.400 ;
        RECT 63.600 334.300 64.400 334.400 ;
        RECT 62.100 333.700 64.400 334.300 ;
        RECT 52.500 332.400 53.100 333.600 ;
        RECT 41.200 331.600 42.000 332.400 ;
        RECT 47.600 331.600 48.400 332.400 ;
        RECT 52.400 331.600 53.200 332.400 ;
        RECT 57.200 331.600 58.000 332.400 ;
        RECT 58.800 331.600 59.600 332.400 ;
        RECT 42.800 329.600 43.600 330.400 ;
        RECT 44.400 329.600 45.200 330.400 ;
        RECT 42.900 328.400 43.500 329.600 ;
        RECT 42.800 327.600 43.600 328.400 ;
        RECT 44.500 318.400 45.100 329.600 ;
        RECT 47.700 326.400 48.300 331.600 ;
        RECT 57.300 330.400 57.900 331.600 ;
        RECT 58.900 330.400 59.500 331.600 ;
        RECT 50.800 329.600 51.600 330.400 ;
        RECT 57.200 329.600 58.000 330.400 ;
        RECT 58.800 329.600 59.600 330.400 ;
        RECT 54.000 327.600 54.800 328.400 ;
        RECT 58.900 328.300 59.500 329.600 ;
        RECT 57.300 327.700 59.500 328.300 ;
        RECT 47.600 325.600 48.400 326.400 ;
        RECT 52.400 325.600 53.200 326.400 ;
        RECT 44.400 317.600 45.200 318.400 ;
        RECT 54.100 316.400 54.700 327.600 ;
        RECT 57.300 318.400 57.900 327.700 ;
        RECT 60.400 327.600 61.200 328.400 ;
        RECT 57.200 317.600 58.000 318.400 ;
        RECT 60.500 316.400 61.100 327.600 ;
        RECT 47.600 315.600 48.400 316.400 ;
        RECT 52.400 315.600 53.200 316.400 ;
        RECT 54.000 315.600 54.800 316.400 ;
        RECT 60.400 315.600 61.200 316.400 ;
        RECT 41.200 313.600 42.000 314.400 ;
        RECT 42.800 311.600 43.600 312.400 ;
        RECT 44.400 311.600 45.200 312.400 ;
        RECT 41.200 309.600 42.000 310.400 ;
        RECT 38.100 303.700 40.300 304.300 ;
        RECT 33.200 295.600 34.000 296.400 ;
        RECT 36.400 295.600 37.200 296.400 ;
        RECT 33.200 293.600 34.000 294.400 ;
        RECT 10.800 291.600 11.600 292.400 ;
        RECT 14.000 291.600 14.800 292.400 ;
        RECT 22.000 291.600 22.800 292.400 ;
        RECT 23.600 291.600 24.400 292.400 ;
        RECT 14.100 290.400 14.700 291.600 ;
        RECT 22.100 290.400 22.700 291.600 ;
        RECT 14.000 289.600 14.800 290.400 ;
        RECT 22.000 289.600 22.800 290.400 ;
        RECT 28.400 289.600 29.200 290.400 ;
        RECT 4.500 287.700 8.300 288.300 ;
        RECT 4.400 283.600 5.200 284.400 ;
        RECT 2.800 277.600 3.600 278.400 ;
        RECT 4.500 256.400 5.100 283.600 ;
        RECT 1.200 255.600 2.000 256.400 ;
        RECT 4.400 255.600 5.200 256.400 ;
        RECT 4.400 251.600 5.200 252.400 ;
        RECT 4.400 229.600 5.200 230.400 ;
        RECT 2.800 224.300 3.600 224.400 ;
        RECT 4.500 224.300 5.100 229.600 ;
        RECT 2.800 223.700 5.100 224.300 ;
        RECT 2.800 223.600 3.600 223.700 ;
        RECT 4.500 214.400 5.100 223.700 ;
        RECT 6.100 222.400 6.700 287.700 ;
        RECT 18.800 287.600 19.600 288.400 ;
        RECT 25.200 287.600 26.000 288.400 ;
        RECT 23.600 283.600 24.400 284.400 ;
        RECT 18.800 281.600 19.600 282.400 ;
        RECT 12.400 264.200 13.200 277.800 ;
        RECT 14.000 264.200 14.800 277.800 ;
        RECT 15.600 264.200 16.400 277.800 ;
        RECT 17.200 264.200 18.000 275.800 ;
        RECT 18.900 266.400 19.500 281.600 ;
        RECT 23.700 278.400 24.300 283.600 ;
        RECT 23.600 277.600 24.400 278.400 ;
        RECT 18.800 265.600 19.600 266.400 ;
        RECT 9.200 255.600 10.000 256.400 ;
        RECT 14.000 255.600 14.800 256.400 ;
        RECT 9.300 254.400 9.900 255.600 ;
        RECT 14.100 254.400 14.700 255.600 ;
        RECT 9.200 253.600 10.000 254.400 ;
        RECT 14.000 253.600 14.800 254.400 ;
        RECT 7.600 251.600 8.400 252.400 ;
        RECT 12.400 251.600 13.200 252.400 ;
        RECT 15.600 251.600 16.400 252.400 ;
        RECT 12.500 250.400 13.100 251.600 ;
        RECT 12.400 249.600 13.200 250.400 ;
        RECT 10.800 247.600 11.600 248.400 ;
        RECT 18.900 246.400 19.500 265.600 ;
        RECT 20.400 264.200 21.200 275.800 ;
        RECT 22.000 273.600 22.800 274.400 ;
        RECT 22.100 268.400 22.700 273.600 ;
        RECT 22.000 267.600 22.800 268.400 ;
        RECT 23.600 264.200 24.400 275.800 ;
        RECT 25.200 264.200 26.000 277.800 ;
        RECT 26.800 264.200 27.600 277.800 ;
        RECT 28.500 272.400 29.100 289.600 ;
        RECT 30.000 275.600 30.800 276.400 ;
        RECT 28.400 271.600 29.200 272.400 ;
        RECT 30.100 270.400 30.700 275.600 ;
        RECT 28.400 269.600 29.200 270.400 ;
        RECT 30.000 269.600 30.800 270.400 ;
        RECT 23.600 257.600 24.400 258.400 ;
        RECT 23.700 256.400 24.300 257.600 ;
        RECT 23.600 255.600 24.400 256.400 ;
        RECT 20.400 253.600 21.200 254.400 ;
        RECT 25.200 253.600 26.000 254.400 ;
        RECT 20.500 252.400 21.100 253.600 ;
        RECT 20.400 251.600 21.200 252.400 ;
        RECT 23.600 251.600 24.400 252.400 ;
        RECT 26.800 251.600 27.600 252.400 ;
        RECT 18.800 245.600 19.600 246.400 ;
        RECT 7.600 243.600 8.400 244.400 ;
        RECT 18.800 243.600 19.600 244.400 ;
        RECT 6.000 221.600 6.800 222.400 ;
        RECT 6.100 216.400 6.700 221.600 ;
        RECT 7.700 216.400 8.300 243.600 ;
        RECT 12.400 224.200 13.200 237.800 ;
        RECT 14.000 224.200 14.800 237.800 ;
        RECT 15.600 224.200 16.400 237.800 ;
        RECT 17.200 224.200 18.000 235.800 ;
        RECT 18.900 228.400 19.500 243.600 ;
        RECT 18.800 227.600 19.600 228.400 ;
        RECT 18.800 225.600 19.600 226.400 ;
        RECT 20.400 224.200 21.200 235.800 ;
        RECT 22.000 231.600 22.800 232.400 ;
        RECT 22.100 228.400 22.700 231.600 ;
        RECT 22.000 227.600 22.800 228.400 ;
        RECT 22.000 225.600 22.800 226.400 ;
        RECT 22.100 222.300 22.700 225.600 ;
        RECT 23.600 224.200 24.400 235.800 ;
        RECT 25.200 224.200 26.000 237.800 ;
        RECT 26.800 224.200 27.600 237.800 ;
        RECT 28.500 230.400 29.100 269.600 ;
        RECT 30.000 267.600 30.800 268.400 ;
        RECT 30.100 258.400 30.700 267.600 ;
        RECT 30.000 257.600 30.800 258.400 ;
        RECT 31.600 255.600 32.400 256.400 ;
        RECT 31.700 254.400 32.300 255.600 ;
        RECT 31.600 253.600 32.400 254.400 ;
        RECT 31.600 251.600 32.400 252.400 ;
        RECT 30.000 243.600 30.800 244.400 ;
        RECT 28.400 229.600 29.200 230.400 ;
        RECT 30.100 224.400 30.700 243.600 ;
        RECT 30.000 223.600 30.800 224.400 ;
        RECT 20.500 221.700 22.700 222.300 ;
        RECT 15.600 217.600 16.400 218.400 ;
        RECT 6.000 215.600 6.800 216.400 ;
        RECT 7.600 215.600 8.400 216.400 ;
        RECT 17.200 215.600 18.000 216.400 ;
        RECT 4.400 213.600 5.200 214.400 ;
        RECT 6.100 212.400 6.700 215.600 ;
        RECT 17.300 214.400 17.900 215.600 ;
        RECT 9.200 213.600 10.000 214.400 ;
        RECT 12.400 213.600 13.200 214.400 ;
        RECT 15.600 213.600 16.400 214.400 ;
        RECT 17.200 213.600 18.000 214.400 ;
        RECT 18.800 213.600 19.600 214.400 ;
        RECT 9.300 212.400 9.900 213.600 ;
        RECT 6.000 211.600 6.800 212.400 ;
        RECT 9.200 211.600 10.000 212.400 ;
        RECT 12.500 208.400 13.100 213.600 ;
        RECT 12.400 207.600 13.200 208.400 ;
        RECT 2.800 203.600 3.600 204.400 ;
        RECT 1.200 187.600 2.000 188.400 ;
        RECT 1.300 176.400 1.900 187.600 ;
        RECT 1.200 175.600 2.000 176.400 ;
        RECT 2.900 152.400 3.500 203.600 ;
        RECT 4.400 191.600 5.200 192.400 ;
        RECT 6.000 191.600 6.800 192.400 ;
        RECT 10.800 191.600 11.600 192.400 ;
        RECT 4.500 190.400 5.100 191.600 ;
        RECT 10.900 190.400 11.500 191.600 ;
        RECT 4.400 189.600 5.200 190.400 ;
        RECT 6.000 189.600 6.800 190.400 ;
        RECT 10.800 189.600 11.600 190.400 ;
        RECT 4.400 183.600 5.200 184.400 ;
        RECT 4.500 176.400 5.100 183.600 ;
        RECT 4.400 175.600 5.200 176.400 ;
        RECT 6.100 170.300 6.700 189.600 ;
        RECT 9.200 187.600 10.000 188.400 ;
        RECT 9.300 186.400 9.900 187.600 ;
        RECT 9.200 185.600 10.000 186.400 ;
        RECT 7.600 183.600 8.400 184.400 ;
        RECT 7.700 176.400 8.300 183.600 ;
        RECT 10.900 176.400 11.500 189.600 ;
        RECT 12.500 176.400 13.100 207.600 ;
        RECT 14.000 185.600 14.800 186.400 ;
        RECT 7.600 175.600 8.400 176.400 ;
        RECT 9.200 175.600 10.000 176.400 ;
        RECT 10.800 175.600 11.600 176.400 ;
        RECT 12.400 175.600 13.200 176.400 ;
        RECT 9.200 171.600 10.000 172.400 ;
        RECT 12.400 172.300 13.200 172.400 ;
        RECT 10.900 171.700 13.200 172.300 ;
        RECT 6.100 169.700 8.300 170.300 ;
        RECT 4.400 157.600 5.200 158.400 ;
        RECT 2.800 151.600 3.600 152.400 ;
        RECT 4.500 150.400 5.100 157.600 ;
        RECT 7.700 154.400 8.300 169.700 ;
        RECT 7.600 153.600 8.400 154.400 ;
        RECT 6.000 151.600 6.800 152.400 ;
        RECT 4.400 149.600 5.200 150.400 ;
        RECT 7.600 149.600 8.400 150.400 ;
        RECT 7.600 143.600 8.400 144.400 ;
        RECT 7.700 138.400 8.300 143.600 ;
        RECT 2.800 137.600 3.600 138.400 ;
        RECT 7.600 137.600 8.400 138.400 ;
        RECT 2.900 134.400 3.500 137.600 ;
        RECT 4.400 135.600 5.200 136.400 ;
        RECT 7.600 135.600 8.400 136.400 ;
        RECT 2.800 133.600 3.600 134.400 ;
        RECT 4.500 132.400 5.100 135.600 ;
        RECT 6.000 133.600 6.800 134.400 ;
        RECT 4.400 131.600 5.200 132.400 ;
        RECT 7.700 130.400 8.300 135.600 ;
        RECT 9.200 131.600 10.000 132.400 ;
        RECT 7.600 129.600 8.400 130.400 ;
        RECT 10.900 130.300 11.500 171.700 ;
        RECT 12.400 171.600 13.200 171.700 ;
        RECT 14.000 172.300 14.800 172.400 ;
        RECT 15.700 172.300 16.300 213.600 ;
        RECT 17.200 211.600 18.000 212.400 ;
        RECT 18.800 210.300 19.600 210.400 ;
        RECT 20.500 210.300 21.100 221.700 ;
        RECT 22.000 219.600 22.800 220.400 ;
        RECT 28.400 219.600 29.200 220.400 ;
        RECT 31.600 219.600 32.400 220.400 ;
        RECT 22.100 214.400 22.700 219.600 ;
        RECT 26.800 215.600 27.600 216.400 ;
        RECT 22.000 213.600 22.800 214.400 ;
        RECT 26.900 212.400 27.500 215.600 ;
        RECT 26.800 211.600 27.600 212.400 ;
        RECT 28.500 210.400 29.100 219.600 ;
        RECT 30.000 215.600 30.800 216.400 ;
        RECT 30.100 214.400 30.700 215.600 ;
        RECT 30.000 213.600 30.800 214.400 ;
        RECT 18.800 209.700 21.100 210.300 ;
        RECT 18.800 209.600 19.600 209.700 ;
        RECT 26.800 209.600 27.600 210.400 ;
        RECT 28.400 209.600 29.200 210.400 ;
        RECT 25.200 207.600 26.000 208.400 ;
        RECT 26.900 206.400 27.500 209.600 ;
        RECT 30.100 208.400 30.700 213.600 ;
        RECT 31.700 212.400 32.300 219.600 ;
        RECT 31.600 211.600 32.400 212.400 ;
        RECT 30.000 207.600 30.800 208.400 ;
        RECT 26.800 205.600 27.600 206.400 ;
        RECT 33.300 200.400 33.900 293.600 ;
        RECT 36.500 292.400 37.100 295.600 ;
        RECT 38.100 292.400 38.700 303.700 ;
        RECT 39.600 301.600 40.400 302.400 ;
        RECT 39.700 298.400 40.300 301.600 ;
        RECT 39.600 297.600 40.400 298.400 ;
        RECT 41.300 296.400 41.900 309.600 ;
        RECT 42.900 308.400 43.500 311.600 ;
        RECT 44.500 310.400 45.100 311.600 ;
        RECT 47.700 310.400 48.300 315.600 ;
        RECT 57.200 313.600 58.000 314.400 ;
        RECT 54.000 311.600 54.800 312.400 ;
        RECT 55.600 311.600 56.400 312.400 ;
        RECT 44.400 309.600 45.200 310.400 ;
        RECT 47.600 309.600 48.400 310.400 ;
        RECT 44.500 308.400 45.100 309.600 ;
        RECT 42.800 307.600 43.600 308.400 ;
        RECT 44.400 307.600 45.200 308.400 ;
        RECT 49.200 307.600 50.000 308.400 ;
        RECT 50.800 307.600 51.600 308.400 ;
        RECT 42.800 299.600 43.600 300.400 ;
        RECT 41.200 295.600 42.000 296.400 ;
        RECT 36.400 291.600 37.200 292.400 ;
        RECT 38.000 291.600 38.800 292.400 ;
        RECT 34.800 287.600 35.600 288.400 ;
        RECT 34.900 268.300 35.500 287.600 ;
        RECT 36.400 283.600 37.200 284.400 ;
        RECT 39.600 283.600 40.400 284.400 ;
        RECT 36.500 272.400 37.100 283.600 ;
        RECT 38.000 273.600 38.800 274.400 ;
        RECT 36.400 271.600 37.200 272.400 ;
        RECT 38.000 269.600 38.800 270.400 ;
        RECT 36.400 268.300 37.200 268.400 ;
        RECT 34.900 267.700 37.200 268.300 ;
        RECT 36.400 267.600 37.200 267.700 ;
        RECT 38.000 267.600 38.800 268.400 ;
        RECT 36.400 265.600 37.200 266.400 ;
        RECT 36.500 254.400 37.100 265.600 ;
        RECT 36.400 253.600 37.200 254.400 ;
        RECT 34.800 251.600 35.600 252.400 ;
        RECT 36.500 250.400 37.100 253.600 ;
        RECT 38.100 252.400 38.700 267.600 ;
        RECT 38.000 251.600 38.800 252.400 ;
        RECT 36.400 249.600 37.200 250.400 ;
        RECT 36.500 246.300 37.100 249.600 ;
        RECT 38.100 248.400 38.700 251.600 ;
        RECT 38.000 247.600 38.800 248.400 ;
        RECT 34.900 245.700 37.100 246.300 ;
        RECT 34.900 212.400 35.500 245.700 ;
        RECT 38.100 236.400 38.700 247.600 ;
        RECT 39.700 246.400 40.300 283.600 ;
        RECT 41.200 269.600 42.000 270.400 ;
        RECT 41.300 262.400 41.900 269.600 ;
        RECT 42.900 268.400 43.500 299.600 ;
        RECT 44.500 286.400 45.100 307.600 ;
        RECT 49.300 300.400 49.900 307.600 ;
        RECT 50.900 306.400 51.500 307.600 ;
        RECT 50.800 305.600 51.600 306.400 ;
        RECT 54.100 304.400 54.700 311.600 ;
        RECT 55.700 310.400 56.300 311.600 ;
        RECT 57.300 310.400 57.900 313.600 ;
        RECT 62.100 310.400 62.700 333.700 ;
        RECT 63.600 333.600 64.400 333.700 ;
        RECT 63.600 331.600 64.400 332.400 ;
        RECT 66.800 331.600 67.600 332.400 ;
        RECT 63.600 329.600 64.400 330.400 ;
        RECT 63.700 318.400 64.300 329.600 ;
        RECT 65.200 327.600 66.000 328.400 ;
        RECT 63.600 317.600 64.400 318.400 ;
        RECT 65.300 312.400 65.900 327.600 ;
        RECT 68.500 318.400 69.100 341.600 ;
        RECT 70.000 329.600 70.800 330.400 ;
        RECT 68.400 317.600 69.200 318.400 ;
        RECT 65.200 311.600 66.000 312.400 ;
        RECT 66.800 311.600 67.600 312.400 ;
        RECT 65.300 310.400 65.900 311.600 ;
        RECT 66.900 310.400 67.500 311.600 ;
        RECT 55.600 309.600 56.400 310.400 ;
        RECT 57.200 309.600 58.000 310.400 ;
        RECT 58.800 309.600 59.600 310.400 ;
        RECT 62.000 309.600 62.800 310.400 ;
        RECT 65.200 309.600 66.000 310.400 ;
        RECT 66.800 309.600 67.600 310.400 ;
        RECT 54.000 303.600 54.800 304.400 ;
        RECT 57.200 303.600 58.000 304.400 ;
        RECT 57.300 300.400 57.900 303.600 ;
        RECT 49.200 299.600 50.000 300.400 ;
        RECT 57.200 299.600 58.000 300.400 ;
        RECT 47.600 291.600 48.400 292.400 ;
        RECT 44.400 285.600 45.200 286.400 ;
        RECT 47.700 276.400 48.300 291.600 ;
        RECT 49.200 284.200 50.000 297.800 ;
        RECT 50.800 284.200 51.600 297.800 ;
        RECT 52.400 284.200 53.200 297.800 ;
        RECT 54.000 286.200 54.800 297.800 ;
        RECT 55.600 295.600 56.400 296.400 ;
        RECT 55.700 282.400 56.300 295.600 ;
        RECT 57.200 286.200 58.000 297.800 ;
        RECT 58.900 294.400 59.500 309.600 ;
        RECT 62.000 307.600 62.800 308.400 ;
        RECT 62.100 302.400 62.700 307.600 ;
        RECT 65.300 304.400 65.900 309.600 ;
        RECT 66.800 307.600 67.600 308.400 ;
        RECT 66.900 306.400 67.500 307.600 ;
        RECT 66.800 305.600 67.600 306.400 ;
        RECT 65.200 303.600 66.000 304.400 ;
        RECT 62.000 301.600 62.800 302.400 ;
        RECT 66.800 301.600 67.600 302.400 ;
        RECT 58.800 293.600 59.600 294.400 ;
        RECT 60.400 286.200 61.200 297.800 ;
        RECT 62.000 284.200 62.800 297.800 ;
        RECT 63.600 284.200 64.400 297.800 ;
        RECT 55.600 281.600 56.400 282.400 ;
        RECT 66.900 278.400 67.500 301.600 ;
        RECT 70.100 294.400 70.700 329.600 ;
        RECT 71.700 322.400 72.300 347.600 ;
        RECT 73.200 344.200 74.000 355.800 ;
        RECT 74.800 345.600 75.600 346.400 ;
        RECT 74.900 344.400 75.500 345.600 ;
        RECT 74.800 343.600 75.600 344.400 ;
        RECT 76.400 344.200 77.200 355.800 ;
        RECT 78.000 344.200 78.800 357.800 ;
        RECT 79.600 344.200 80.400 357.800 ;
        RECT 81.200 344.200 82.000 357.800 ;
        RECT 82.800 349.600 83.600 350.400 ;
        RECT 89.300 344.400 89.900 375.600 ;
        RECT 90.800 366.200 91.600 377.800 ;
        RECT 92.400 373.600 93.200 374.400 ;
        RECT 92.400 365.600 93.200 366.400 ;
        RECT 94.000 366.200 94.800 377.800 ;
        RECT 92.500 350.400 93.100 365.600 ;
        RECT 95.600 364.200 96.400 377.800 ;
        RECT 97.200 364.200 98.000 377.800 ;
        RECT 100.400 371.600 101.200 372.400 ;
        RECT 97.200 357.600 98.000 358.400 ;
        RECT 92.400 349.600 93.200 350.400 ;
        RECT 89.200 343.600 90.000 344.400 ;
        RECT 73.200 337.600 74.000 338.400 ;
        RECT 73.300 334.400 73.900 337.600 ;
        RECT 92.500 336.400 93.100 349.600 ;
        RECT 97.300 346.400 97.900 357.600 ;
        RECT 100.500 350.400 101.100 371.600 ;
        RECT 114.800 365.600 115.600 366.400 ;
        RECT 124.400 364.200 125.200 377.800 ;
        RECT 126.000 364.200 126.800 377.800 ;
        RECT 127.600 364.200 128.400 377.800 ;
        RECT 129.200 366.200 130.000 377.800 ;
        RECT 130.800 375.600 131.600 376.400 ;
        RECT 130.900 364.300 131.500 375.600 ;
        RECT 132.400 366.200 133.200 377.800 ;
        RECT 134.000 375.600 134.800 376.400 ;
        RECT 134.100 374.400 134.700 375.600 ;
        RECT 134.000 373.600 134.800 374.400 ;
        RECT 135.600 366.200 136.400 377.800 ;
        RECT 129.300 363.700 131.500 364.300 ;
        RECT 137.200 364.200 138.000 377.800 ;
        RECT 138.800 364.200 139.600 377.800 ;
        RECT 140.400 371.600 141.200 372.400 ;
        RECT 153.200 371.600 154.000 372.400 ;
        RECT 100.400 349.600 101.200 350.400 ;
        RECT 94.000 345.600 94.800 346.400 ;
        RECT 97.200 345.600 98.000 346.400 ;
        RECT 74.800 335.600 75.600 336.400 ;
        RECT 79.600 335.600 80.400 336.400 ;
        RECT 92.400 335.600 93.200 336.400 ;
        RECT 79.700 334.400 80.300 335.600 ;
        RECT 73.200 333.600 74.000 334.400 ;
        RECT 79.600 333.600 80.400 334.400 ;
        RECT 89.200 333.600 90.000 334.400 ;
        RECT 82.800 331.600 83.600 332.400 ;
        RECT 87.600 331.600 88.400 332.400 ;
        RECT 89.300 330.400 89.900 333.600 ;
        RECT 90.800 331.600 91.600 332.400 ;
        RECT 74.800 329.600 75.600 330.400 ;
        RECT 86.000 329.600 86.800 330.400 ;
        RECT 89.200 329.600 90.000 330.400 ;
        RECT 86.100 328.400 86.700 329.600 ;
        RECT 94.100 328.400 94.700 345.600 ;
        RECT 95.600 343.600 96.400 344.400 ;
        RECT 95.700 338.400 96.300 343.600 ;
        RECT 95.600 337.600 96.400 338.400 ;
        RECT 97.300 334.400 97.900 345.600 ;
        RECT 106.800 344.200 107.600 357.800 ;
        RECT 108.400 344.200 109.200 357.800 ;
        RECT 110.000 344.200 110.800 355.800 ;
        RECT 111.600 347.600 112.400 348.400 ;
        RECT 113.200 344.200 114.000 355.800 ;
        RECT 114.800 345.600 115.600 346.400 ;
        RECT 114.900 342.400 115.500 345.600 ;
        RECT 116.400 344.200 117.200 355.800 ;
        RECT 118.000 344.200 118.800 357.800 ;
        RECT 119.600 344.200 120.400 357.800 ;
        RECT 121.200 344.200 122.000 357.800 ;
        RECT 122.800 349.600 123.600 350.400 ;
        RECT 111.600 341.600 112.400 342.400 ;
        RECT 114.800 341.600 115.600 342.400 ;
        RECT 97.200 333.600 98.000 334.400 ;
        RECT 103.600 329.600 104.400 330.400 ;
        RECT 86.000 327.600 86.800 328.400 ;
        RECT 94.000 327.600 94.800 328.400 ;
        RECT 92.400 325.600 93.200 326.400 ;
        RECT 87.600 323.600 88.400 324.400 ;
        RECT 71.600 321.600 72.400 322.400 ;
        RECT 73.200 313.600 74.000 314.400 ;
        RECT 71.600 309.600 72.400 310.400 ;
        RECT 71.700 302.400 72.300 309.600 ;
        RECT 73.300 308.400 73.900 313.600 ;
        RECT 73.200 307.600 74.000 308.400 ;
        RECT 87.700 306.400 88.300 323.600 ;
        RECT 92.500 310.400 93.100 325.600 ;
        RECT 95.600 323.600 96.400 324.400 ;
        RECT 95.700 312.400 96.300 323.600 ;
        RECT 94.000 311.600 94.800 312.400 ;
        RECT 95.600 311.600 96.400 312.400 ;
        RECT 98.800 311.600 99.600 312.400 ;
        RECT 92.400 309.600 93.200 310.400 ;
        RECT 90.800 307.600 91.600 308.400 ;
        RECT 92.400 307.600 93.200 308.400 ;
        RECT 74.800 305.600 75.600 306.400 ;
        RECT 76.400 305.600 77.200 306.400 ;
        RECT 79.600 305.600 80.400 306.400 ;
        RECT 87.600 305.600 88.400 306.400 ;
        RECT 74.900 304.400 75.500 305.600 ;
        RECT 74.800 303.600 75.600 304.400 ;
        RECT 71.600 301.600 72.400 302.400 ;
        RECT 70.000 293.600 70.800 294.400 ;
        RECT 68.400 291.600 69.200 292.400 ;
        RECT 74.800 283.600 75.600 284.400 ;
        RECT 66.800 277.600 67.600 278.400 ;
        RECT 47.600 275.600 48.400 276.400 ;
        RECT 44.400 271.600 45.200 272.400 ;
        RECT 47.600 271.600 48.400 272.400 ;
        RECT 60.400 271.600 61.200 272.400 ;
        RECT 65.200 271.600 66.000 272.400 ;
        RECT 70.000 271.600 70.800 272.400 ;
        RECT 42.800 267.600 43.600 268.400 ;
        RECT 41.200 261.600 42.000 262.400 ;
        RECT 42.900 258.400 43.500 267.600 ;
        RECT 44.500 266.400 45.100 271.600 ;
        RECT 47.700 268.400 48.300 271.600 ;
        RECT 79.700 270.400 80.300 305.600 ;
        RECT 82.800 291.600 83.600 292.400 ;
        RECT 84.400 284.200 85.200 297.800 ;
        RECT 86.000 284.200 86.800 297.800 ;
        RECT 87.600 284.200 88.400 297.800 ;
        RECT 89.200 286.200 90.000 297.800 ;
        RECT 90.900 296.400 91.500 307.600 ;
        RECT 92.500 306.400 93.100 307.600 ;
        RECT 92.400 305.600 93.200 306.400 ;
        RECT 90.800 295.600 91.600 296.400 ;
        RECT 49.200 269.600 50.000 270.400 ;
        RECT 52.400 269.600 53.200 270.400 ;
        RECT 55.600 269.600 56.400 270.400 ;
        RECT 63.600 269.600 64.400 270.400 ;
        RECT 73.200 269.600 74.000 270.400 ;
        RECT 79.600 269.600 80.400 270.400 ;
        RECT 82.800 269.600 83.600 270.400 ;
        RECT 86.000 269.600 86.800 270.400 ;
        RECT 49.300 268.400 49.900 269.600 ;
        RECT 63.700 268.400 64.300 269.600 ;
        RECT 47.600 267.600 48.400 268.400 ;
        RECT 49.200 267.600 50.000 268.400 ;
        RECT 54.000 267.600 54.800 268.400 ;
        RECT 60.400 267.600 61.200 268.400 ;
        RECT 63.600 267.600 64.400 268.400 ;
        RECT 68.400 267.600 69.200 268.400 ;
        RECT 74.800 267.600 75.600 268.400 ;
        RECT 44.400 265.600 45.200 266.400 ;
        RECT 52.400 265.600 53.200 266.400 ;
        RECT 55.600 265.600 56.400 266.400 ;
        RECT 52.500 264.400 53.100 265.600 ;
        RECT 46.000 263.600 46.800 264.400 ;
        RECT 52.400 263.600 53.200 264.400 ;
        RECT 42.800 257.600 43.600 258.400 ;
        RECT 46.100 256.400 46.700 263.600 ;
        RECT 41.200 255.600 42.000 256.400 ;
        RECT 44.400 255.600 45.200 256.400 ;
        RECT 46.000 255.600 46.800 256.400 ;
        RECT 42.800 253.600 43.600 254.400 ;
        RECT 54.000 253.600 54.800 254.400 ;
        RECT 39.600 245.600 40.400 246.400 ;
        RECT 41.200 245.600 42.000 246.400 ;
        RECT 39.600 243.600 40.400 244.400 ;
        RECT 39.700 238.400 40.300 243.600 ;
        RECT 41.300 238.400 41.900 245.600 ;
        RECT 39.600 237.600 40.400 238.400 ;
        RECT 41.200 237.600 42.000 238.400 ;
        RECT 38.000 235.600 38.800 236.400 ;
        RECT 38.000 233.600 38.800 234.400 ;
        RECT 39.600 233.600 40.400 234.400 ;
        RECT 36.400 231.600 37.200 232.400 ;
        RECT 36.500 230.400 37.100 231.600 ;
        RECT 38.100 230.400 38.700 233.600 ;
        RECT 36.400 229.600 37.200 230.400 ;
        RECT 38.000 229.600 38.800 230.400 ;
        RECT 38.100 216.400 38.700 229.600 ;
        RECT 39.700 228.400 40.300 233.600 ;
        RECT 42.900 228.400 43.500 253.600 ;
        RECT 49.200 251.600 50.000 252.400 ;
        RECT 46.000 249.600 46.800 250.400 ;
        RECT 47.600 249.600 48.400 250.400 ;
        RECT 46.100 248.400 46.700 249.600 ;
        RECT 46.000 247.600 46.800 248.400 ;
        RECT 47.700 246.400 48.300 249.600 ;
        RECT 47.600 245.600 48.400 246.400 ;
        RECT 49.300 242.400 49.900 251.600 ;
        RECT 50.800 249.600 51.600 250.400 ;
        RECT 50.900 248.400 51.500 249.600 ;
        RECT 50.800 247.600 51.600 248.400 ;
        RECT 52.400 243.600 53.200 244.400 ;
        RECT 55.700 244.300 56.300 265.600 ;
        RECT 57.200 263.600 58.000 264.400 ;
        RECT 57.300 258.400 57.900 263.600 ;
        RECT 57.200 257.600 58.000 258.400 ;
        RECT 57.200 249.600 58.000 250.400 ;
        RECT 58.800 249.600 59.600 250.400 ;
        RECT 57.300 246.400 57.900 249.600 ;
        RECT 57.200 245.600 58.000 246.400 ;
        RECT 58.800 245.600 59.600 246.400 ;
        RECT 55.700 243.700 57.900 244.300 ;
        RECT 46.000 241.600 46.800 242.400 ;
        RECT 49.200 241.600 50.000 242.400 ;
        RECT 44.400 231.600 45.200 232.400 ;
        RECT 44.400 229.600 45.200 230.400 ;
        RECT 39.600 227.600 40.400 228.400 ;
        RECT 42.800 227.600 43.600 228.400 ;
        RECT 39.600 223.600 40.400 224.400 ;
        RECT 38.000 215.600 38.800 216.400 ;
        RECT 39.700 214.400 40.300 223.600 ;
        RECT 42.900 222.400 43.500 227.600 ;
        RECT 42.800 221.600 43.600 222.400 ;
        RECT 36.400 213.600 37.200 214.400 ;
        RECT 39.600 213.600 40.400 214.400 ;
        RECT 44.500 212.400 45.100 229.600 ;
        RECT 46.100 212.400 46.700 241.600 ;
        RECT 49.200 239.600 50.000 240.400 ;
        RECT 47.600 229.600 48.400 230.400 ;
        RECT 49.300 228.400 49.900 239.600 ;
        RECT 52.500 236.400 53.100 243.600 ;
        RECT 50.800 235.600 51.600 236.400 ;
        RECT 52.400 235.600 53.200 236.400 ;
        RECT 50.900 230.400 51.500 235.600 ;
        RECT 50.800 229.600 51.600 230.400 ;
        RECT 49.200 227.600 50.000 228.400 ;
        RECT 50.800 227.600 51.600 228.400 ;
        RECT 34.800 211.600 35.600 212.400 ;
        RECT 38.000 211.600 38.800 212.400 ;
        RECT 39.600 211.600 40.400 212.400 ;
        RECT 44.400 211.600 45.200 212.400 ;
        RECT 46.000 211.600 46.800 212.400 ;
        RECT 47.600 211.600 48.400 212.400 ;
        RECT 38.100 210.400 38.700 211.600 ;
        RECT 38.000 209.600 38.800 210.400 ;
        RECT 38.100 204.400 38.700 209.600 ;
        RECT 38.000 203.600 38.800 204.400 ;
        RECT 33.200 199.600 34.000 200.400 ;
        RECT 31.600 195.600 32.400 196.400 ;
        RECT 31.600 193.600 32.400 194.400 ;
        RECT 36.400 193.600 37.200 194.400 ;
        RECT 22.000 189.600 22.800 190.400 ;
        RECT 25.200 189.600 26.000 190.400 ;
        RECT 17.200 187.600 18.000 188.800 ;
        RECT 14.000 171.700 16.300 172.300 ;
        RECT 14.000 171.600 14.800 171.700 ;
        RECT 14.100 152.400 14.700 171.600 ;
        RECT 15.600 169.600 16.400 170.400 ;
        RECT 14.000 151.600 14.800 152.400 ;
        RECT 17.300 150.400 17.900 187.600 ;
        RECT 22.000 185.600 22.800 186.400 ;
        RECT 20.400 183.600 21.200 184.400 ;
        RECT 20.500 180.400 21.100 183.600 ;
        RECT 20.400 179.600 21.200 180.400 ;
        RECT 25.300 180.300 25.900 189.600 ;
        RECT 26.800 187.600 27.600 188.400 ;
        RECT 28.400 187.600 29.200 188.400 ;
        RECT 26.900 186.400 27.500 187.600 ;
        RECT 26.800 185.600 27.600 186.400 ;
        RECT 28.500 182.400 29.100 187.600 ;
        RECT 28.400 181.600 29.200 182.400 ;
        RECT 23.700 179.700 25.900 180.300 ;
        RECT 23.700 178.400 24.300 179.700 ;
        RECT 28.400 179.600 29.200 180.400 ;
        RECT 23.600 177.600 24.400 178.400 ;
        RECT 23.700 176.400 24.300 177.600 ;
        RECT 18.800 175.600 19.600 176.400 ;
        RECT 22.000 175.600 22.800 176.400 ;
        RECT 23.600 175.600 24.400 176.400 ;
        RECT 18.900 172.300 19.500 175.600 ;
        RECT 20.400 173.600 21.200 174.400 ;
        RECT 28.500 172.400 29.100 179.600 ;
        RECT 30.000 173.600 30.800 174.400 ;
        RECT 18.900 171.700 21.100 172.300 ;
        RECT 18.800 151.600 19.600 152.400 ;
        RECT 18.900 150.400 19.500 151.600 ;
        RECT 17.200 149.600 18.000 150.400 ;
        RECT 18.800 149.600 19.600 150.400 ;
        RECT 20.500 148.400 21.100 171.700 ;
        RECT 28.400 171.600 29.200 172.400 ;
        RECT 30.100 170.400 30.700 173.600 ;
        RECT 30.000 169.600 30.800 170.400 ;
        RECT 31.700 168.400 32.300 193.600 ;
        RECT 33.200 191.600 34.000 192.400 ;
        RECT 34.800 191.600 35.600 192.400 ;
        RECT 33.300 186.300 33.900 191.600 ;
        RECT 34.900 190.400 35.500 191.600 ;
        RECT 34.800 189.600 35.600 190.400 ;
        RECT 34.800 187.600 35.600 188.400 ;
        RECT 33.300 185.700 35.500 186.300 ;
        RECT 33.200 171.600 34.000 172.400 ;
        RECT 30.000 167.600 30.800 168.400 ;
        RECT 31.600 167.600 32.400 168.400 ;
        RECT 28.400 163.600 29.200 164.400 ;
        RECT 25.200 153.600 26.000 154.400 ;
        RECT 20.400 147.600 21.200 148.400 ;
        RECT 20.500 146.400 21.100 147.600 ;
        RECT 25.300 146.400 25.900 153.600 ;
        RECT 28.400 149.600 29.200 150.400 ;
        RECT 20.400 145.600 21.200 146.400 ;
        RECT 25.200 145.600 26.000 146.400 ;
        RECT 28.400 145.600 29.200 146.400 ;
        RECT 20.400 143.600 21.200 144.400 ;
        RECT 12.400 141.600 13.200 142.400 ;
        RECT 20.500 142.300 21.100 143.600 ;
        RECT 28.500 142.400 29.100 145.600 ;
        RECT 20.500 141.700 22.700 142.300 ;
        RECT 12.500 136.400 13.100 141.600 ;
        RECT 20.400 139.600 21.200 140.400 ;
        RECT 12.400 135.600 13.200 136.400 ;
        RECT 15.600 135.600 16.400 136.400 ;
        RECT 15.700 132.400 16.300 135.600 ;
        RECT 20.500 134.400 21.100 139.600 ;
        RECT 17.200 133.600 18.000 134.400 ;
        RECT 18.800 133.600 19.600 134.400 ;
        RECT 20.400 133.600 21.200 134.400 ;
        RECT 17.300 132.400 17.900 133.600 ;
        RECT 18.900 132.400 19.500 133.600 ;
        RECT 15.600 131.600 16.400 132.400 ;
        RECT 17.200 131.600 18.000 132.400 ;
        RECT 18.800 131.600 19.600 132.400 ;
        RECT 22.100 130.400 22.700 141.700 ;
        RECT 28.400 141.600 29.200 142.400 ;
        RECT 26.800 131.600 27.600 132.400 ;
        RECT 28.400 131.600 29.200 132.400 ;
        RECT 28.500 130.400 29.100 131.600 ;
        RECT 9.300 129.700 11.500 130.300 ;
        RECT 1.200 123.600 2.000 124.400 ;
        RECT 1.300 94.400 1.900 123.600 ;
        RECT 4.400 121.600 5.200 122.400 ;
        RECT 4.500 118.400 5.100 121.600 ;
        RECT 9.300 118.400 9.900 129.700 ;
        RECT 22.000 129.600 22.800 130.400 ;
        RECT 28.400 129.600 29.200 130.400 ;
        RECT 22.100 128.400 22.700 129.600 ;
        RECT 22.000 127.600 22.800 128.400 ;
        RECT 25.200 127.600 26.000 128.400 ;
        RECT 22.000 125.600 22.800 126.400 ;
        RECT 22.100 118.400 22.700 125.600 ;
        RECT 26.800 123.600 27.600 124.400 ;
        RECT 30.100 124.300 30.700 167.600 ;
        RECT 34.900 164.400 35.500 185.700 ;
        RECT 36.500 178.400 37.100 193.600 ;
        RECT 36.400 177.600 37.200 178.400 ;
        RECT 36.500 174.400 37.100 177.600 ;
        RECT 38.000 175.600 38.800 176.400 ;
        RECT 38.100 174.400 38.700 175.600 ;
        RECT 36.400 173.600 37.200 174.400 ;
        RECT 38.000 173.600 38.800 174.400 ;
        RECT 39.700 172.400 40.300 211.600 ;
        RECT 47.700 210.400 48.300 211.600 ;
        RECT 46.000 209.600 46.800 210.400 ;
        RECT 47.600 209.600 48.400 210.400 ;
        RECT 44.400 208.300 45.200 208.400 ;
        RECT 42.900 207.700 45.200 208.300 ;
        RECT 42.900 206.400 43.500 207.700 ;
        RECT 44.400 207.600 45.200 207.700 ;
        RECT 42.800 205.600 43.600 206.400 ;
        RECT 44.400 205.600 45.200 206.400 ;
        RECT 41.200 203.600 42.000 204.400 ;
        RECT 41.300 194.400 41.900 203.600 ;
        RECT 42.800 201.600 43.600 202.400 ;
        RECT 42.900 198.400 43.500 201.600 ;
        RECT 42.800 197.600 43.600 198.400 ;
        RECT 41.200 193.600 42.000 194.400 ;
        RECT 44.500 192.400 45.100 205.600 ;
        RECT 46.100 204.400 46.700 209.600 ;
        RECT 46.000 203.600 46.800 204.400 ;
        RECT 44.400 191.600 45.200 192.400 ;
        RECT 42.800 190.300 43.600 190.400 ;
        RECT 41.300 189.700 43.600 190.300 ;
        RECT 39.600 172.300 40.400 172.400 ;
        RECT 38.100 171.700 40.400 172.300 ;
        RECT 34.800 163.600 35.600 164.400 ;
        RECT 36.400 153.600 37.200 154.400 ;
        RECT 36.400 151.600 37.200 152.400 ;
        RECT 36.500 150.400 37.100 151.600 ;
        RECT 31.600 149.600 32.400 150.400 ;
        RECT 36.400 149.600 37.200 150.400 ;
        RECT 31.700 146.400 32.300 149.600 ;
        RECT 31.600 145.600 32.400 146.400 ;
        RECT 33.200 145.600 34.000 146.400 ;
        RECT 36.400 145.600 37.200 146.400 ;
        RECT 33.300 138.400 33.900 145.600 ;
        RECT 33.200 137.600 34.000 138.400 ;
        RECT 36.500 136.400 37.100 145.600 ;
        RECT 36.400 135.600 37.200 136.400 ;
        RECT 36.500 134.400 37.100 135.600 ;
        RECT 33.200 133.600 34.000 134.400 ;
        RECT 36.400 133.600 37.200 134.400 ;
        RECT 33.300 132.400 33.900 133.600 ;
        RECT 38.100 132.400 38.700 171.700 ;
        RECT 39.600 171.600 40.400 171.700 ;
        RECT 41.300 166.400 41.900 189.700 ;
        RECT 42.800 189.600 43.600 189.700 ;
        RECT 46.100 186.400 46.700 203.600 ;
        RECT 49.300 200.300 49.900 227.600 ;
        RECT 54.000 225.600 54.800 226.400 ;
        RECT 55.600 223.600 56.400 224.400 ;
        RECT 55.700 220.400 56.300 223.600 ;
        RECT 55.600 219.600 56.400 220.400 ;
        RECT 57.300 218.400 57.900 243.700 ;
        RECT 58.900 230.400 59.500 245.600 ;
        RECT 60.500 234.400 61.100 267.600 ;
        RECT 68.400 265.600 69.200 266.400 ;
        RECT 74.800 265.600 75.600 266.400 ;
        RECT 76.400 265.600 77.200 266.400 ;
        RECT 62.000 263.600 62.800 264.400 ;
        RECT 62.100 262.400 62.700 263.600 ;
        RECT 62.000 261.600 62.800 262.400 ;
        RECT 63.600 255.600 64.400 256.400 ;
        RECT 68.500 252.400 69.100 265.600 ;
        RECT 70.000 263.600 70.800 264.400 ;
        RECT 70.100 254.400 70.700 263.600 ;
        RECT 73.200 257.600 74.000 258.400 ;
        RECT 73.300 254.400 73.900 257.600 ;
        RECT 74.900 256.400 75.500 265.600 ;
        RECT 76.500 256.400 77.100 265.600 ;
        RECT 74.800 255.600 75.600 256.400 ;
        RECT 76.400 255.600 77.200 256.400 ;
        RECT 81.200 256.300 82.000 256.400 ;
        RECT 82.900 256.300 83.500 269.600 ;
        RECT 86.100 268.400 86.700 269.600 ;
        RECT 86.000 267.600 86.800 268.400 ;
        RECT 87.600 265.600 88.400 266.400 ;
        RECT 89.200 263.600 90.000 264.400 ;
        RECT 81.200 255.700 83.500 256.300 ;
        RECT 81.200 255.600 82.000 255.700 ;
        RECT 70.000 253.600 70.800 254.400 ;
        RECT 73.200 253.600 74.000 254.400 ;
        RECT 74.800 253.600 75.600 254.400 ;
        RECT 63.600 251.600 64.400 252.400 ;
        RECT 66.800 251.600 67.600 252.400 ;
        RECT 68.400 251.600 69.200 252.400 ;
        RECT 70.000 251.600 70.800 252.400 ;
        RECT 71.600 251.600 72.400 252.400 ;
        RECT 66.900 250.300 67.500 251.600 ;
        RECT 68.400 250.300 69.200 250.400 ;
        RECT 66.900 249.700 69.200 250.300 ;
        RECT 68.400 249.600 69.200 249.700 ;
        RECT 65.200 247.600 66.000 248.400 ;
        RECT 62.000 245.600 62.800 246.400 ;
        RECT 60.400 233.600 61.200 234.400 ;
        RECT 62.100 232.400 62.700 245.600 ;
        RECT 65.300 244.400 65.900 247.600 ;
        RECT 65.200 243.600 66.000 244.400 ;
        RECT 62.000 231.600 62.800 232.400 ;
        RECT 65.300 230.400 65.900 243.600 ;
        RECT 70.000 237.600 70.800 238.400 ;
        RECT 68.400 233.600 69.200 234.400 ;
        RECT 70.100 230.400 70.700 237.600 ;
        RECT 71.700 234.400 72.300 251.600 ;
        RECT 73.300 240.400 73.900 253.600 ;
        RECT 73.200 239.600 74.000 240.400 ;
        RECT 74.900 240.300 75.500 253.600 ;
        RECT 79.600 251.600 80.400 252.400 ;
        RECT 76.400 245.600 77.200 246.400 ;
        RECT 74.900 239.700 77.100 240.300 ;
        RECT 74.800 237.600 75.600 238.400 ;
        RECT 71.600 233.600 72.400 234.400 ;
        RECT 73.200 233.600 74.000 234.400 ;
        RECT 71.600 231.600 72.400 232.400 ;
        RECT 58.800 229.600 59.600 230.400 ;
        RECT 60.400 229.600 61.200 230.400 ;
        RECT 65.200 229.600 66.000 230.400 ;
        RECT 70.000 229.600 70.800 230.400 ;
        RECT 60.500 228.400 61.100 229.600 ;
        RECT 65.300 228.400 65.900 229.600 ;
        RECT 73.300 228.400 73.900 233.600 ;
        RECT 74.900 230.400 75.500 237.600 ;
        RECT 74.800 229.600 75.600 230.400 ;
        RECT 60.400 227.600 61.200 228.400 ;
        RECT 65.200 227.600 66.000 228.400 ;
        RECT 73.200 227.600 74.000 228.400 ;
        RECT 62.000 225.600 62.800 226.400 ;
        RECT 66.800 223.600 67.600 224.400 ;
        RECT 57.200 217.600 58.000 218.400 ;
        RECT 65.200 217.600 66.000 218.400 ;
        RECT 50.800 215.600 51.600 216.400 ;
        RECT 50.900 202.400 51.500 215.600 ;
        RECT 52.400 213.600 53.200 214.400 ;
        RECT 63.600 213.600 64.400 214.400 ;
        RECT 52.500 210.400 53.100 213.600 ;
        RECT 63.700 212.400 64.300 213.600 ;
        RECT 54.000 211.600 54.800 212.400 ;
        RECT 63.600 211.600 64.400 212.400 ;
        RECT 52.400 209.600 53.200 210.400 ;
        RECT 50.800 201.600 51.600 202.400 ;
        RECT 47.700 199.700 49.900 200.300 ;
        RECT 47.700 186.400 48.300 199.700 ;
        RECT 54.100 196.400 54.700 211.600 ;
        RECT 62.000 209.600 62.800 210.400 ;
        RECT 62.100 208.400 62.700 209.600 ;
        RECT 62.000 207.600 62.800 208.400 ;
        RECT 63.700 206.400 64.300 211.600 ;
        RECT 65.300 208.400 65.900 217.600 ;
        RECT 65.200 207.600 66.000 208.400 ;
        RECT 63.600 205.600 64.400 206.400 ;
        RECT 63.600 203.600 64.400 204.400 ;
        RECT 63.700 202.400 64.300 203.600 ;
        RECT 60.400 201.600 61.200 202.400 ;
        RECT 63.600 201.600 64.400 202.400 ;
        RECT 57.200 197.600 58.000 198.400 ;
        RECT 54.000 195.600 54.800 196.400 ;
        RECT 52.400 193.600 53.200 194.400 ;
        RECT 55.600 193.600 56.400 194.400 ;
        RECT 52.500 192.400 53.100 193.600 ;
        RECT 52.400 191.600 53.200 192.400 ;
        RECT 49.200 189.600 50.000 190.400 ;
        RECT 49.300 188.400 49.900 189.600 ;
        RECT 49.200 187.600 50.000 188.400 ;
        RECT 44.400 185.600 45.200 186.400 ;
        RECT 46.000 185.600 46.800 186.400 ;
        RECT 47.600 185.600 48.400 186.400 ;
        RECT 49.200 185.600 50.000 186.400 ;
        RECT 42.800 175.600 43.600 176.400 ;
        RECT 44.500 174.400 45.100 185.600 ;
        RECT 47.600 183.600 48.400 184.400 ;
        RECT 42.800 173.600 43.600 174.400 ;
        RECT 44.400 173.600 45.200 174.400 ;
        RECT 46.000 173.600 46.800 174.400 ;
        RECT 42.900 172.400 43.500 173.600 ;
        RECT 42.800 171.600 43.600 172.400 ;
        RECT 42.800 167.600 43.600 168.400 ;
        RECT 41.200 165.600 42.000 166.400 ;
        RECT 42.900 158.400 43.500 167.600 ;
        RECT 44.500 162.400 45.100 173.600 ;
        RECT 46.100 172.400 46.700 173.600 ;
        RECT 46.000 171.600 46.800 172.400 ;
        RECT 44.400 161.600 45.200 162.400 ;
        RECT 42.800 157.600 43.600 158.400 ;
        RECT 42.800 155.600 43.600 156.400 ;
        RECT 41.200 147.600 42.000 148.400 ;
        RECT 39.600 145.600 40.400 146.400 ;
        RECT 41.200 133.600 42.000 134.400 ;
        RECT 33.200 131.600 34.000 132.400 ;
        RECT 34.800 131.600 35.600 132.400 ;
        RECT 38.000 132.300 38.800 132.400 ;
        RECT 36.500 131.700 38.800 132.300 ;
        RECT 34.900 130.400 35.500 131.600 ;
        RECT 34.800 129.600 35.600 130.400 ;
        RECT 31.600 127.600 32.400 128.400 ;
        RECT 33.200 127.600 34.000 128.400 ;
        RECT 33.300 126.400 33.900 127.600 ;
        RECT 33.200 125.600 34.000 126.400 ;
        RECT 28.500 123.700 30.700 124.300 ;
        RECT 4.400 117.600 5.200 118.400 ;
        RECT 9.200 117.600 10.000 118.400 ;
        RECT 22.000 117.600 22.800 118.400 ;
        RECT 15.600 115.600 16.400 116.400 ;
        RECT 20.400 115.600 21.200 116.400 ;
        RECT 20.500 114.400 21.100 115.600 ;
        RECT 6.000 113.600 6.800 114.400 ;
        RECT 14.000 113.600 14.800 114.400 ;
        RECT 18.800 113.600 19.600 114.400 ;
        RECT 20.400 113.600 21.200 114.400 ;
        RECT 6.100 112.400 6.700 113.600 ;
        RECT 4.400 111.600 5.200 112.400 ;
        RECT 6.000 111.600 6.800 112.400 ;
        RECT 10.800 111.600 11.600 112.400 ;
        RECT 17.200 111.600 18.000 112.400 ;
        RECT 4.400 110.300 5.200 110.400 ;
        RECT 2.900 109.700 5.200 110.300 ;
        RECT 1.200 93.600 2.000 94.400 ;
        RECT 1.300 90.400 1.900 93.600 ;
        RECT 1.200 89.600 2.000 90.400 ;
        RECT 2.900 78.400 3.500 109.700 ;
        RECT 4.400 109.600 5.200 109.700 ;
        RECT 4.500 108.400 5.100 109.600 ;
        RECT 4.400 107.600 5.200 108.400 ;
        RECT 4.400 89.600 5.200 90.400 ;
        RECT 4.500 88.400 5.100 89.600 ;
        RECT 4.400 87.600 5.200 88.400 ;
        RECT 2.800 77.600 3.600 78.400 ;
        RECT 4.400 69.600 5.200 70.400 ;
        RECT 1.200 65.600 2.000 66.400 ;
        RECT 2.800 65.600 3.600 66.400 ;
        RECT 1.300 56.400 1.900 65.600 ;
        RECT 4.500 56.400 5.100 69.600 ;
        RECT 6.100 68.400 6.700 111.600 ;
        RECT 14.000 109.600 14.800 110.400 ;
        RECT 15.600 109.600 16.400 110.400 ;
        RECT 7.600 107.600 8.400 108.400 ;
        RECT 9.200 103.600 10.000 104.400 ;
        RECT 9.300 96.400 9.900 103.600 ;
        RECT 14.100 98.400 14.700 109.600 ;
        RECT 14.000 97.600 14.800 98.400 ;
        RECT 9.200 95.600 10.000 96.400 ;
        RECT 14.000 95.600 14.800 96.400 ;
        RECT 14.100 92.400 14.700 95.600 ;
        RECT 15.700 94.400 16.300 109.600 ;
        RECT 15.600 93.600 16.400 94.400 ;
        RECT 14.000 91.600 14.800 92.400 ;
        RECT 12.400 87.600 13.200 88.400 ;
        RECT 7.600 83.600 8.400 84.400 ;
        RECT 10.800 83.600 11.600 84.400 ;
        RECT 7.700 74.400 8.300 83.600 ;
        RECT 7.600 73.600 8.400 74.400 ;
        RECT 9.200 69.600 10.000 70.400 ;
        RECT 6.000 67.600 6.800 68.400 ;
        RECT 6.100 66.400 6.700 67.600 ;
        RECT 6.000 65.600 6.800 66.400 ;
        RECT 9.200 66.300 10.000 66.400 ;
        RECT 7.700 65.700 10.000 66.300 ;
        RECT 7.700 58.400 8.300 65.700 ;
        RECT 9.200 65.600 10.000 65.700 ;
        RECT 10.900 58.400 11.500 83.600 ;
        RECT 12.400 69.600 13.200 70.400 ;
        RECT 14.100 68.400 14.700 91.600 ;
        RECT 17.300 90.400 17.900 111.600 ;
        RECT 15.600 89.600 16.400 90.400 ;
        RECT 17.200 89.600 18.000 90.400 ;
        RECT 18.900 88.400 19.500 113.600 ;
        RECT 26.900 112.400 27.500 123.600 ;
        RECT 28.500 114.400 29.100 123.700 ;
        RECT 30.000 121.600 30.800 122.400 ;
        RECT 30.100 118.400 30.700 121.600 ;
        RECT 30.000 117.600 30.800 118.400 ;
        RECT 28.400 113.600 29.200 114.400 ;
        RECT 23.600 111.600 24.400 112.400 ;
        RECT 25.200 111.600 26.000 112.400 ;
        RECT 26.800 111.600 27.600 112.400 ;
        RECT 31.600 111.600 32.400 112.400 ;
        RECT 22.000 109.600 22.800 110.400 ;
        RECT 23.700 100.300 24.300 111.600 ;
        RECT 36.500 110.400 37.100 131.700 ;
        RECT 38.000 131.600 38.800 131.700 ;
        RECT 38.000 129.600 38.800 130.400 ;
        RECT 41.200 129.600 42.000 130.400 ;
        RECT 26.800 109.600 27.600 110.400 ;
        RECT 36.400 109.600 37.200 110.400 ;
        RECT 23.700 99.700 25.900 100.300 ;
        RECT 23.600 95.600 24.400 96.400 ;
        RECT 23.700 94.400 24.300 95.600 ;
        RECT 23.600 93.600 24.400 94.400 ;
        RECT 20.400 91.600 21.200 92.400 ;
        RECT 23.600 91.600 24.400 92.400 ;
        RECT 23.700 90.400 24.300 91.600 ;
        RECT 22.000 89.600 22.800 90.400 ;
        RECT 23.600 89.600 24.400 90.400 ;
        RECT 18.800 87.600 19.600 88.400 ;
        RECT 20.400 87.600 21.200 88.400 ;
        RECT 20.500 84.400 21.100 87.600 ;
        RECT 20.400 83.600 21.200 84.400 ;
        RECT 15.600 81.600 16.400 82.400 ;
        RECT 15.700 78.400 16.300 81.600 ;
        RECT 15.600 77.600 16.400 78.400 ;
        RECT 14.000 67.600 14.800 68.400 ;
        RECT 17.200 66.300 18.000 66.400 ;
        RECT 15.700 65.700 18.000 66.300 ;
        RECT 15.700 58.400 16.300 65.700 ;
        RECT 17.200 65.600 18.000 65.700 ;
        RECT 18.800 65.600 19.600 66.400 ;
        RECT 7.600 57.600 8.400 58.400 ;
        RECT 10.800 57.600 11.600 58.400 ;
        RECT 15.600 57.600 16.400 58.400 ;
        RECT 20.500 56.400 21.100 83.600 ;
        RECT 23.700 78.400 24.300 89.600 ;
        RECT 25.300 88.400 25.900 99.700 ;
        RECT 26.900 92.400 27.500 109.600 ;
        RECT 33.200 107.600 34.000 108.400 ;
        RECT 36.400 107.600 37.200 108.400 ;
        RECT 33.300 106.400 33.900 107.600 ;
        RECT 33.200 105.600 34.000 106.400 ;
        RECT 31.600 101.600 32.400 102.400 ;
        RECT 28.400 97.600 29.200 98.400 ;
        RECT 26.800 91.600 27.600 92.400 ;
        RECT 25.200 87.600 26.000 88.400 ;
        RECT 26.900 78.400 27.500 91.600 ;
        RECT 28.500 90.400 29.100 97.600 ;
        RECT 30.000 93.600 30.800 94.400 ;
        RECT 30.000 91.600 30.800 92.400 ;
        RECT 28.400 89.600 29.200 90.400 ;
        RECT 30.100 88.400 30.700 91.600 ;
        RECT 30.000 87.600 30.800 88.400 ;
        RECT 23.600 77.600 24.400 78.400 ;
        RECT 26.800 77.600 27.600 78.400 ;
        RECT 31.700 70.400 32.300 101.600 ;
        RECT 33.200 97.600 34.000 98.400 ;
        RECT 33.300 90.400 33.900 97.600 ;
        RECT 33.200 89.600 34.000 90.400 ;
        RECT 36.500 72.400 37.100 107.600 ;
        RECT 38.100 98.400 38.700 129.600 ;
        RECT 41.300 128.400 41.900 129.600 ;
        RECT 41.200 127.600 42.000 128.400 ;
        RECT 41.200 107.600 42.000 108.400 ;
        RECT 39.600 103.600 40.400 104.400 ;
        RECT 38.000 97.600 38.800 98.400 ;
        RECT 39.700 96.400 40.300 103.600 ;
        RECT 39.600 95.600 40.400 96.400 ;
        RECT 42.900 94.400 43.500 155.600 ;
        RECT 44.400 153.600 45.200 154.400 ;
        RECT 44.500 152.400 45.100 153.600 ;
        RECT 44.400 151.600 45.200 152.400 ;
        RECT 44.400 147.600 45.200 148.400 ;
        RECT 44.500 130.400 45.100 147.600 ;
        RECT 47.700 134.300 48.300 183.600 ;
        RECT 49.300 178.400 49.900 185.600 ;
        RECT 52.400 183.600 53.200 184.400 ;
        RECT 55.700 182.400 56.300 193.600 ;
        RECT 58.800 191.600 59.600 192.400 ;
        RECT 57.200 189.600 58.000 190.400 ;
        RECT 57.300 186.400 57.900 189.600 ;
        RECT 60.500 188.400 61.100 201.600 ;
        RECT 62.000 199.600 62.800 200.400 ;
        RECT 63.600 199.600 64.400 200.400 ;
        RECT 62.100 190.400 62.700 199.600 ;
        RECT 62.000 189.600 62.800 190.400 ;
        RECT 60.400 187.600 61.200 188.400 ;
        RECT 57.200 185.600 58.000 186.400 ;
        RECT 52.400 181.600 53.200 182.400 ;
        RECT 55.600 181.600 56.400 182.400 ;
        RECT 52.500 178.400 53.100 181.600 ;
        RECT 54.000 179.600 54.800 180.400 ;
        RECT 49.200 177.600 50.000 178.400 ;
        RECT 52.400 177.600 53.200 178.400 ;
        RECT 54.100 174.400 54.700 179.600 ;
        RECT 57.200 177.600 58.000 178.400 ;
        RECT 54.000 173.600 54.800 174.400 ;
        RECT 49.200 169.600 50.000 170.400 ;
        RECT 58.800 163.600 59.600 164.400 ;
        RECT 57.200 161.600 58.000 162.400 ;
        RECT 49.200 159.600 50.000 160.400 ;
        RECT 49.300 146.400 49.900 159.600 ;
        RECT 50.800 153.600 51.600 154.400 ;
        RECT 50.900 150.400 51.500 153.600 ;
        RECT 52.400 151.600 53.200 152.400 ;
        RECT 50.800 149.600 51.600 150.400 ;
        RECT 49.200 145.600 50.000 146.400 ;
        RECT 50.800 145.600 51.600 146.400 ;
        RECT 49.200 143.600 50.000 144.400 ;
        RECT 46.100 133.700 48.300 134.300 ;
        RECT 46.100 132.400 46.700 133.700 ;
        RECT 46.000 131.600 46.800 132.400 ;
        RECT 44.400 129.600 45.200 130.400 ;
        RECT 47.600 129.600 48.400 130.400 ;
        RECT 49.300 128.400 49.900 143.600 ;
        RECT 50.900 138.400 51.500 145.600 ;
        RECT 50.800 137.600 51.600 138.400 ;
        RECT 49.200 127.600 50.000 128.400 ;
        RECT 46.000 123.600 46.800 124.400 ;
        RECT 44.400 103.600 45.200 104.400 ;
        RECT 44.500 102.400 45.100 103.600 ;
        RECT 44.400 101.600 45.200 102.400 ;
        RECT 46.100 98.400 46.700 123.600 ;
        RECT 52.500 108.400 53.100 151.600 ;
        RECT 57.300 148.400 57.900 161.600 ;
        RECT 58.900 150.400 59.500 163.600 ;
        RECT 60.500 154.400 61.100 187.600 ;
        RECT 60.400 153.600 61.200 154.400 ;
        RECT 58.800 149.600 59.600 150.400 ;
        RECT 62.100 148.400 62.700 189.600 ;
        RECT 63.700 156.400 64.300 199.600 ;
        RECT 66.900 192.400 67.500 223.600 ;
        RECT 68.400 217.600 69.200 218.400 ;
        RECT 68.500 210.400 69.100 217.600 ;
        RECT 76.500 212.400 77.100 239.700 ;
        RECT 78.000 233.600 78.800 234.400 ;
        RECT 79.700 230.400 80.300 251.600 ;
        RECT 84.400 233.600 85.200 234.400 ;
        RECT 87.600 233.600 88.400 234.400 ;
        RECT 82.800 231.600 83.600 232.400 ;
        RECT 79.600 229.600 80.400 230.400 ;
        RECT 82.900 228.400 83.500 231.600 ;
        RECT 84.500 230.400 85.100 233.600 ;
        RECT 84.400 229.600 85.200 230.400 ;
        RECT 86.000 229.600 86.800 230.400 ;
        RECT 82.800 227.600 83.600 228.400 ;
        RECT 86.100 226.400 86.700 229.600 ;
        RECT 79.600 225.600 80.400 226.400 ;
        RECT 86.000 225.600 86.800 226.400 ;
        RECT 79.700 224.400 80.300 225.600 ;
        RECT 79.600 223.600 80.400 224.400 ;
        RECT 81.200 223.600 82.000 224.400 ;
        RECT 86.000 223.600 86.800 224.400 ;
        RECT 78.000 217.600 78.800 218.400 ;
        RECT 70.000 211.600 70.800 212.400 ;
        RECT 76.400 211.600 77.200 212.400 ;
        RECT 68.400 209.600 69.200 210.400 ;
        RECT 70.100 200.400 70.700 211.600 ;
        RECT 71.600 209.600 72.400 210.400 ;
        RECT 74.800 209.600 75.600 210.400 ;
        RECT 71.700 208.400 72.300 209.600 ;
        RECT 71.600 207.600 72.400 208.400 ;
        RECT 74.900 204.400 75.500 209.600 ;
        RECT 78.100 208.400 78.700 217.600 ;
        RECT 81.300 210.400 81.900 223.600 ;
        RECT 86.100 218.400 86.700 223.600 ;
        RECT 86.000 217.600 86.800 218.400 ;
        RECT 82.800 213.600 83.600 214.400 ;
        RECT 81.200 209.600 82.000 210.400 ;
        RECT 78.000 207.600 78.800 208.400 ;
        RECT 73.200 203.600 74.000 204.400 ;
        RECT 74.800 203.600 75.600 204.400 ;
        RECT 73.300 200.400 73.900 203.600 ;
        RECT 70.000 199.600 70.800 200.400 ;
        RECT 73.200 199.600 74.000 200.400 ;
        RECT 82.900 198.400 83.500 213.600 ;
        RECT 87.700 212.400 88.300 233.600 ;
        RECT 89.300 230.400 89.900 263.600 ;
        RECT 90.900 260.400 91.500 295.600 ;
        RECT 92.400 286.200 93.200 297.800 ;
        RECT 94.100 294.400 94.700 311.600 ;
        RECT 98.900 310.400 99.500 311.600 ;
        RECT 98.800 309.600 99.600 310.400 ;
        RECT 103.700 308.400 104.300 329.600 ;
        RECT 105.200 324.200 106.000 337.800 ;
        RECT 106.800 324.200 107.600 337.800 ;
        RECT 108.400 324.200 109.200 337.800 ;
        RECT 110.000 326.200 110.800 337.800 ;
        RECT 111.700 336.400 112.300 341.600 ;
        RECT 111.600 335.600 112.400 336.400 ;
        RECT 111.600 327.600 112.400 328.400 ;
        RECT 106.800 321.600 107.600 322.400 ;
        RECT 105.200 313.600 106.000 314.400 ;
        RECT 102.000 307.600 102.800 308.400 ;
        RECT 103.600 307.600 104.400 308.400 ;
        RECT 94.000 293.600 94.800 294.400 ;
        RECT 95.600 286.200 96.400 297.800 ;
        RECT 97.200 284.200 98.000 297.800 ;
        RECT 98.800 284.200 99.600 297.800 ;
        RECT 102.100 284.400 102.700 307.600 ;
        RECT 106.900 296.300 107.500 321.600 ;
        RECT 108.400 311.600 109.200 312.400 ;
        RECT 110.000 311.600 110.800 312.400 ;
        RECT 108.500 306.400 109.100 311.600 ;
        RECT 111.700 306.400 112.300 327.600 ;
        RECT 113.200 326.200 114.000 337.800 ;
        RECT 114.800 333.600 115.600 334.400 ;
        RECT 114.900 330.400 115.500 333.600 ;
        RECT 114.800 329.600 115.600 330.400 ;
        RECT 116.400 326.200 117.200 337.800 ;
        RECT 118.000 324.200 118.800 337.800 ;
        RECT 119.600 324.200 120.400 337.800 ;
        RECT 122.900 332.400 123.500 349.600 ;
        RECT 129.300 342.400 129.900 363.700 ;
        RECT 140.500 350.400 141.100 371.600 ;
        RECT 140.400 349.600 141.200 350.400 ;
        RECT 143.600 349.600 144.400 350.400 ;
        RECT 130.800 343.600 131.600 344.400 ;
        RECT 129.200 341.600 130.000 342.400 ;
        RECT 122.800 331.600 123.600 332.400 ;
        RECT 129.200 311.600 130.000 312.400 ;
        RECT 114.800 309.600 115.600 310.400 ;
        RECT 121.200 309.600 122.000 310.400 ;
        RECT 119.600 307.600 120.400 308.400 ;
        RECT 108.400 305.600 109.200 306.400 ;
        RECT 111.600 305.600 112.400 306.400 ;
        RECT 118.000 305.600 118.800 306.400 ;
        RECT 108.500 298.400 109.100 305.600 ;
        RECT 108.400 297.600 109.200 298.400 ;
        RECT 108.400 296.300 109.200 296.400 ;
        RECT 106.900 295.700 109.200 296.300 ;
        RECT 108.400 295.600 109.200 295.700 ;
        RECT 118.100 294.400 118.700 305.600 ;
        RECT 119.700 300.400 120.300 307.600 ;
        RECT 122.800 305.600 123.600 306.400 ;
        RECT 119.600 299.600 120.400 300.400 ;
        RECT 119.600 297.600 120.400 298.400 ;
        RECT 119.700 296.400 120.300 297.600 ;
        RECT 119.600 295.600 120.400 296.400 ;
        RECT 118.000 293.600 118.800 294.400 ;
        RECT 122.900 292.400 123.500 305.600 ;
        RECT 126.000 303.600 126.800 304.400 ;
        RECT 126.100 292.400 126.700 303.600 ;
        RECT 129.300 294.400 129.900 311.600 ;
        RECT 130.900 304.400 131.500 343.600 ;
        RECT 140.500 332.400 141.100 349.600 ;
        RECT 148.400 344.200 149.200 357.800 ;
        RECT 150.000 344.200 150.800 357.800 ;
        RECT 151.600 344.200 152.400 355.800 ;
        RECT 153.300 350.400 153.900 371.600 ;
        RECT 156.400 364.200 157.200 377.800 ;
        RECT 158.000 364.200 158.800 377.800 ;
        RECT 159.600 366.200 160.400 377.800 ;
        RECT 161.200 373.600 162.000 374.400 ;
        RECT 161.300 372.400 161.900 373.600 ;
        RECT 161.200 371.600 162.000 372.400 ;
        RECT 162.800 366.200 163.600 377.800 ;
        RECT 164.400 375.600 165.200 376.400 ;
        RECT 153.200 349.600 154.000 350.400 ;
        RECT 153.200 347.600 154.000 348.400 ;
        RECT 151.600 341.600 152.400 342.400 ;
        RECT 140.400 331.600 141.200 332.400 ;
        RECT 140.400 329.600 141.200 330.400 ;
        RECT 140.500 318.400 141.100 329.600 ;
        RECT 143.600 324.200 144.400 337.800 ;
        RECT 145.200 324.200 146.000 337.800 ;
        RECT 146.800 326.200 147.600 337.800 ;
        RECT 148.400 333.600 149.200 334.400 ;
        RECT 148.500 318.400 149.100 333.600 ;
        RECT 150.000 326.200 150.800 337.800 ;
        RECT 151.700 336.400 152.300 341.600 ;
        RECT 153.300 340.400 153.900 347.600 ;
        RECT 154.800 344.200 155.600 355.800 ;
        RECT 156.400 345.600 157.200 346.400 ;
        RECT 156.500 342.400 157.100 345.600 ;
        RECT 158.000 344.200 158.800 355.800 ;
        RECT 159.600 344.200 160.400 357.800 ;
        RECT 161.200 344.200 162.000 357.800 ;
        RECT 162.800 344.200 163.600 357.800 ;
        RECT 164.500 342.400 165.100 375.600 ;
        RECT 166.000 366.200 166.800 377.800 ;
        RECT 167.600 364.200 168.400 377.800 ;
        RECT 169.200 364.200 170.000 377.800 ;
        RECT 170.800 364.200 171.600 377.800 ;
        RECT 172.400 371.600 173.200 372.400 ;
        RECT 175.600 371.600 176.400 372.400 ;
        RECT 186.800 371.600 187.600 372.400 ;
        RECT 172.500 370.400 173.100 371.600 ;
        RECT 172.400 369.600 173.200 370.400 ;
        RECT 170.800 347.600 171.600 348.400 ;
        RECT 156.400 341.600 157.200 342.400 ;
        RECT 164.400 341.600 165.200 342.400 ;
        RECT 153.200 339.600 154.000 340.400 ;
        RECT 151.600 335.600 152.400 336.400 ;
        RECT 151.700 322.400 152.300 335.600 ;
        RECT 153.200 326.200 154.000 337.800 ;
        RECT 154.800 324.200 155.600 337.800 ;
        RECT 156.400 324.200 157.200 337.800 ;
        RECT 158.000 324.200 158.800 337.800 ;
        RECT 159.600 333.600 160.400 334.400 ;
        RECT 169.200 333.600 170.000 334.400 ;
        RECT 159.700 332.400 160.300 333.600 ;
        RECT 159.600 331.600 160.400 332.400 ;
        RECT 167.600 323.600 168.400 324.400 ;
        RECT 151.600 321.600 152.400 322.400 ;
        RECT 156.400 321.600 157.200 322.400 ;
        RECT 156.500 318.400 157.100 321.600 ;
        RECT 167.700 320.400 168.300 323.600 ;
        RECT 159.600 319.600 160.400 320.400 ;
        RECT 167.600 319.600 168.400 320.400 ;
        RECT 140.400 317.600 141.200 318.400 ;
        RECT 148.400 317.600 149.200 318.400 ;
        RECT 156.400 317.600 157.200 318.400 ;
        RECT 134.000 313.600 134.800 314.400 ;
        RECT 140.400 313.600 141.200 314.400 ;
        RECT 130.800 303.600 131.600 304.400 ;
        RECT 134.100 300.400 134.700 313.600 ;
        RECT 137.200 311.600 138.000 312.400 ;
        RECT 140.500 310.400 141.100 313.600 ;
        RECT 143.600 311.600 144.400 312.400 ;
        RECT 135.600 309.600 136.400 310.400 ;
        RECT 140.400 309.600 141.200 310.400 ;
        RECT 135.600 305.600 136.400 306.400 ;
        RECT 135.700 304.400 136.300 305.600 ;
        RECT 135.600 303.600 136.400 304.400 ;
        RECT 134.000 299.600 134.800 300.400 ;
        RECT 135.700 296.300 136.300 303.600 ;
        RECT 137.200 296.300 138.000 296.400 ;
        RECT 135.700 295.700 138.000 296.300 ;
        RECT 137.200 295.600 138.000 295.700 ;
        RECT 143.700 294.400 144.300 311.600 ;
        RECT 159.700 310.400 160.300 319.600 ;
        RECT 167.600 317.600 168.400 318.400 ;
        RECT 166.000 311.600 166.800 312.400 ;
        RECT 159.600 309.600 160.400 310.400 ;
        RECT 164.400 309.600 165.200 310.400 ;
        RECT 156.400 303.600 157.200 304.400 ;
        RECT 156.500 296.400 157.100 303.600 ;
        RECT 156.400 295.600 157.200 296.400 ;
        RECT 159.700 294.400 160.300 309.600 ;
        RECT 161.200 307.600 162.000 308.400 ;
        RECT 161.300 306.400 161.900 307.600 ;
        RECT 161.200 305.600 162.000 306.400 ;
        RECT 164.400 306.300 165.200 306.400 ;
        RECT 162.900 305.700 165.200 306.300 ;
        RECT 129.200 293.600 130.000 294.400 ;
        RECT 143.600 293.600 144.400 294.400 ;
        RECT 153.200 293.600 154.000 294.400 ;
        RECT 158.000 293.600 158.800 294.400 ;
        RECT 159.600 293.600 160.400 294.400 ;
        RECT 153.300 292.400 153.900 293.600 ;
        RECT 103.600 291.600 104.400 292.400 ;
        RECT 116.400 291.600 117.200 292.400 ;
        RECT 122.800 291.600 123.600 292.400 ;
        RECT 126.000 291.600 126.800 292.400 ;
        RECT 137.200 291.600 138.000 292.400 ;
        RECT 142.000 291.600 142.800 292.400 ;
        RECT 150.000 291.600 150.800 292.400 ;
        RECT 153.200 291.600 154.000 292.400 ;
        RECT 154.800 291.600 155.600 292.400 ;
        RECT 159.600 292.300 160.400 292.400 ;
        RECT 161.300 292.300 161.900 305.600 ;
        RECT 162.900 298.400 163.500 305.700 ;
        RECT 164.400 305.600 165.200 305.700 ;
        RECT 166.100 298.400 166.700 311.600 ;
        RECT 167.700 310.400 168.300 317.600 ;
        RECT 170.900 310.400 171.500 347.600 ;
        RECT 172.400 343.600 173.200 344.400 ;
        RECT 172.500 318.400 173.100 343.600 ;
        RECT 175.700 338.400 176.300 371.600 ;
        RECT 186.900 370.400 187.500 371.600 ;
        RECT 186.800 369.600 187.600 370.400 ;
        RECT 182.000 367.600 182.800 368.400 ;
        RECT 177.200 343.600 178.000 344.400 ;
        RECT 177.300 340.400 177.900 343.600 ;
        RECT 177.200 339.600 178.000 340.400 ;
        RECT 175.600 337.600 176.400 338.400 ;
        RECT 182.100 336.400 182.700 367.600 ;
        RECT 191.600 364.200 192.400 377.800 ;
        RECT 193.200 364.200 194.000 377.800 ;
        RECT 194.800 366.200 195.600 377.800 ;
        RECT 196.400 377.600 197.200 378.400 ;
        RECT 196.500 374.400 197.100 377.600 ;
        RECT 196.400 373.600 197.200 374.400 ;
        RECT 198.000 366.200 198.800 377.800 ;
        RECT 199.600 375.600 200.400 376.400 ;
        RECT 199.700 362.400 200.300 375.600 ;
        RECT 201.200 366.200 202.000 377.800 ;
        RECT 202.800 364.200 203.600 377.800 ;
        RECT 204.400 364.200 205.200 377.800 ;
        RECT 206.000 364.200 206.800 377.800 ;
        RECT 218.800 377.600 219.600 378.400 ;
        RECT 249.200 375.600 250.000 376.400 ;
        RECT 228.400 373.600 229.200 374.400 ;
        RECT 234.800 373.600 235.600 374.400 ;
        RECT 236.400 373.600 237.200 374.400 ;
        RECT 239.600 373.600 240.400 374.400 ;
        RECT 242.800 373.600 243.600 374.400 ;
        RECT 246.000 373.600 246.800 374.400 ;
        RECT 247.600 373.600 248.400 374.400 ;
        RECT 228.500 372.400 229.100 373.600 ;
        RECT 234.900 372.400 235.500 373.600 ;
        RECT 226.800 371.600 227.600 372.400 ;
        RECT 228.400 371.600 229.200 372.400 ;
        RECT 233.200 371.600 234.000 372.400 ;
        RECT 234.800 371.600 235.600 372.400 ;
        RECT 226.900 370.400 227.500 371.600 ;
        RECT 233.300 370.400 233.900 371.600 ;
        RECT 215.600 369.600 216.400 370.400 ;
        RECT 218.800 369.600 219.600 370.400 ;
        RECT 222.000 369.600 222.800 370.400 ;
        RECT 226.800 369.600 227.600 370.400 ;
        RECT 233.200 369.600 234.000 370.400 ;
        RECT 236.400 369.600 237.200 370.400 ;
        RECT 239.700 370.300 240.300 373.600 ;
        RECT 246.100 372.400 246.700 373.600 ;
        RECT 244.400 371.600 245.200 372.400 ;
        RECT 246.000 371.600 246.800 372.400 ;
        RECT 244.500 370.400 245.100 371.600 ;
        RECT 239.700 369.700 241.900 370.300 ;
        RECT 193.200 361.600 194.000 362.400 ;
        RECT 199.600 361.600 200.400 362.400 ;
        RECT 186.800 344.200 187.600 357.800 ;
        RECT 188.400 344.200 189.200 357.800 ;
        RECT 190.000 344.200 190.800 357.800 ;
        RECT 191.600 344.200 192.400 355.800 ;
        RECT 193.300 346.400 193.900 361.600 ;
        RECT 193.200 345.600 194.000 346.400 ;
        RECT 193.300 342.400 193.900 345.600 ;
        RECT 194.800 344.200 195.600 355.800 ;
        RECT 196.400 347.600 197.200 348.400 ;
        RECT 196.500 342.400 197.100 347.600 ;
        RECT 198.000 344.200 198.800 355.800 ;
        RECT 199.600 344.200 200.400 357.800 ;
        RECT 201.200 344.200 202.000 357.800 ;
        RECT 215.700 352.400 216.300 369.600 ;
        RECT 218.900 364.400 219.500 369.600 ;
        RECT 236.500 368.400 237.100 369.600 ;
        RECT 230.000 367.600 230.800 368.400 ;
        RECT 233.200 367.600 234.000 368.400 ;
        RECT 236.400 367.600 237.200 368.400 ;
        RECT 239.600 367.600 240.400 368.400 ;
        RECT 239.700 366.400 240.300 367.600 ;
        RECT 241.300 366.400 241.900 369.700 ;
        RECT 244.400 369.600 245.200 370.400 ;
        RECT 250.800 369.600 251.600 370.400 ;
        RECT 250.900 368.400 251.500 369.600 ;
        RECT 250.800 367.600 251.600 368.400 ;
        RECT 239.600 365.600 240.400 366.400 ;
        RECT 241.200 365.600 242.000 366.400 ;
        RECT 252.400 365.600 253.200 366.400 ;
        RECT 255.600 365.600 256.400 366.400 ;
        RECT 218.800 363.600 219.600 364.400 ;
        RECT 246.000 363.600 246.800 364.400 ;
        RECT 246.100 358.400 246.700 363.600 ;
        RECT 252.500 358.400 253.100 365.600 ;
        RECT 254.000 363.600 254.800 364.400 ;
        RECT 254.100 358.400 254.700 363.600 ;
        RECT 215.600 351.600 216.400 352.400 ;
        RECT 206.000 349.600 206.800 350.400 ;
        RECT 209.200 349.600 210.000 350.400 ;
        RECT 220.400 349.600 221.200 350.400 ;
        RECT 193.200 341.600 194.000 342.400 ;
        RECT 196.400 341.600 197.200 342.400 ;
        RECT 199.600 341.600 200.400 342.400 ;
        RECT 191.600 339.600 192.400 340.400 ;
        RECT 191.700 336.400 192.300 339.600 ;
        RECT 199.700 338.400 200.300 341.600 ;
        RECT 209.300 338.400 209.900 349.600 ;
        RECT 212.400 344.300 213.200 344.400 ;
        RECT 212.400 343.700 214.700 344.300 ;
        RECT 212.400 343.600 213.200 343.700 ;
        RECT 194.800 337.600 195.600 338.400 ;
        RECT 199.600 337.600 200.400 338.400 ;
        RECT 209.200 337.600 210.000 338.400 ;
        RECT 182.000 335.600 182.800 336.400 ;
        RECT 191.600 335.600 192.400 336.400 ;
        RECT 180.400 331.600 181.200 332.400 ;
        RECT 175.600 329.600 176.400 330.400 ;
        RECT 172.400 317.600 173.200 318.400 ;
        RECT 175.600 313.600 176.400 314.400 ;
        RECT 172.400 311.600 173.200 312.400 ;
        RECT 175.700 310.400 176.300 313.600 ;
        RECT 177.200 311.600 178.000 312.400 ;
        RECT 167.600 309.600 168.400 310.400 ;
        RECT 169.200 309.600 170.000 310.400 ;
        RECT 170.800 309.600 171.600 310.400 ;
        RECT 175.600 309.600 176.400 310.400 ;
        RECT 170.800 307.600 171.600 308.400 ;
        RECT 169.200 301.600 170.000 302.400 ;
        RECT 162.800 297.600 163.600 298.400 ;
        RECT 166.000 297.600 166.800 298.400 ;
        RECT 169.300 296.400 169.900 301.600 ;
        RECT 169.200 295.600 170.000 296.400 ;
        RECT 164.400 293.600 165.200 294.400 ;
        RECT 167.600 292.300 168.400 292.400 ;
        RECT 159.600 291.700 161.900 292.300 ;
        RECT 166.100 291.700 168.400 292.300 ;
        RECT 159.600 291.600 160.400 291.700 ;
        RECT 102.000 283.600 102.800 284.400 ;
        RECT 98.800 264.200 99.600 277.800 ;
        RECT 100.400 264.200 101.200 277.800 ;
        RECT 102.000 264.200 102.800 275.800 ;
        RECT 103.700 270.400 104.300 291.600 ;
        RECT 122.900 290.400 123.500 291.600 ;
        RECT 108.400 289.600 109.200 290.400 ;
        RECT 113.200 290.300 114.000 290.400 ;
        RECT 113.200 289.700 115.500 290.300 ;
        RECT 113.200 289.600 114.000 289.700 ;
        RECT 108.500 284.400 109.100 289.600 ;
        RECT 108.400 283.600 109.200 284.400 ;
        RECT 103.600 269.600 104.400 270.400 ;
        RECT 103.600 267.600 104.400 268.400 ;
        RECT 103.700 264.400 104.300 267.600 ;
        RECT 103.600 263.600 104.400 264.400 ;
        RECT 105.200 264.200 106.000 275.800 ;
        RECT 106.800 265.600 107.600 266.400 ;
        RECT 106.900 260.400 107.500 265.600 ;
        RECT 108.400 264.200 109.200 275.800 ;
        RECT 110.000 264.200 110.800 277.800 ;
        RECT 111.600 264.200 112.400 277.800 ;
        RECT 113.200 264.200 114.000 277.800 ;
        RECT 114.900 272.400 115.500 289.700 ;
        RECT 122.800 289.600 123.600 290.400 ;
        RECT 132.400 289.600 133.200 290.400 ;
        RECT 135.600 289.600 136.400 290.400 ;
        RECT 145.200 289.600 146.000 290.400 ;
        RECT 151.600 289.600 152.400 290.400 ;
        RECT 162.800 289.600 163.600 290.400 ;
        RECT 129.200 287.600 130.000 288.400 ;
        RECT 114.800 271.600 115.600 272.400 ;
        RECT 132.500 270.400 133.100 289.600 ;
        RECT 135.700 284.400 136.300 289.600 ;
        RECT 134.000 283.600 134.800 284.400 ;
        RECT 135.600 283.600 136.400 284.400 ;
        RECT 134.100 278.400 134.700 283.600 ;
        RECT 134.000 277.600 134.800 278.400 ;
        RECT 145.300 276.400 145.900 289.600 ;
        RECT 148.400 287.600 149.200 288.400 ;
        RECT 150.000 283.600 150.800 284.400 ;
        RECT 145.200 275.600 146.000 276.400 ;
        RECT 150.100 274.400 150.700 283.600 ;
        RECT 150.000 273.600 150.800 274.400 ;
        RECT 140.400 271.600 141.200 272.400 ;
        RECT 145.200 271.600 146.000 272.400 ;
        RECT 114.800 269.600 115.600 270.400 ;
        RECT 132.400 269.600 133.200 270.400 ;
        RECT 138.800 269.600 139.600 270.400 ;
        RECT 90.800 259.600 91.600 260.400 ;
        RECT 97.200 259.600 98.000 260.400 ;
        RECT 106.800 259.600 107.600 260.400 ;
        RECT 90.800 244.200 91.600 257.800 ;
        RECT 92.400 244.200 93.200 257.800 ;
        RECT 94.000 244.200 94.800 257.800 ;
        RECT 95.600 246.200 96.400 257.800 ;
        RECT 97.300 256.400 97.900 259.600 ;
        RECT 97.200 255.600 98.000 256.400 ;
        RECT 98.800 246.200 99.600 257.800 ;
        RECT 100.400 253.600 101.200 254.400 ;
        RECT 100.500 252.400 101.100 253.600 ;
        RECT 100.400 251.600 101.200 252.400 ;
        RECT 102.000 246.200 102.800 257.800 ;
        RECT 103.600 244.200 104.400 257.800 ;
        RECT 105.200 244.200 106.000 257.800 ;
        RECT 110.000 251.600 110.800 252.400 ;
        RECT 110.100 248.400 110.700 251.600 ;
        RECT 114.900 248.400 115.500 269.600 ;
        RECT 122.800 267.600 123.600 268.400 ;
        RECT 132.400 267.600 133.200 268.400 ;
        RECT 134.000 267.600 134.800 268.400 ;
        RECT 138.800 267.600 139.600 268.400 ;
        RECT 119.600 259.600 120.400 260.400 ;
        RECT 110.000 247.600 110.800 248.400 ;
        RECT 114.800 247.600 115.600 248.400 ;
        RECT 103.600 239.600 104.400 240.400 ;
        RECT 102.000 237.600 102.800 238.400 ;
        RECT 100.400 235.600 101.200 236.400 ;
        RECT 89.200 229.600 90.000 230.400 ;
        RECT 92.400 229.600 93.200 230.400 ;
        RECT 92.500 214.400 93.100 229.600 ;
        RECT 100.500 228.400 101.100 235.600 ;
        RECT 102.100 230.400 102.700 237.600 ;
        RECT 102.000 229.600 102.800 230.400 ;
        RECT 100.400 227.600 101.200 228.400 ;
        RECT 102.000 227.600 102.800 228.400 ;
        RECT 97.200 225.600 98.000 226.400 ;
        RECT 97.300 224.400 97.900 225.600 ;
        RECT 95.600 223.600 96.400 224.400 ;
        RECT 97.200 223.600 98.000 224.400 ;
        RECT 98.800 223.600 99.600 224.400 ;
        RECT 95.700 220.300 96.300 223.600 ;
        RECT 94.100 219.700 96.300 220.300 ;
        RECT 94.100 214.400 94.700 219.700 ;
        RECT 95.600 217.600 96.400 218.400 ;
        RECT 97.200 216.300 98.000 216.400 ;
        RECT 95.700 215.700 98.000 216.300 ;
        RECT 89.200 213.600 90.000 214.400 ;
        RECT 92.400 213.600 93.200 214.400 ;
        RECT 94.000 213.600 94.800 214.400 ;
        RECT 87.600 211.600 88.400 212.400 ;
        RECT 92.400 211.600 93.200 212.400 ;
        RECT 87.700 210.400 88.300 211.600 ;
        RECT 87.600 209.600 88.400 210.400 ;
        RECT 66.800 191.600 67.600 192.400 ;
        RECT 65.200 189.600 66.000 190.400 ;
        RECT 65.300 188.400 65.900 189.600 ;
        RECT 65.200 187.600 66.000 188.400 ;
        RECT 74.800 184.200 75.600 197.800 ;
        RECT 76.400 184.200 77.200 197.800 ;
        RECT 82.800 197.600 83.600 198.400 ;
        RECT 78.000 184.200 78.800 195.800 ;
        RECT 79.600 187.600 80.400 188.400 ;
        RECT 81.200 184.200 82.000 195.800 ;
        RECT 82.800 185.600 83.600 186.400 ;
        RECT 82.900 178.400 83.500 185.600 ;
        RECT 84.400 184.200 85.200 195.800 ;
        RECT 86.000 184.200 86.800 197.800 ;
        RECT 87.600 184.200 88.400 197.800 ;
        RECT 89.200 184.200 90.000 197.800 ;
        RECT 95.700 196.400 96.300 215.700 ;
        RECT 97.200 215.600 98.000 215.700 ;
        RECT 97.200 213.600 98.000 214.400 ;
        RECT 98.900 200.400 99.500 223.600 ;
        RECT 102.100 210.400 102.700 227.600 ;
        RECT 103.700 214.400 104.300 239.600 ;
        RECT 119.700 238.300 120.300 259.600 ;
        RECT 122.900 258.400 123.500 267.600 ;
        RECT 122.800 257.600 123.600 258.400 ;
        RECT 132.500 256.400 133.100 267.600 ;
        RECT 134.100 266.400 134.700 267.600 ;
        RECT 134.000 265.600 134.800 266.400 ;
        RECT 132.400 255.600 133.200 256.400 ;
        RECT 122.800 253.600 123.600 254.400 ;
        RECT 121.200 251.600 122.000 252.400 ;
        RECT 122.900 250.400 123.500 253.600 ;
        RECT 132.500 252.400 133.100 255.600 ;
        RECT 134.100 254.300 134.700 265.600 ;
        RECT 137.200 261.600 138.000 262.400 ;
        RECT 137.300 258.400 137.900 261.600 ;
        RECT 137.200 257.600 138.000 258.400 ;
        RECT 138.900 254.400 139.500 267.600 ;
        RECT 140.500 262.400 141.100 271.600 ;
        RECT 142.000 269.600 142.800 270.400 ;
        RECT 142.000 263.600 142.800 264.400 ;
        RECT 140.400 261.600 141.200 262.400 ;
        RECT 142.100 258.400 142.700 263.600 ;
        RECT 142.000 257.600 142.800 258.400 ;
        RECT 143.600 255.600 144.400 256.400 ;
        RECT 135.600 254.300 136.400 254.400 ;
        RECT 134.100 253.700 136.400 254.300 ;
        RECT 135.600 253.600 136.400 253.700 ;
        RECT 138.800 253.600 139.600 254.400 ;
        RECT 132.400 251.600 133.200 252.400 ;
        RECT 122.800 249.600 123.600 250.400 ;
        RECT 134.000 247.600 134.800 248.400 ;
        RECT 105.000 229.600 106.000 230.400 ;
        RECT 113.200 223.600 114.000 224.400 ;
        RECT 114.800 224.200 115.600 237.800 ;
        RECT 116.400 224.200 117.200 237.800 ;
        RECT 118.000 224.200 118.800 237.800 ;
        RECT 119.700 237.700 121.900 238.300 ;
        RECT 119.600 224.200 120.400 235.800 ;
        RECT 121.300 226.400 121.900 237.700 ;
        RECT 121.200 225.600 122.000 226.400 ;
        RECT 122.800 224.200 123.600 235.800 ;
        RECT 124.400 227.600 125.200 228.400 ;
        RECT 124.500 224.400 125.100 227.600 ;
        RECT 124.400 223.600 125.200 224.400 ;
        RECT 126.000 224.200 126.800 235.800 ;
        RECT 127.600 224.200 128.400 237.800 ;
        RECT 129.200 224.200 130.000 237.800 ;
        RECT 134.100 230.400 134.700 247.600 ;
        RECT 135.700 246.400 136.300 253.600 ;
        RECT 135.600 245.600 136.400 246.400 ;
        RECT 134.000 229.600 134.800 230.400 ;
        RECT 138.900 228.400 139.500 253.600 ;
        RECT 140.400 252.300 141.200 252.400 ;
        RECT 140.400 251.700 142.700 252.300 ;
        RECT 140.400 251.600 141.200 251.700 ;
        RECT 140.400 247.600 141.200 248.400 ;
        RECT 138.800 227.600 139.600 228.400 ;
        RECT 113.300 218.400 113.900 223.600 ;
        RECT 113.200 217.600 114.000 218.400 ;
        RECT 103.600 213.600 104.400 214.400 ;
        RECT 105.200 211.600 106.000 212.400 ;
        RECT 100.400 209.600 101.200 210.400 ;
        RECT 102.000 209.600 102.800 210.400 ;
        RECT 98.800 199.600 99.600 200.400 ;
        RECT 98.800 197.600 99.600 198.400 ;
        RECT 95.600 195.600 96.400 196.400 ;
        RECT 98.800 195.600 99.600 196.400 ;
        RECT 90.800 191.600 91.600 192.400 ;
        RECT 90.900 190.400 91.500 191.600 ;
        RECT 90.800 189.600 91.600 190.400 ;
        RECT 66.800 164.200 67.600 177.800 ;
        RECT 68.400 164.200 69.200 177.800 ;
        RECT 70.000 164.200 70.800 177.800 ;
        RECT 71.600 166.200 72.400 177.800 ;
        RECT 73.200 177.600 74.000 178.400 ;
        RECT 73.300 176.400 73.900 177.600 ;
        RECT 73.200 175.600 74.000 176.400 ;
        RECT 63.600 155.600 64.400 156.400 ;
        RECT 65.200 151.600 66.000 152.400 ;
        RECT 57.200 147.600 58.000 148.400 ;
        RECT 58.800 147.600 59.600 148.400 ;
        RECT 62.000 147.600 62.800 148.400 ;
        RECT 65.200 147.600 66.000 148.400 ;
        RECT 57.300 120.400 57.900 147.600 ;
        RECT 58.900 130.400 59.500 147.600 ;
        RECT 73.300 146.400 73.900 175.600 ;
        RECT 74.800 166.200 75.600 177.800 ;
        RECT 76.400 175.600 77.200 176.400 ;
        RECT 76.500 174.400 77.100 175.600 ;
        RECT 76.400 173.600 77.200 174.400 ;
        RECT 78.000 166.200 78.800 177.800 ;
        RECT 79.600 164.200 80.400 177.800 ;
        RECT 81.200 164.200 82.000 177.800 ;
        RECT 82.800 177.600 83.600 178.400 ;
        RECT 90.900 176.400 91.500 189.600 ;
        RECT 92.400 185.600 93.200 186.400 ;
        RECT 86.000 175.600 86.800 176.400 ;
        RECT 90.800 175.600 91.600 176.400 ;
        RECT 86.100 172.400 86.700 175.600 ;
        RECT 90.800 173.600 91.600 174.400 ;
        RECT 86.000 171.600 86.800 172.400 ;
        RECT 90.900 162.400 91.500 173.600 ;
        RECT 92.500 172.400 93.100 185.600 ;
        RECT 98.900 176.300 99.500 195.600 ;
        RECT 100.400 176.300 101.200 176.400 ;
        RECT 98.900 175.700 101.200 176.300 ;
        RECT 92.400 171.600 93.200 172.400 ;
        RECT 97.200 171.600 98.000 172.400 ;
        RECT 95.600 169.600 96.400 170.400 ;
        RECT 95.700 168.400 96.300 169.600 ;
        RECT 95.600 167.600 96.400 168.400 ;
        RECT 90.800 161.600 91.600 162.400 ;
        RECT 79.600 149.600 80.400 150.400 ;
        RECT 66.800 145.600 67.600 146.400 ;
        RECT 73.200 145.600 74.000 146.400 ;
        RECT 58.800 129.600 59.600 130.400 ;
        RECT 60.400 124.200 61.200 137.800 ;
        RECT 62.000 124.200 62.800 137.800 ;
        RECT 63.600 124.200 64.400 137.800 ;
        RECT 65.200 126.200 66.000 137.800 ;
        RECT 66.900 136.400 67.500 145.600 ;
        RECT 71.600 143.600 72.400 144.400 ;
        RECT 71.700 142.400 72.300 143.600 ;
        RECT 71.600 141.600 72.400 142.400 ;
        RECT 66.800 135.600 67.600 136.400 ;
        RECT 66.900 120.400 67.500 135.600 ;
        RECT 68.400 126.200 69.200 137.800 ;
        RECT 70.000 133.600 70.800 134.400 ;
        RECT 70.000 131.600 70.800 132.400 ;
        RECT 57.200 119.600 58.000 120.400 ;
        RECT 60.400 119.600 61.200 120.400 ;
        RECT 66.800 119.600 67.600 120.400 ;
        RECT 52.400 107.600 53.200 108.400 ;
        RECT 54.000 104.200 54.800 117.800 ;
        RECT 55.600 104.200 56.400 117.800 ;
        RECT 57.200 104.200 58.000 117.800 ;
        RECT 58.800 104.200 59.600 115.800 ;
        RECT 60.500 106.400 61.100 119.600 ;
        RECT 60.400 105.600 61.200 106.400 ;
        RECT 60.500 102.300 61.100 105.600 ;
        RECT 62.000 104.200 62.800 115.800 ;
        RECT 63.600 107.600 64.400 108.400 ;
        RECT 63.700 106.400 64.300 107.600 ;
        RECT 63.600 105.600 64.400 106.400 ;
        RECT 65.200 104.200 66.000 115.800 ;
        RECT 66.800 104.200 67.600 117.800 ;
        RECT 68.400 104.200 69.200 117.800 ;
        RECT 70.100 110.400 70.700 131.600 ;
        RECT 71.600 126.200 72.400 137.800 ;
        RECT 73.200 124.200 74.000 137.800 ;
        RECT 74.800 124.200 75.600 137.800 ;
        RECT 78.000 135.600 78.800 136.400 ;
        RECT 70.000 109.600 70.800 110.400 ;
        RECT 78.100 108.400 78.700 135.600 ;
        RECT 79.700 132.400 80.300 149.600 ;
        RECT 81.200 144.200 82.000 157.800 ;
        RECT 82.800 144.200 83.600 157.800 ;
        RECT 84.400 144.200 85.200 157.800 ;
        RECT 86.000 144.200 86.800 155.800 ;
        RECT 87.600 145.600 88.400 146.400 ;
        RECT 89.200 144.200 90.000 155.800 ;
        RECT 90.800 147.600 91.600 148.400 ;
        RECT 92.400 144.200 93.200 155.800 ;
        RECT 94.000 144.200 94.800 157.800 ;
        RECT 95.600 144.200 96.400 157.800 ;
        RECT 97.200 143.600 98.000 144.400 ;
        RECT 89.200 141.600 90.000 142.400 ;
        RECT 89.300 138.400 89.900 141.600 ;
        RECT 89.200 137.600 90.000 138.400 ;
        RECT 97.300 136.400 97.900 143.600 ;
        RECT 98.900 142.400 99.500 175.700 ;
        RECT 100.400 175.600 101.200 175.700 ;
        RECT 100.400 173.600 101.200 174.400 ;
        RECT 100.500 172.400 101.100 173.600 ;
        RECT 100.400 171.600 101.200 172.400 ;
        RECT 102.100 152.400 102.700 209.600 ;
        RECT 105.300 208.400 105.900 211.600 ;
        RECT 108.400 209.600 109.200 210.400 ;
        RECT 105.200 207.600 106.000 208.400 ;
        RECT 124.400 204.200 125.200 217.800 ;
        RECT 126.000 204.200 126.800 217.800 ;
        RECT 127.600 206.200 128.400 217.800 ;
        RECT 129.200 213.600 130.000 214.400 ;
        RECT 129.200 211.600 130.000 212.400 ;
        RECT 103.600 183.600 104.400 184.400 ;
        RECT 113.200 184.200 114.000 197.800 ;
        RECT 114.800 184.200 115.600 197.800 ;
        RECT 116.400 184.200 117.200 197.800 ;
        RECT 118.000 184.200 118.800 195.800 ;
        RECT 119.600 185.600 120.400 186.400 ;
        RECT 103.700 156.400 104.300 183.600 ;
        RECT 119.700 178.400 120.300 185.600 ;
        RECT 121.200 184.200 122.000 195.800 ;
        RECT 122.800 187.600 123.600 188.400 ;
        RECT 124.400 184.200 125.200 195.800 ;
        RECT 126.000 184.200 126.800 197.800 ;
        RECT 127.600 184.200 128.400 197.800 ;
        RECT 129.300 192.400 129.900 211.600 ;
        RECT 130.800 206.200 131.600 217.800 ;
        RECT 132.400 215.600 133.200 216.400 ;
        RECT 132.500 204.300 133.100 215.600 ;
        RECT 134.000 206.200 134.800 217.800 ;
        RECT 132.500 203.700 134.700 204.300 ;
        RECT 135.600 204.200 136.400 217.800 ;
        RECT 137.200 204.200 138.000 217.800 ;
        RECT 138.800 204.200 139.600 217.800 ;
        RECT 140.500 212.400 141.100 247.600 ;
        RECT 140.400 211.600 141.200 212.400 ;
        RECT 129.200 191.200 130.000 192.400 ;
        RECT 134.100 178.400 134.700 203.700 ;
        RECT 142.100 196.400 142.700 251.700 ;
        RECT 145.300 232.400 145.900 271.600 ;
        RECT 148.400 269.600 149.200 270.400 ;
        RECT 148.500 268.400 149.100 269.600 ;
        RECT 151.700 268.400 152.300 289.600 ;
        RECT 162.900 284.400 163.500 289.600 ;
        RECT 162.800 283.600 163.600 284.400 ;
        RECT 161.200 273.600 162.000 274.400 ;
        RECT 161.300 270.400 161.900 273.600 ;
        RECT 156.400 269.600 157.200 270.400 ;
        RECT 161.200 269.600 162.000 270.400 ;
        RECT 162.900 268.400 163.500 283.600 ;
        RECT 166.100 272.400 166.700 291.700 ;
        RECT 167.600 291.600 168.400 291.700 ;
        RECT 167.600 289.600 168.400 290.400 ;
        RECT 167.700 282.400 168.300 289.600 ;
        RECT 169.200 287.600 170.000 288.400 ;
        RECT 167.600 281.600 168.400 282.400 ;
        RECT 167.600 273.600 168.400 274.400 ;
        RECT 166.000 271.600 166.800 272.400 ;
        RECT 166.100 270.400 166.700 271.600 ;
        RECT 166.000 269.600 166.800 270.400 ;
        RECT 148.400 267.600 149.200 268.400 ;
        RECT 151.600 267.600 152.400 268.400 ;
        RECT 154.800 267.600 155.600 268.400 ;
        RECT 162.800 267.600 163.600 268.400 ;
        RECT 167.600 267.600 168.400 268.400 ;
        RECT 151.600 265.600 152.400 266.400 ;
        RECT 158.000 265.600 158.800 266.400 ;
        RECT 151.700 264.400 152.300 265.600 ;
        RECT 151.600 263.600 152.400 264.400 ;
        RECT 150.000 249.600 150.800 250.400 ;
        RECT 146.800 245.600 147.600 246.400 ;
        RECT 146.900 238.400 147.500 245.600 ;
        RECT 146.800 237.600 147.600 238.400 ;
        RECT 150.100 234.400 150.700 249.600 ;
        RECT 153.200 244.200 154.000 257.800 ;
        RECT 154.800 244.200 155.600 257.800 ;
        RECT 156.400 246.200 157.200 257.800 ;
        RECT 158.100 256.400 158.700 265.600 ;
        RECT 166.000 263.600 166.800 264.400 ;
        RECT 166.100 260.400 166.700 263.600 ;
        RECT 167.700 262.400 168.300 267.600 ;
        RECT 167.600 261.600 168.400 262.400 ;
        RECT 166.000 259.600 166.800 260.400 ;
        RECT 158.000 255.600 158.800 256.400 ;
        RECT 158.000 253.600 158.800 254.400 ;
        RECT 158.000 251.600 158.800 252.400 ;
        RECT 158.100 248.400 158.700 251.600 ;
        RECT 158.000 247.600 158.800 248.400 ;
        RECT 159.600 246.200 160.400 257.800 ;
        RECT 161.200 255.600 162.000 256.400 ;
        RECT 161.300 254.400 161.900 255.600 ;
        RECT 161.200 253.600 162.000 254.400 ;
        RECT 162.800 246.200 163.600 257.800 ;
        RECT 164.400 244.200 165.200 257.800 ;
        RECT 166.000 244.200 166.800 257.800 ;
        RECT 167.600 244.200 168.400 257.800 ;
        RECT 169.300 252.400 169.900 287.600 ;
        RECT 170.900 280.400 171.500 307.600 ;
        RECT 175.700 306.400 176.300 309.600 ;
        RECT 175.600 305.600 176.400 306.400 ;
        RECT 177.300 298.400 177.900 311.600 ;
        RECT 180.500 310.400 181.100 331.600 ;
        RECT 182.100 322.400 182.700 335.600 ;
        RECT 186.800 333.600 187.600 334.400 ;
        RECT 186.900 332.400 187.500 333.600 ;
        RECT 186.800 331.600 187.600 332.400 ;
        RECT 188.400 329.600 189.200 330.400 ;
        RECT 188.500 328.400 189.100 329.600 ;
        RECT 188.400 327.600 189.200 328.400 ;
        RECT 186.800 323.600 187.600 324.400 ;
        RECT 182.000 321.600 182.800 322.400 ;
        RECT 182.000 317.600 182.800 318.400 ;
        RECT 182.100 312.400 182.700 317.600 ;
        RECT 182.000 311.600 182.800 312.400 ;
        RECT 180.400 309.600 181.200 310.400 ;
        RECT 180.500 306.400 181.100 309.600 ;
        RECT 186.900 306.400 187.500 323.600 ;
        RECT 191.700 318.400 192.300 335.600 ;
        RECT 193.200 333.600 194.000 334.400 ;
        RECT 194.900 318.400 195.500 337.600 ;
        RECT 214.100 336.400 214.700 343.700 ;
        RECT 214.000 335.600 214.800 336.400 ;
        RECT 201.200 333.600 202.000 334.400 ;
        RECT 212.400 333.600 213.200 334.400 ;
        RECT 196.400 331.600 197.200 332.400 ;
        RECT 191.600 317.600 192.400 318.400 ;
        RECT 194.800 317.600 195.600 318.400 ;
        RECT 191.600 311.600 192.400 312.400 ;
        RECT 190.000 309.600 190.800 310.400 ;
        RECT 178.800 305.600 179.600 306.400 ;
        RECT 180.400 305.600 181.200 306.400 ;
        RECT 186.800 305.600 187.600 306.400 ;
        RECT 178.900 302.400 179.500 305.600 ;
        RECT 183.600 303.600 184.400 304.400 ;
        RECT 178.800 301.600 179.600 302.400 ;
        RECT 177.200 297.600 178.000 298.400 ;
        RECT 175.600 293.600 176.400 294.400 ;
        RECT 180.400 293.600 181.200 294.400 ;
        RECT 172.400 291.600 173.200 292.400 ;
        RECT 174.000 291.600 174.800 292.400 ;
        RECT 172.500 284.400 173.100 291.600 ;
        RECT 174.100 290.400 174.700 291.600 ;
        RECT 174.000 289.600 174.800 290.400 ;
        RECT 172.400 283.600 173.200 284.400 ;
        RECT 170.800 279.600 171.600 280.400 ;
        RECT 174.000 277.600 174.800 278.400 ;
        RECT 175.700 276.300 176.300 293.600 ;
        RECT 178.800 281.600 179.600 282.400 ;
        RECT 174.100 275.700 176.300 276.300 ;
        RECT 174.100 274.400 174.700 275.700 ;
        RECT 172.400 273.600 173.200 274.400 ;
        RECT 174.000 273.600 174.800 274.400 ;
        RECT 175.600 273.600 176.400 274.400 ;
        RECT 172.500 272.400 173.100 273.600 ;
        RECT 178.900 272.400 179.500 281.600 ;
        RECT 180.500 272.400 181.100 293.600 ;
        RECT 182.000 290.300 182.800 290.400 ;
        RECT 183.700 290.300 184.300 303.600 ;
        RECT 185.200 301.600 186.000 302.400 ;
        RECT 185.300 290.400 185.900 301.600 ;
        RECT 186.900 294.400 187.500 305.600 ;
        RECT 186.800 293.600 187.600 294.400 ;
        RECT 190.100 292.400 190.700 309.600 ;
        RECT 191.700 306.400 192.300 311.600 ;
        RECT 194.800 310.300 195.600 310.400 ;
        RECT 196.500 310.300 197.100 331.600 ;
        RECT 212.500 330.400 213.100 333.600 ;
        RECT 199.600 329.600 200.400 330.400 ;
        RECT 204.400 329.600 205.200 330.400 ;
        RECT 212.400 329.600 213.200 330.400 ;
        RECT 199.700 316.400 200.300 329.600 ;
        RECT 202.800 323.600 203.600 324.400 ;
        RECT 210.800 323.600 211.600 324.400 ;
        RECT 199.600 315.600 200.400 316.400 ;
        RECT 201.200 311.600 202.000 312.400 ;
        RECT 194.800 309.700 197.100 310.300 ;
        RECT 194.800 309.600 195.600 309.700 ;
        RECT 196.400 307.600 197.200 308.400 ;
        RECT 199.600 308.300 200.400 308.400 ;
        RECT 198.100 307.700 200.400 308.300 ;
        RECT 191.600 305.600 192.400 306.400 ;
        RECT 196.500 296.300 197.100 307.600 ;
        RECT 198.100 296.400 198.700 307.700 ;
        RECT 199.600 307.600 200.400 307.700 ;
        RECT 199.600 306.300 200.400 306.400 ;
        RECT 201.300 306.300 201.900 311.600 ;
        RECT 202.900 310.400 203.500 323.600 ;
        RECT 206.000 321.600 206.800 322.400 ;
        RECT 210.900 322.300 211.500 323.600 ;
        RECT 209.300 321.700 211.500 322.300 ;
        RECT 206.100 312.400 206.700 321.600 ;
        RECT 209.300 314.400 209.900 321.700 ;
        RECT 212.400 321.600 213.200 322.400 ;
        RECT 210.800 317.600 211.600 318.400 ;
        RECT 209.200 313.600 210.000 314.400 ;
        RECT 206.000 311.600 206.800 312.400 ;
        RECT 209.300 310.400 209.900 313.600 ;
        RECT 202.800 309.600 203.600 310.400 ;
        RECT 209.200 309.600 210.000 310.400 ;
        RECT 210.900 308.400 211.500 317.600 ;
        RECT 212.500 308.400 213.100 321.600 ;
        RECT 214.100 318.400 214.700 335.600 ;
        RECT 220.500 332.400 221.100 349.600 ;
        RECT 222.000 344.200 222.800 357.800 ;
        RECT 223.600 344.200 224.400 357.800 ;
        RECT 225.200 344.200 226.000 357.800 ;
        RECT 226.800 344.200 227.600 355.800 ;
        RECT 228.400 345.600 229.200 346.400 ;
        RECT 228.500 336.400 229.100 345.600 ;
        RECT 230.000 344.200 230.800 355.800 ;
        RECT 231.600 347.600 232.400 348.400 ;
        RECT 231.700 344.400 232.300 347.600 ;
        RECT 231.600 343.600 232.400 344.400 ;
        RECT 233.200 344.200 234.000 355.800 ;
        RECT 234.800 344.200 235.600 357.800 ;
        RECT 236.400 344.200 237.200 357.800 ;
        RECT 246.000 357.600 246.800 358.400 ;
        RECT 252.400 357.600 253.200 358.400 ;
        RECT 254.000 357.600 254.800 358.400 ;
        RECT 249.200 355.600 250.000 356.400 ;
        RECT 254.000 355.600 254.800 356.400 ;
        RECT 247.600 353.600 248.400 354.400 ;
        RECT 242.800 349.600 243.600 350.400 ;
        RECT 228.400 335.600 229.200 336.400 ;
        RECT 220.400 331.600 221.200 332.400 ;
        RECT 228.400 331.600 229.200 332.400 ;
        RECT 220.400 323.600 221.200 324.400 ;
        RECT 230.000 324.200 230.800 337.800 ;
        RECT 231.600 324.200 232.400 337.800 ;
        RECT 233.200 324.200 234.000 337.800 ;
        RECT 234.800 326.200 235.600 337.800 ;
        RECT 236.400 335.600 237.200 336.400 ;
        RECT 214.000 317.600 214.800 318.400 ;
        RECT 218.800 313.600 219.600 314.400 ;
        RECT 218.900 312.400 219.500 313.600 ;
        RECT 215.600 311.600 216.400 312.400 ;
        RECT 217.200 311.600 218.000 312.400 ;
        RECT 218.800 311.600 219.600 312.400 ;
        RECT 220.500 312.300 221.100 323.600 ;
        RECT 233.200 319.600 234.000 320.400 ;
        RECT 226.800 317.600 227.600 318.400 ;
        RECT 222.000 312.300 222.800 312.400 ;
        RECT 220.500 311.700 222.800 312.300 ;
        RECT 222.000 311.600 222.800 311.700 ;
        RECT 214.000 309.600 214.800 310.400 ;
        RECT 210.800 307.600 211.600 308.400 ;
        RECT 212.400 307.600 213.200 308.400 ;
        RECT 199.600 305.700 201.900 306.300 ;
        RECT 199.600 305.600 200.400 305.700 ;
        RECT 202.800 303.600 203.600 304.400 ;
        RECT 202.900 302.400 203.500 303.600 ;
        RECT 199.600 301.600 200.400 302.400 ;
        RECT 202.800 301.600 203.600 302.400 ;
        RECT 194.900 295.700 197.100 296.300 ;
        RECT 191.600 293.600 192.400 294.400 ;
        RECT 190.000 292.300 190.800 292.400 ;
        RECT 191.600 292.300 192.400 292.400 ;
        RECT 190.000 291.700 192.400 292.300 ;
        RECT 190.000 291.600 190.800 291.700 ;
        RECT 191.600 291.600 192.400 291.700 ;
        RECT 182.000 289.700 184.300 290.300 ;
        RECT 182.000 289.600 182.800 289.700 ;
        RECT 185.200 289.600 186.000 290.400 ;
        RECT 182.100 288.400 182.700 289.600 ;
        RECT 182.000 287.600 182.800 288.400 ;
        RECT 193.200 283.600 194.000 284.400 ;
        RECT 185.200 279.600 186.000 280.400 ;
        RECT 170.800 271.600 171.600 272.400 ;
        RECT 172.400 271.600 173.200 272.400 ;
        RECT 178.800 271.600 179.600 272.400 ;
        RECT 180.400 271.600 181.200 272.400 ;
        RECT 183.600 271.600 184.400 272.400 ;
        RECT 169.200 251.600 170.000 252.400 ;
        RECT 151.600 241.600 152.400 242.400 ;
        RECT 150.000 233.600 150.800 234.400 ;
        RECT 145.200 231.600 146.000 232.400 ;
        RECT 145.200 227.600 146.000 228.400 ;
        RECT 145.300 226.400 145.900 227.600 ;
        RECT 151.700 226.400 152.300 241.600 ;
        RECT 161.200 233.600 162.000 234.400 ;
        RECT 153.200 231.600 154.000 232.400 ;
        RECT 156.400 231.600 157.200 232.400 ;
        RECT 158.000 231.600 158.800 232.400 ;
        RECT 145.200 225.600 146.000 226.400 ;
        RECT 151.600 225.600 152.400 226.400 ;
        RECT 146.800 223.600 147.600 224.400 ;
        RECT 146.900 220.400 147.500 223.600 ;
        RECT 146.800 219.600 147.600 220.400 ;
        RECT 151.700 216.400 152.300 225.600 ;
        RECT 151.600 215.600 152.400 216.400 ;
        RECT 154.800 215.600 155.600 216.400 ;
        RECT 154.900 212.400 155.500 215.600 ;
        RECT 156.500 214.400 157.100 231.600 ;
        RECT 158.100 230.400 158.700 231.600 ;
        RECT 161.300 230.400 161.900 233.600 ;
        RECT 162.800 231.600 163.600 232.400 ;
        RECT 164.400 231.600 165.200 232.400 ;
        RECT 166.000 231.600 166.800 232.400 ;
        RECT 162.900 230.400 163.500 231.600 ;
        RECT 158.000 229.600 158.800 230.400 ;
        RECT 159.600 229.600 160.400 230.400 ;
        RECT 161.200 229.600 162.000 230.400 ;
        RECT 162.800 229.600 163.600 230.400 ;
        RECT 159.700 228.400 160.300 229.600 ;
        RECT 158.000 227.600 158.800 228.400 ;
        RECT 159.600 227.600 160.400 228.400 ;
        RECT 159.700 222.400 160.300 227.600 ;
        RECT 159.600 221.600 160.400 222.400 ;
        RECT 162.800 221.600 163.600 222.400 ;
        RECT 156.400 213.600 157.200 214.400 ;
        RECT 158.000 213.600 158.800 214.400 ;
        RECT 159.600 213.600 160.400 214.400 ;
        RECT 161.200 213.600 162.000 214.400 ;
        RECT 151.600 211.600 152.400 212.400 ;
        RECT 154.800 211.600 155.600 212.400 ;
        RECT 151.700 210.400 152.300 211.600 ;
        RECT 159.700 210.400 160.300 213.600 ;
        RECT 161.300 212.400 161.900 213.600 ;
        RECT 162.900 212.400 163.500 221.600 ;
        RECT 164.500 214.400 165.100 231.600 ;
        RECT 169.300 230.400 169.900 251.600 ;
        RECT 170.900 234.400 171.500 271.600 ;
        RECT 174.000 269.600 174.800 270.400 ;
        RECT 177.200 269.600 178.000 270.400 ;
        RECT 174.100 264.400 174.700 269.600 ;
        RECT 175.600 267.600 176.400 268.400 ;
        RECT 174.000 263.600 174.800 264.400 ;
        RECT 175.700 238.400 176.300 267.600 ;
        RECT 177.300 258.400 177.900 269.600 ;
        RECT 178.900 266.400 179.500 271.600 ;
        RECT 178.800 265.600 179.600 266.400 ;
        RECT 180.500 266.300 181.100 271.600 ;
        RECT 182.000 269.600 182.800 270.400 ;
        RECT 182.100 268.400 182.700 269.600 ;
        RECT 182.000 267.600 182.800 268.400 ;
        RECT 183.700 266.300 184.300 271.600 ;
        RECT 180.500 265.700 184.300 266.300 ;
        RECT 178.800 263.600 179.600 264.400 ;
        RECT 182.100 258.400 182.700 265.700 ;
        RECT 177.200 257.600 178.000 258.400 ;
        RECT 182.000 257.600 182.800 258.400 ;
        RECT 182.000 247.600 182.800 248.400 ;
        RECT 182.100 238.400 182.700 247.600 ;
        RECT 175.600 237.600 176.400 238.400 ;
        RECT 182.000 237.600 182.800 238.400 ;
        RECT 170.800 233.600 171.600 234.400 ;
        RECT 177.200 233.600 178.000 234.400 ;
        RECT 180.400 233.600 181.200 234.400 ;
        RECT 180.500 232.400 181.100 233.600 ;
        RECT 170.800 231.600 171.600 232.400 ;
        RECT 178.800 231.600 179.600 232.400 ;
        RECT 180.400 231.600 181.200 232.400 ;
        RECT 169.200 229.600 170.000 230.400 ;
        RECT 170.900 228.400 171.500 231.600 ;
        RECT 166.000 227.600 166.800 228.400 ;
        RECT 169.200 227.600 170.000 228.400 ;
        RECT 170.800 227.600 171.600 228.400 ;
        RECT 172.400 228.000 173.200 228.800 ;
        RECT 169.300 224.400 169.900 227.600 ;
        RECT 172.500 224.400 173.100 228.000 ;
        RECT 174.000 227.600 174.800 228.400 ;
        RECT 177.200 227.600 178.000 228.400 ;
        RECT 169.200 223.600 170.000 224.400 ;
        RECT 172.400 223.600 173.200 224.400 ;
        RECT 167.600 219.600 168.400 220.400 ;
        RECT 167.700 214.400 168.300 219.600 ;
        RECT 169.200 215.600 170.000 216.400 ;
        RECT 169.300 214.400 169.900 215.600 ;
        RECT 174.100 214.400 174.700 227.600 ;
        RECT 175.600 223.600 176.400 224.400 ;
        RECT 175.700 218.400 176.300 223.600 ;
        RECT 175.600 217.600 176.400 218.400 ;
        RECT 177.300 216.400 177.900 227.600 ;
        RECT 178.900 226.400 179.500 231.600 ;
        RECT 178.800 225.600 179.600 226.400 ;
        RECT 178.800 221.600 179.600 222.400 ;
        RECT 177.200 215.600 178.000 216.400 ;
        RECT 164.400 213.600 165.200 214.400 ;
        RECT 167.600 213.600 168.400 214.400 ;
        RECT 169.200 213.600 170.000 214.400 ;
        RECT 174.000 213.600 174.800 214.400 ;
        RECT 161.200 211.600 162.000 212.400 ;
        RECT 162.800 211.600 163.600 212.400 ;
        RECT 174.000 211.600 174.800 212.400 ;
        RECT 151.600 209.600 152.400 210.400 ;
        RECT 159.600 209.600 160.400 210.400 ;
        RECT 166.000 209.600 166.800 210.400 ;
        RECT 150.000 199.600 150.800 200.400 ;
        RECT 142.000 195.600 142.800 196.400 ;
        RECT 148.400 191.600 149.200 192.400 ;
        RECT 148.500 190.400 149.100 191.600 ;
        RECT 148.400 189.600 149.200 190.400 ;
        RECT 119.600 177.600 120.400 178.400 ;
        RECT 105.200 173.600 106.000 174.400 ;
        RECT 106.800 173.600 107.600 174.400 ;
        RECT 106.900 172.400 107.500 173.600 ;
        RECT 106.800 171.600 107.600 172.400 ;
        RECT 110.000 171.600 110.800 172.400 ;
        RECT 110.100 156.400 110.700 171.600 ;
        RECT 118.000 164.300 118.800 164.400 ;
        RECT 118.000 163.700 120.300 164.300 ;
        RECT 127.600 164.200 128.400 177.800 ;
        RECT 129.200 164.200 130.000 177.800 ;
        RECT 130.800 164.200 131.600 177.800 ;
        RECT 132.400 166.200 133.200 177.800 ;
        RECT 134.000 177.600 134.800 178.400 ;
        RECT 134.100 176.400 134.700 177.600 ;
        RECT 134.000 175.600 134.800 176.400 ;
        RECT 118.000 163.600 118.800 163.700 ;
        RECT 119.700 158.400 120.300 163.700 ;
        RECT 119.600 157.600 120.400 158.400 ;
        RECT 103.600 155.600 104.400 156.400 ;
        RECT 108.400 155.600 109.200 156.400 ;
        RECT 110.000 155.600 110.800 156.400 ;
        RECT 102.000 151.600 102.800 152.400 ;
        RECT 106.800 151.600 107.600 152.400 ;
        RECT 100.400 149.600 101.200 150.400 ;
        RECT 105.200 149.600 106.000 150.400 ;
        RECT 98.800 141.600 99.600 142.400 ;
        RECT 84.400 135.600 85.200 136.400 ;
        RECT 92.400 135.600 93.200 136.400 ;
        RECT 97.200 135.600 98.000 136.400 ;
        RECT 90.800 133.600 91.600 134.400 ;
        RECT 79.600 131.600 80.400 132.400 ;
        RECT 86.000 129.600 86.800 130.400 ;
        RECT 86.000 121.600 86.800 122.400 ;
        RECT 82.800 111.600 83.600 112.400 ;
        RECT 79.600 109.600 80.400 110.400 ;
        RECT 79.700 108.400 80.300 109.600 ;
        RECT 78.000 107.600 78.800 108.400 ;
        RECT 79.600 107.600 80.400 108.400 ;
        RECT 84.400 107.600 85.200 108.400 ;
        RECT 81.200 103.600 82.000 104.400 ;
        RECT 82.800 103.600 83.600 104.400 ;
        RECT 60.500 101.700 62.700 102.300 ;
        RECT 44.400 97.600 45.200 98.400 ;
        RECT 46.000 97.600 46.800 98.400 ;
        RECT 49.200 97.600 50.000 98.400 ;
        RECT 39.600 93.600 40.400 94.400 ;
        RECT 42.800 93.600 43.600 94.400 ;
        RECT 39.700 92.400 40.300 93.600 ;
        RECT 39.600 91.600 40.400 92.400 ;
        RECT 41.200 91.600 42.000 92.400 ;
        RECT 41.300 90.400 41.900 91.600 ;
        RECT 44.500 90.400 45.100 97.600 ;
        RECT 46.000 95.600 46.800 96.400 ;
        RECT 38.000 89.600 38.800 90.400 ;
        RECT 41.200 89.600 42.000 90.400 ;
        RECT 44.400 89.600 45.200 90.400 ;
        RECT 38.100 88.400 38.700 89.600 ;
        RECT 38.000 87.600 38.800 88.400 ;
        RECT 36.400 71.600 37.200 72.400 ;
        RECT 39.600 71.600 40.400 72.400 ;
        RECT 46.100 70.400 46.700 95.600 ;
        RECT 47.600 89.600 48.400 90.400 ;
        RECT 22.000 69.600 22.800 70.400 ;
        RECT 26.800 69.600 27.600 70.400 ;
        RECT 28.400 69.600 29.200 70.400 ;
        RECT 31.600 69.600 32.400 70.400 ;
        RECT 46.000 69.600 46.800 70.400 ;
        RECT 25.200 65.600 26.000 66.400 ;
        RECT 25.300 64.400 25.900 65.600 ;
        RECT 25.200 63.600 26.000 64.400 ;
        RECT 22.000 57.600 22.800 58.400 ;
        RECT 1.200 55.600 2.000 56.400 ;
        RECT 4.400 55.600 5.200 56.400 ;
        RECT 9.200 55.600 10.000 56.400 ;
        RECT 12.400 55.600 13.200 56.400 ;
        RECT 20.400 55.600 21.200 56.400 ;
        RECT 1.300 54.400 1.900 55.600 ;
        RECT 1.200 53.600 2.000 54.400 ;
        RECT 2.800 53.600 3.600 54.400 ;
        RECT 4.400 53.600 5.200 54.400 ;
        RECT 2.900 38.400 3.500 53.600 ;
        RECT 4.400 49.600 5.200 50.400 ;
        RECT 2.800 37.600 3.600 38.400 ;
        RECT 9.300 20.400 9.900 55.600 ;
        RECT 12.500 54.400 13.100 55.600 ;
        RECT 10.800 53.600 11.600 54.400 ;
        RECT 12.400 53.600 13.200 54.400 ;
        RECT 17.200 53.600 18.000 54.400 ;
        RECT 22.100 52.400 22.700 57.600 ;
        RECT 23.600 53.600 24.400 54.400 ;
        RECT 25.200 53.600 26.000 54.400 ;
        RECT 18.800 51.600 19.600 52.400 ;
        RECT 22.000 51.600 22.800 52.400 ;
        RECT 25.300 50.400 25.900 53.600 ;
        RECT 26.800 52.300 27.600 52.400 ;
        RECT 28.500 52.300 29.100 69.600 ;
        RECT 31.700 68.400 32.300 69.600 ;
        RECT 30.000 67.600 30.800 68.400 ;
        RECT 31.600 67.600 32.400 68.400 ;
        RECT 39.600 67.600 40.400 68.400 ;
        RECT 42.800 67.600 43.600 68.400 ;
        RECT 44.400 67.600 45.200 68.400 ;
        RECT 47.700 68.300 48.300 89.600 ;
        RECT 49.300 70.400 49.900 97.600 ;
        RECT 50.800 93.600 51.600 94.400 ;
        RECT 49.200 69.600 50.000 70.400 ;
        RECT 50.900 68.400 51.500 93.600 ;
        RECT 54.000 84.200 54.800 97.800 ;
        RECT 55.600 84.200 56.400 97.800 ;
        RECT 57.200 86.200 58.000 97.800 ;
        RECT 58.800 93.600 59.600 94.400 ;
        RECT 60.400 86.200 61.200 97.800 ;
        RECT 62.100 96.400 62.700 101.700 ;
        RECT 81.300 98.400 81.900 103.600 ;
        RECT 62.000 95.600 62.800 96.400 ;
        RECT 62.100 82.400 62.700 95.600 ;
        RECT 63.600 86.200 64.400 97.800 ;
        RECT 65.200 84.200 66.000 97.800 ;
        RECT 66.800 84.200 67.600 97.800 ;
        RECT 68.400 84.200 69.200 97.800 ;
        RECT 81.200 97.600 82.000 98.400 ;
        RECT 79.600 95.600 80.400 96.400 ;
        RECT 79.700 88.400 80.300 95.600 ;
        RECT 82.900 92.400 83.500 103.600 ;
        RECT 84.500 92.400 85.100 107.600 ;
        RECT 82.800 91.600 83.600 92.400 ;
        RECT 84.400 91.600 85.200 92.400 ;
        RECT 81.200 90.300 82.000 90.400 ;
        RECT 81.200 89.700 83.500 90.300 ;
        RECT 81.200 89.600 82.000 89.700 ;
        RECT 79.600 87.600 80.400 88.400 ;
        RECT 62.000 81.600 62.800 82.400 ;
        RECT 65.200 81.600 66.000 82.400 ;
        RECT 65.300 78.400 65.900 81.600 ;
        RECT 65.200 77.600 66.000 78.400 ;
        RECT 52.400 73.600 53.200 74.400 ;
        RECT 52.500 68.400 53.100 73.600 ;
        RECT 58.800 71.600 59.600 72.400 ;
        RECT 79.700 70.400 80.300 87.600 ;
        RECT 82.900 78.400 83.500 89.700 ;
        RECT 82.800 77.600 83.600 78.400 ;
        RECT 84.500 74.400 85.100 91.600 ;
        RECT 86.100 74.400 86.700 121.600 ;
        RECT 90.900 112.400 91.500 133.600 ;
        RECT 92.500 132.400 93.100 135.600 ;
        RECT 94.000 133.600 94.800 134.400 ;
        RECT 92.400 131.600 93.200 132.400 ;
        RECT 94.100 122.400 94.700 133.600 ;
        RECT 100.500 132.400 101.100 149.600 ;
        RECT 105.300 142.400 105.900 149.600 ;
        RECT 108.500 148.400 109.100 155.600 ;
        RECT 114.800 153.600 115.600 154.400 ;
        RECT 114.900 150.400 115.500 153.600 ;
        RECT 118.000 151.600 118.800 152.400 ;
        RECT 114.800 149.600 115.600 150.400 ;
        RECT 108.400 147.600 109.200 148.400 ;
        RECT 116.400 147.600 117.200 148.400 ;
        RECT 116.500 144.400 117.100 147.600 ;
        RECT 118.100 146.400 118.700 151.600 ;
        RECT 119.700 150.400 120.300 157.600 ;
        RECT 121.200 155.600 122.000 156.400 ;
        RECT 119.600 149.600 120.400 150.400 ;
        RECT 119.700 146.400 120.300 149.600 ;
        RECT 118.000 145.600 118.800 146.400 ;
        RECT 119.600 145.600 120.400 146.400 ;
        RECT 129.200 146.200 130.000 151.800 ;
        RECT 111.600 143.600 112.400 144.400 ;
        RECT 116.400 143.600 117.200 144.400 ;
        RECT 132.400 144.200 133.200 155.800 ;
        RECT 134.100 148.400 134.700 175.600 ;
        RECT 135.600 166.200 136.400 177.800 ;
        RECT 137.200 173.600 138.000 174.400 ;
        RECT 138.800 166.200 139.600 177.800 ;
        RECT 140.400 164.200 141.200 177.800 ;
        RECT 142.000 164.200 142.800 177.800 ;
        RECT 146.800 169.600 147.600 170.400 ;
        RECT 135.600 149.600 136.400 150.400 ;
        RECT 134.000 147.600 134.800 148.400 ;
        RECT 105.200 141.600 106.000 142.400 ;
        RECT 102.000 139.600 102.800 140.400 ;
        RECT 97.200 131.600 98.000 132.400 ;
        RECT 100.400 131.600 101.200 132.400 ;
        RECT 94.000 121.600 94.800 122.400 ;
        RECT 102.100 118.400 102.700 139.600 ;
        RECT 106.800 124.200 107.600 137.800 ;
        RECT 108.400 124.200 109.200 137.800 ;
        RECT 110.000 126.200 110.800 137.800 ;
        RECT 111.700 136.400 112.300 143.600 ;
        RECT 111.600 135.600 112.400 136.400 ;
        RECT 111.600 133.600 112.400 134.400 ;
        RECT 111.700 132.400 112.300 133.600 ;
        RECT 111.600 131.600 112.400 132.400 ;
        RECT 113.200 126.200 114.000 137.800 ;
        RECT 114.800 135.600 115.600 136.400 ;
        RECT 90.800 111.600 91.600 112.400 ;
        RECT 87.600 109.600 88.400 110.400 ;
        RECT 92.400 104.200 93.200 117.800 ;
        RECT 94.000 104.200 94.800 117.800 ;
        RECT 102.000 117.600 102.800 118.400 ;
        RECT 95.600 104.200 96.400 115.800 ;
        RECT 97.200 107.600 98.000 108.400 ;
        RECT 97.300 104.400 97.900 107.600 ;
        RECT 97.200 103.600 98.000 104.400 ;
        RECT 98.800 104.200 99.600 115.800 ;
        RECT 100.400 105.600 101.200 106.400 ;
        RECT 102.000 104.200 102.800 115.800 ;
        RECT 103.600 104.200 104.400 117.800 ;
        RECT 105.200 104.200 106.000 117.800 ;
        RECT 106.800 104.200 107.600 117.800 ;
        RECT 108.400 109.600 109.200 110.400 ;
        RECT 108.500 100.400 109.100 109.600 ;
        RECT 114.900 106.400 115.500 135.600 ;
        RECT 116.400 126.200 117.200 137.800 ;
        RECT 116.400 123.600 117.200 124.400 ;
        RECT 118.000 124.200 118.800 137.800 ;
        RECT 119.600 124.200 120.400 137.800 ;
        RECT 121.200 124.200 122.000 137.800 ;
        RECT 134.100 136.400 134.700 147.600 ;
        RECT 142.000 144.200 142.800 155.800 ;
        RECT 145.200 155.600 146.000 156.400 ;
        RECT 143.600 143.600 144.400 144.400 ;
        RECT 134.000 135.600 134.800 136.400 ;
        RECT 142.000 135.600 142.800 136.400 ;
        RECT 143.700 134.400 144.300 143.600 ;
        RECT 122.800 133.600 123.600 134.400 ;
        RECT 143.600 133.600 144.400 134.400 ;
        RECT 122.900 132.400 123.500 133.600 ;
        RECT 145.300 132.400 145.900 155.600 ;
        RECT 146.800 143.600 147.600 144.400 ;
        RECT 122.800 131.600 123.600 132.400 ;
        RECT 145.200 132.300 146.000 132.400 ;
        RECT 143.700 131.700 146.000 132.300 ;
        RECT 130.800 124.300 131.600 124.400 ;
        RECT 129.300 123.700 131.600 124.300 ;
        RECT 116.500 118.400 117.100 123.600 ;
        RECT 119.600 121.600 120.400 122.400 ;
        RECT 119.700 118.400 120.300 121.600 ;
        RECT 116.400 117.600 117.200 118.400 ;
        RECT 119.600 117.600 120.400 118.400 ;
        RECT 116.500 110.400 117.100 117.600 ;
        RECT 116.400 109.600 117.200 110.400 ;
        RECT 127.600 109.600 128.400 110.400 ;
        RECT 129.300 106.400 129.900 123.700 ;
        RECT 130.800 123.600 131.600 123.700 ;
        RECT 137.200 123.600 138.000 124.400 ;
        RECT 130.800 111.600 131.600 112.400 ;
        RECT 134.000 111.600 134.800 112.400 ;
        RECT 134.100 106.400 134.700 111.600 ;
        RECT 137.300 108.400 137.900 123.600 ;
        RECT 143.700 110.400 144.300 131.700 ;
        RECT 145.200 131.600 146.000 131.700 ;
        RECT 150.100 130.400 150.700 199.600 ;
        RECT 151.600 184.200 152.400 197.800 ;
        RECT 153.200 184.200 154.000 197.800 ;
        RECT 154.800 184.200 155.600 195.800 ;
        RECT 156.400 187.600 157.200 188.400 ;
        RECT 153.200 171.600 154.000 172.400 ;
        RECT 153.300 170.400 153.900 171.600 ;
        RECT 153.200 169.600 154.000 170.400 ;
        RECT 156.500 162.300 157.100 187.600 ;
        RECT 158.000 184.200 158.800 195.800 ;
        RECT 159.600 185.600 160.400 186.400 ;
        RECT 161.200 184.200 162.000 195.800 ;
        RECT 162.800 184.200 163.600 197.800 ;
        RECT 164.400 184.200 165.200 197.800 ;
        RECT 166.000 184.200 166.800 197.800 ;
        RECT 167.600 185.600 168.400 186.400 ;
        RECT 159.600 164.200 160.400 177.800 ;
        RECT 161.200 164.200 162.000 177.800 ;
        RECT 162.800 166.200 163.600 177.800 ;
        RECT 164.400 175.600 165.200 176.400 ;
        RECT 164.500 174.400 165.100 175.600 ;
        RECT 164.400 173.600 165.200 174.400 ;
        RECT 164.400 171.600 165.200 172.400 ;
        RECT 154.900 161.700 157.100 162.300 ;
        RECT 151.600 149.600 152.400 150.400 ;
        RECT 151.700 134.400 152.300 149.600 ;
        RECT 154.900 138.400 155.500 161.700 ;
        RECT 156.400 144.200 157.200 157.800 ;
        RECT 158.000 144.200 158.800 157.800 ;
        RECT 159.600 144.200 160.400 155.800 ;
        RECT 161.200 147.600 162.000 148.400 ;
        RECT 161.200 143.600 162.000 144.400 ;
        RECT 162.800 144.200 163.600 155.800 ;
        RECT 164.500 146.400 165.100 171.600 ;
        RECT 166.000 166.200 166.800 177.800 ;
        RECT 167.700 176.400 168.300 185.600 ;
        RECT 174.100 182.400 174.700 211.600 ;
        RECT 175.600 203.600 176.400 204.400 ;
        RECT 175.700 200.400 176.300 203.600 ;
        RECT 175.600 199.600 176.400 200.400 ;
        RECT 175.600 198.300 176.400 198.400 ;
        RECT 177.300 198.300 177.900 215.600 ;
        RECT 178.900 214.400 179.500 221.600 ;
        RECT 183.700 216.400 184.300 265.700 ;
        RECT 185.300 256.400 185.900 279.600 ;
        RECT 188.400 277.600 189.200 278.400 ;
        RECT 186.800 273.600 187.600 274.400 ;
        RECT 188.500 270.400 189.100 277.600 ;
        RECT 193.300 274.400 193.900 283.600 ;
        RECT 190.000 273.600 190.800 274.400 ;
        RECT 193.200 273.600 194.000 274.400 ;
        RECT 190.100 272.400 190.700 273.600 ;
        RECT 190.000 271.600 190.800 272.400 ;
        RECT 194.900 272.300 195.500 295.700 ;
        RECT 198.000 295.600 198.800 296.400 ;
        RECT 198.100 294.400 198.700 295.600 ;
        RECT 196.400 293.600 197.200 294.400 ;
        RECT 198.000 293.600 198.800 294.400 ;
        RECT 196.500 292.400 197.100 293.600 ;
        RECT 199.700 292.400 200.300 301.600 ;
        RECT 201.200 299.600 202.000 300.400 ;
        RECT 201.300 298.400 201.900 299.600 ;
        RECT 201.200 297.600 202.000 298.400 ;
        RECT 212.400 295.600 213.200 296.400 ;
        RECT 201.200 294.300 202.000 294.400 ;
        RECT 201.200 293.700 203.500 294.300 ;
        RECT 201.200 293.600 202.000 293.700 ;
        RECT 202.900 292.400 203.500 293.700 ;
        RECT 204.400 293.600 205.200 294.400 ;
        RECT 196.400 292.300 197.200 292.400 ;
        RECT 196.400 291.700 198.700 292.300 ;
        RECT 196.400 291.600 197.200 291.700 ;
        RECT 198.100 278.400 198.700 291.700 ;
        RECT 199.600 291.600 200.400 292.400 ;
        RECT 202.800 291.600 203.600 292.400 ;
        RECT 206.000 291.600 206.800 292.400 ;
        RECT 201.200 289.600 202.000 290.400 ;
        RECT 198.000 277.600 198.800 278.400 ;
        RECT 199.600 273.600 200.400 274.400 ;
        RECT 196.400 272.300 197.200 272.400 ;
        RECT 194.900 271.700 197.200 272.300 ;
        RECT 196.400 271.600 197.200 271.700 ;
        RECT 188.400 269.600 189.200 270.400 ;
        RECT 193.200 269.600 194.000 270.400 ;
        RECT 194.800 269.600 195.600 270.400 ;
        RECT 198.000 269.600 198.800 270.400 ;
        RECT 194.900 268.400 195.500 269.600 ;
        RECT 188.400 268.300 189.200 268.400 ;
        RECT 188.400 267.700 190.700 268.300 ;
        RECT 188.400 267.600 189.200 267.700 ;
        RECT 188.400 263.600 189.200 264.400 ;
        RECT 188.500 258.400 189.100 263.600 ;
        RECT 190.100 258.400 190.700 267.700 ;
        RECT 191.600 267.600 192.400 268.400 ;
        RECT 194.800 267.600 195.600 268.400 ;
        RECT 188.400 257.600 189.200 258.400 ;
        RECT 190.000 257.600 190.800 258.400 ;
        RECT 185.200 255.600 186.000 256.400 ;
        RECT 185.200 254.300 186.000 254.400 ;
        RECT 185.200 253.700 187.500 254.300 ;
        RECT 185.200 253.600 186.000 253.700 ;
        RECT 186.900 228.400 187.500 253.700 ;
        RECT 188.400 249.600 189.200 250.400 ;
        RECT 188.500 234.400 189.100 249.600 ;
        RECT 188.400 233.600 189.200 234.400 ;
        RECT 191.700 234.300 192.300 267.600 ;
        RECT 193.200 265.600 194.000 266.400 ;
        RECT 193.300 258.400 193.900 265.600 ;
        RECT 201.300 260.300 201.900 289.600 ;
        RECT 202.900 272.400 203.500 291.600 ;
        RECT 206.100 276.400 206.700 291.600 ;
        RECT 207.600 289.600 208.400 290.400 ;
        RECT 207.600 277.600 208.400 278.400 ;
        RECT 206.000 275.600 206.800 276.400 ;
        RECT 210.800 273.600 211.600 274.400 ;
        RECT 202.800 271.600 203.600 272.400 ;
        RECT 209.200 271.600 210.000 272.400 ;
        RECT 209.300 270.400 209.900 271.600 ;
        RECT 202.800 269.600 203.600 270.400 ;
        RECT 209.200 269.600 210.000 270.400 ;
        RECT 210.800 269.600 211.600 270.400 ;
        RECT 212.500 270.300 213.100 295.600 ;
        RECT 214.000 294.300 214.800 294.400 ;
        RECT 215.700 294.300 216.300 311.600 ;
        RECT 222.100 310.400 222.700 311.600 ;
        RECT 222.000 309.600 222.800 310.400 ;
        RECT 226.900 308.400 227.500 317.600 ;
        RECT 230.000 315.600 230.800 316.400 ;
        RECT 228.400 311.600 229.200 312.400 ;
        RECT 226.800 307.600 227.600 308.400 ;
        RECT 220.400 305.600 221.200 306.400 ;
        RECT 217.200 303.600 218.000 304.400 ;
        RECT 218.800 303.600 219.600 304.400 ;
        RECT 217.300 294.400 217.900 303.600 ;
        RECT 218.900 296.400 219.500 303.600 ;
        RECT 220.500 298.400 221.100 305.600 ;
        RECT 228.400 303.600 229.200 304.400 ;
        RECT 220.400 297.600 221.200 298.400 ;
        RECT 218.800 295.600 219.600 296.400 ;
        RECT 228.500 296.300 229.100 303.600 ;
        RECT 230.100 298.400 230.700 315.600 ;
        RECT 233.300 312.400 233.900 319.600 ;
        RECT 236.500 316.400 237.100 335.600 ;
        RECT 238.000 326.200 238.800 337.800 ;
        RECT 239.600 333.600 240.400 334.400 ;
        RECT 241.200 326.200 242.000 337.800 ;
        RECT 242.800 324.200 243.600 337.800 ;
        RECT 244.400 324.200 245.200 337.800 ;
        RECT 247.700 336.400 248.300 353.600 ;
        RECT 249.300 350.400 249.900 355.600 ;
        RECT 254.100 354.400 254.700 355.600 ;
        RECT 254.000 353.600 254.800 354.400 ;
        RECT 255.700 352.400 256.300 365.600 ;
        RECT 263.600 364.200 264.400 377.800 ;
        RECT 265.200 364.200 266.000 377.800 ;
        RECT 266.800 364.200 267.600 377.800 ;
        RECT 268.400 366.200 269.200 377.800 ;
        RECT 270.000 375.600 270.800 376.400 ;
        RECT 270.100 352.400 270.700 375.600 ;
        RECT 271.600 366.200 272.400 377.800 ;
        RECT 273.200 375.600 274.000 376.400 ;
        RECT 273.300 374.400 273.900 375.600 ;
        RECT 273.200 373.600 274.000 374.400 ;
        RECT 274.800 366.200 275.600 377.800 ;
        RECT 276.400 364.200 277.200 377.800 ;
        RECT 278.000 364.200 278.800 377.800 ;
        RECT 327.600 377.600 328.400 378.400 ;
        RECT 342.000 377.600 342.800 378.400 ;
        RECT 302.000 375.600 302.800 376.400 ;
        RECT 314.800 375.600 315.600 376.400 ;
        RECT 295.600 373.600 296.400 374.400 ;
        RECT 298.800 373.600 299.600 374.400 ;
        RECT 300.400 373.600 301.200 374.400 ;
        RECT 306.800 373.600 307.600 374.400 ;
        RECT 319.600 373.600 320.400 374.400 ;
        RECT 298.900 372.400 299.500 373.600 ;
        RECT 281.200 371.600 282.000 372.400 ;
        RECT 297.200 371.600 298.000 372.400 ;
        RECT 298.800 371.600 299.600 372.400 ;
        RECT 250.800 351.600 251.600 352.400 ;
        RECT 255.600 351.600 256.400 352.400 ;
        RECT 257.200 351.600 258.000 352.400 ;
        RECT 266.800 351.600 267.600 352.400 ;
        RECT 270.000 351.600 270.800 352.400 ;
        RECT 255.700 350.400 256.300 351.600 ;
        RECT 249.200 349.600 250.000 350.400 ;
        RECT 255.600 349.600 256.400 350.400 ;
        RECT 257.300 348.400 257.900 351.600 ;
        RECT 257.200 347.600 258.000 348.400 ;
        RECT 265.200 343.600 266.000 344.400 ;
        RECT 265.300 338.400 265.900 343.600 ;
        RECT 265.200 337.600 266.000 338.400 ;
        RECT 247.600 335.600 248.400 336.400 ;
        RECT 255.600 333.600 256.400 334.400 ;
        RECT 244.400 321.600 245.200 322.400 ;
        RECT 244.500 318.400 245.100 321.600 ;
        RECT 238.000 317.600 238.800 318.400 ;
        RECT 244.400 317.600 245.200 318.400 ;
        RECT 236.400 315.600 237.200 316.400 ;
        RECT 233.200 311.600 234.000 312.400 ;
        RECT 236.400 309.600 237.200 310.400 ;
        RECT 238.100 308.400 238.700 317.600 ;
        RECT 247.600 311.600 248.400 312.400 ;
        RECT 244.400 309.600 245.200 310.400 ;
        RECT 238.000 307.600 238.800 308.400 ;
        RECT 238.000 305.600 238.800 306.400 ;
        RECT 238.100 298.400 238.700 305.600 ;
        RECT 230.000 297.600 230.800 298.400 ;
        RECT 238.000 297.600 238.800 298.400 ;
        RECT 242.800 297.600 243.600 298.400 ;
        RECT 226.900 295.700 229.100 296.300 ;
        RECT 214.000 293.700 216.300 294.300 ;
        RECT 214.000 293.600 214.800 293.700 ;
        RECT 214.000 289.600 214.800 290.400 ;
        RECT 214.000 270.300 214.800 270.400 ;
        RECT 212.500 269.700 214.800 270.300 ;
        RECT 214.000 269.600 214.800 269.700 ;
        RECT 204.400 265.600 205.200 266.400 ;
        RECT 206.000 265.600 206.800 266.400 ;
        RECT 199.700 259.700 201.900 260.300 ;
        RECT 193.200 257.600 194.000 258.400 ;
        RECT 193.300 250.400 193.900 257.600 ;
        RECT 199.700 256.400 200.300 259.700 ;
        RECT 201.200 257.600 202.000 258.400 ;
        RECT 194.800 255.600 195.600 256.400 ;
        RECT 199.600 256.300 200.400 256.400 ;
        RECT 198.100 255.700 200.400 256.300 ;
        RECT 193.200 249.600 194.000 250.400 ;
        RECT 194.900 238.400 195.500 255.600 ;
        RECT 198.100 252.400 198.700 255.700 ;
        RECT 199.600 255.600 200.400 255.700 ;
        RECT 201.300 254.400 201.900 257.600 ;
        RECT 201.200 253.600 202.000 254.400 ;
        RECT 198.000 251.600 198.800 252.400 ;
        RECT 194.800 237.600 195.600 238.400 ;
        RECT 204.500 234.400 205.100 265.600 ;
        RECT 207.600 257.600 208.400 258.400 ;
        RECT 209.300 256.400 209.900 269.600 ;
        RECT 210.900 266.400 211.500 269.600 ;
        RECT 215.700 268.400 216.300 293.700 ;
        RECT 217.200 293.600 218.000 294.400 ;
        RECT 220.400 293.600 221.200 294.400 ;
        RECT 223.600 293.600 224.400 294.400 ;
        RECT 220.500 292.400 221.100 293.600 ;
        RECT 226.900 292.400 227.500 295.700 ;
        RECT 234.800 295.600 235.600 296.400 ;
        RECT 228.400 293.600 229.200 294.400 ;
        RECT 231.600 293.600 232.400 294.400 ;
        RECT 228.500 292.400 229.100 293.600 ;
        RECT 234.900 292.400 235.500 295.600 ;
        RECT 242.900 294.400 243.500 297.600 ;
        RECT 236.400 293.600 237.200 294.400 ;
        RECT 239.600 293.600 240.400 294.400 ;
        RECT 242.800 293.600 243.600 294.400 ;
        RECT 236.500 292.400 237.100 293.600 ;
        RECT 220.400 291.600 221.200 292.400 ;
        RECT 225.200 291.600 226.000 292.400 ;
        RECT 226.800 291.600 227.600 292.400 ;
        RECT 228.400 291.600 229.200 292.400 ;
        RECT 233.200 291.600 234.000 292.400 ;
        RECT 234.800 291.600 235.600 292.400 ;
        RECT 236.400 291.600 237.200 292.400 ;
        RECT 225.300 280.400 225.900 291.600 ;
        RECT 233.300 290.400 233.900 291.600 ;
        RECT 233.200 289.600 234.000 290.400 ;
        RECT 231.600 287.600 232.400 288.400 ;
        RECT 225.200 279.600 226.000 280.400 ;
        RECT 220.400 271.600 221.200 272.400 ;
        RECT 225.200 271.600 226.000 272.400 ;
        RECT 215.600 267.600 216.400 268.400 ;
        RECT 220.500 266.400 221.100 271.600 ;
        RECT 231.700 270.400 232.300 287.600 ;
        RECT 234.800 273.600 235.600 274.400 ;
        RECT 234.900 272.400 235.500 273.600 ;
        RECT 234.800 271.600 235.600 272.400 ;
        RECT 236.500 272.300 237.100 291.600 ;
        RECT 239.700 290.300 240.300 293.600 ;
        RECT 244.500 292.400 245.100 309.600 ;
        RECT 247.700 306.400 248.300 311.600 ;
        RECT 249.200 309.600 250.000 310.400 ;
        RECT 247.600 305.600 248.400 306.400 ;
        RECT 246.000 297.600 246.800 298.400 ;
        RECT 241.200 291.600 242.000 292.400 ;
        RECT 244.400 291.600 245.200 292.400 ;
        RECT 239.700 289.700 241.900 290.300 ;
        RECT 238.000 273.600 238.800 274.400 ;
        RECT 236.500 271.700 238.700 272.300 ;
        RECT 226.800 269.600 227.600 270.400 ;
        RECT 231.600 269.600 232.400 270.400 ;
        RECT 236.400 269.600 237.200 270.400 ;
        RECT 231.700 268.400 232.300 269.600 ;
        RECT 238.100 268.400 238.700 271.700 ;
        RECT 241.300 268.400 241.900 289.700 ;
        RECT 244.500 288.400 245.100 291.600 ;
        RECT 244.400 287.600 245.200 288.400 ;
        RECT 242.800 273.600 243.600 274.400 ;
        RECT 242.900 270.400 243.500 273.600 ;
        RECT 242.800 269.600 243.600 270.400 ;
        RECT 231.600 267.600 232.400 268.400 ;
        RECT 238.000 267.600 238.800 268.400 ;
        RECT 241.200 267.600 242.000 268.400 ;
        RECT 244.400 267.600 245.200 268.400 ;
        RECT 210.800 265.600 211.600 266.400 ;
        RECT 214.000 265.600 214.800 266.400 ;
        RECT 220.400 265.600 221.200 266.400 ;
        RECT 226.800 265.600 227.600 266.400 ;
        RECT 214.100 258.400 214.700 265.600 ;
        RECT 234.800 263.600 235.600 264.400 ;
        RECT 214.000 257.600 214.800 258.400 ;
        RECT 206.000 255.600 206.800 256.400 ;
        RECT 209.200 255.600 210.000 256.400 ;
        RECT 217.200 244.200 218.000 257.800 ;
        RECT 218.800 244.200 219.600 257.800 ;
        RECT 220.400 244.200 221.200 257.800 ;
        RECT 222.000 246.200 222.800 257.800 ;
        RECT 223.600 255.600 224.400 256.400 ;
        RECT 223.700 254.400 224.300 255.600 ;
        RECT 223.600 253.600 224.400 254.400 ;
        RECT 212.400 241.600 213.200 242.400 ;
        RECT 190.100 233.700 192.300 234.300 ;
        RECT 190.100 232.400 190.700 233.700 ;
        RECT 194.800 233.600 195.600 234.400 ;
        RECT 204.400 233.600 205.200 234.400 ;
        RECT 190.000 231.600 190.800 232.400 ;
        RECT 191.600 231.600 192.400 232.400 ;
        RECT 194.900 230.400 195.500 233.600 ;
        RECT 202.800 231.600 203.600 232.400 ;
        RECT 209.200 231.600 210.000 232.400 ;
        RECT 191.600 229.600 192.400 230.400 ;
        RECT 194.800 229.600 195.600 230.400 ;
        RECT 199.600 229.600 200.400 230.400 ;
        RECT 186.800 227.600 187.600 228.400 ;
        RECT 196.400 227.600 197.200 228.400 ;
        RECT 198.000 227.600 198.800 228.400 ;
        RECT 186.900 224.400 187.500 227.600 ;
        RECT 186.800 223.600 187.600 224.400 ;
        RECT 196.500 222.400 197.100 227.600 ;
        RECT 204.400 225.600 205.200 226.400 ;
        RECT 206.000 223.600 206.800 224.400 ;
        RECT 185.200 221.600 186.000 222.400 ;
        RECT 196.400 221.600 197.200 222.400 ;
        RECT 183.600 215.600 184.400 216.400 ;
        RECT 178.800 213.600 179.600 214.400 ;
        RECT 185.300 212.400 185.900 221.600 ;
        RECT 199.600 219.600 200.400 220.400 ;
        RECT 188.400 215.600 189.200 216.400 ;
        RECT 194.800 215.600 195.600 216.400 ;
        RECT 188.500 214.400 189.100 215.600 ;
        RECT 188.400 213.600 189.200 214.400 ;
        RECT 180.400 211.600 181.200 212.400 ;
        RECT 183.600 211.600 184.400 212.400 ;
        RECT 185.200 211.600 186.000 212.400 ;
        RECT 191.600 211.600 192.400 212.400 ;
        RECT 180.500 198.400 181.100 211.600 ;
        RECT 194.900 210.400 195.500 215.600 ;
        RECT 199.700 214.400 200.300 219.600 ;
        RECT 201.200 215.600 202.000 216.400 ;
        RECT 196.400 213.600 197.200 214.400 ;
        RECT 199.600 213.600 200.400 214.400 ;
        RECT 198.000 211.600 198.800 212.400 ;
        RECT 199.700 210.400 200.300 213.600 ;
        RECT 194.800 209.600 195.600 210.400 ;
        RECT 199.600 209.600 200.400 210.400 ;
        RECT 191.600 207.600 192.400 208.400 ;
        RECT 201.300 206.300 201.900 215.600 ;
        RECT 204.400 211.600 205.200 212.400 ;
        RECT 206.100 212.300 206.700 223.600 ;
        RECT 209.300 218.400 209.900 231.600 ;
        RECT 212.500 228.400 213.100 241.600 ;
        RECT 223.700 238.300 224.300 253.600 ;
        RECT 225.200 246.200 226.000 257.800 ;
        RECT 226.800 253.600 227.600 254.400 ;
        RECT 228.400 246.200 229.200 257.800 ;
        RECT 230.000 244.200 230.800 257.800 ;
        RECT 231.600 244.200 232.400 257.800 ;
        RECT 234.900 254.400 235.500 263.600 ;
        RECT 234.800 253.600 235.600 254.400 ;
        RECT 233.200 251.600 234.000 252.400 ;
        RECT 212.400 227.600 213.200 228.400 ;
        RECT 209.200 217.600 210.000 218.400 ;
        RECT 212.500 214.400 213.100 227.600 ;
        RECT 215.600 224.200 216.400 237.800 ;
        RECT 217.200 224.200 218.000 237.800 ;
        RECT 218.800 224.200 219.600 237.800 ;
        RECT 222.100 237.700 224.300 238.300 ;
        RECT 220.400 224.200 221.200 235.800 ;
        RECT 222.100 226.400 222.700 237.700 ;
        RECT 222.000 225.600 222.800 226.400 ;
        RECT 220.400 221.600 221.200 222.400 ;
        RECT 220.500 214.400 221.100 221.600 ;
        RECT 222.100 216.400 222.700 225.600 ;
        RECT 223.600 224.200 224.400 235.800 ;
        RECT 225.200 227.600 226.000 228.400 ;
        RECT 225.300 226.400 225.900 227.600 ;
        RECT 225.200 225.600 226.000 226.400 ;
        RECT 226.800 224.200 227.600 235.800 ;
        RECT 228.400 224.200 229.200 237.800 ;
        RECT 230.000 224.200 230.800 237.800 ;
        RECT 233.300 230.400 233.900 251.600 ;
        RECT 241.300 250.400 241.900 267.600 ;
        RECT 244.500 266.400 245.100 267.600 ;
        RECT 242.800 265.600 243.600 266.400 ;
        RECT 244.400 265.600 245.200 266.400 ;
        RECT 242.900 258.400 243.500 265.600 ;
        RECT 242.800 257.600 243.600 258.400 ;
        RECT 241.200 249.600 242.000 250.400 ;
        RECT 241.300 242.400 241.900 249.600 ;
        RECT 241.200 241.600 242.000 242.400 ;
        RECT 233.200 229.600 234.000 230.400 ;
        RECT 234.800 229.600 235.600 230.400 ;
        RECT 244.500 226.400 245.100 265.600 ;
        RECT 246.100 262.400 246.700 297.600 ;
        RECT 249.300 296.400 249.900 309.600 ;
        RECT 250.800 303.600 251.600 304.400 ;
        RECT 255.700 298.400 256.300 333.600 ;
        RECT 258.800 303.600 259.600 304.400 ;
        RECT 260.400 304.200 261.200 317.800 ;
        RECT 262.000 304.200 262.800 317.800 ;
        RECT 263.600 304.200 264.400 317.800 ;
        RECT 266.900 316.400 267.500 351.600 ;
        RECT 268.400 349.600 269.200 350.400 ;
        RECT 270.000 349.600 270.800 350.400 ;
        RECT 265.200 304.200 266.000 315.800 ;
        RECT 266.800 315.600 267.600 316.400 ;
        RECT 266.900 306.400 267.500 315.600 ;
        RECT 266.800 305.600 267.600 306.400 ;
        RECT 255.600 297.600 256.400 298.400 ;
        RECT 258.900 296.400 259.500 303.600 ;
        RECT 266.900 296.400 267.500 305.600 ;
        RECT 268.400 304.200 269.200 315.800 ;
        RECT 270.100 310.400 270.700 349.600 ;
        RECT 273.200 344.200 274.000 357.800 ;
        RECT 274.800 344.200 275.600 357.800 ;
        RECT 276.400 344.200 277.200 355.800 ;
        RECT 278.000 347.600 278.800 348.400 ;
        RECT 278.100 346.400 278.700 347.600 ;
        RECT 278.000 345.600 278.800 346.400 ;
        RECT 279.600 344.200 280.400 355.800 ;
        RECT 281.300 354.400 281.900 371.600 ;
        RECT 297.300 370.400 297.900 371.600 ;
        RECT 297.200 369.600 298.000 370.400 ;
        RECT 292.400 367.600 293.200 368.400 ;
        RECT 292.500 364.400 293.100 367.600 ;
        RECT 292.400 363.600 293.200 364.400 ;
        RECT 298.900 362.400 299.500 371.600 ;
        RECT 303.600 369.600 304.400 370.400 ;
        RECT 298.800 361.600 299.600 362.400 ;
        RECT 302.000 359.600 302.800 360.400 ;
        RECT 281.200 353.600 282.000 354.400 ;
        RECT 281.200 345.600 282.000 346.400 ;
        RECT 281.300 344.400 281.900 345.600 ;
        RECT 281.200 343.600 282.000 344.400 ;
        RECT 282.800 344.200 283.600 355.800 ;
        RECT 284.400 344.200 285.200 357.800 ;
        RECT 286.000 344.200 286.800 357.800 ;
        RECT 287.600 344.200 288.400 357.800 ;
        RECT 302.100 354.400 302.700 359.600 ;
        RECT 303.700 358.400 304.300 369.600 ;
        RECT 305.200 365.600 306.000 366.400 ;
        RECT 305.300 364.400 305.900 365.600 ;
        RECT 305.200 363.600 306.000 364.400 ;
        RECT 303.600 357.600 304.400 358.400 ;
        RECT 303.600 355.600 304.400 356.400 ;
        RECT 302.000 353.600 302.800 354.400 ;
        RECT 303.700 352.400 304.300 355.600 ;
        RECT 305.300 352.400 305.900 363.600 ;
        RECT 306.900 362.400 307.500 373.600 ;
        RECT 327.700 372.400 328.300 377.600 ;
        RECT 342.100 376.400 342.700 377.600 ;
        RECT 330.800 375.600 331.600 376.400 ;
        RECT 335.600 375.600 336.400 376.400 ;
        RECT 342.000 375.600 342.800 376.400 ;
        RECT 310.000 371.600 310.800 372.400 ;
        RECT 314.800 371.600 315.600 372.400 ;
        RECT 318.000 371.600 318.800 372.400 ;
        RECT 319.600 371.600 320.400 372.400 ;
        RECT 322.800 371.600 323.600 372.400 ;
        RECT 327.600 371.600 328.400 372.400 ;
        RECT 308.400 369.600 309.200 370.400 ;
        RECT 308.500 366.400 309.100 369.600 ;
        RECT 310.000 367.600 310.800 368.400 ;
        RECT 313.200 367.600 314.000 368.400 ;
        RECT 308.400 365.600 309.200 366.400 ;
        RECT 306.800 361.600 307.600 362.400 ;
        RECT 310.100 356.400 310.700 367.600 ;
        RECT 311.600 365.600 312.400 366.400 ;
        RECT 311.700 358.400 312.300 365.600 ;
        RECT 311.600 357.600 312.400 358.400 ;
        RECT 310.000 355.600 310.800 356.400 ;
        RECT 311.600 353.600 312.400 354.400 ;
        RECT 303.600 351.600 304.400 352.400 ;
        RECT 305.200 351.600 306.000 352.400 ;
        RECT 303.700 350.400 304.300 351.600 ;
        RECT 297.200 349.600 298.200 350.400 ;
        RECT 303.600 349.600 304.400 350.400 ;
        RECT 306.800 349.600 307.600 350.400 ;
        RECT 310.000 349.600 310.800 350.400 ;
        RECT 306.900 344.400 307.500 349.600 ;
        RECT 310.000 345.600 310.800 346.400 ;
        RECT 290.800 343.600 291.600 344.400 ;
        RECT 306.800 343.600 307.600 344.400 ;
        RECT 290.900 338.400 291.500 343.600 ;
        RECT 281.200 331.600 282.000 332.400 ;
        RECT 270.000 309.600 270.800 310.400 ;
        RECT 270.000 307.600 270.800 308.400 ;
        RECT 270.100 298.400 270.700 307.600 ;
        RECT 271.600 304.200 272.400 315.800 ;
        RECT 273.200 304.200 274.000 317.800 ;
        RECT 274.800 304.200 275.600 317.800 ;
        RECT 281.300 310.400 281.900 331.600 ;
        RECT 282.800 324.200 283.600 337.800 ;
        RECT 284.400 324.200 285.200 337.800 ;
        RECT 286.000 326.200 286.800 337.800 ;
        RECT 287.600 333.600 288.400 334.400 ;
        RECT 287.700 318.400 288.300 333.600 ;
        RECT 289.200 326.200 290.000 337.800 ;
        RECT 290.800 337.600 291.600 338.400 ;
        RECT 290.900 336.400 291.500 337.600 ;
        RECT 290.800 335.600 291.600 336.400 ;
        RECT 292.400 326.200 293.200 337.800 ;
        RECT 294.000 324.200 294.800 337.800 ;
        RECT 295.600 324.200 296.400 337.800 ;
        RECT 297.200 324.200 298.000 337.800 ;
        RECT 306.900 326.400 307.500 343.600 ;
        RECT 308.400 337.600 309.200 338.400 ;
        RECT 306.800 325.600 307.600 326.400 ;
        RECT 306.800 323.600 307.600 324.400 ;
        RECT 306.900 320.400 307.500 323.600 ;
        RECT 306.800 319.600 307.600 320.400 ;
        RECT 287.600 317.600 288.400 318.400 ;
        RECT 281.200 309.600 282.000 310.400 ;
        RECT 270.000 297.600 270.800 298.400 ;
        RECT 249.200 295.600 250.000 296.400 ;
        RECT 257.200 295.600 258.000 296.400 ;
        RECT 258.800 295.600 259.600 296.400 ;
        RECT 266.800 295.600 267.600 296.400 ;
        RECT 254.000 293.600 254.800 294.400 ;
        RECT 249.200 291.600 250.000 292.400 ;
        RECT 247.600 289.600 248.400 290.400 ;
        RECT 247.700 266.400 248.300 289.600 ;
        RECT 250.800 283.600 251.600 284.400 ;
        RECT 250.900 270.400 251.500 283.600 ;
        RECT 254.100 282.400 254.700 293.600 ;
        RECT 254.000 281.600 254.800 282.400 ;
        RECT 257.300 278.400 257.900 295.600 ;
        RECT 263.600 291.600 264.400 292.400 ;
        RECT 266.800 289.600 267.600 290.400 ;
        RECT 276.400 283.600 277.200 284.400 ;
        RECT 281.300 280.400 281.900 309.600 ;
        RECT 292.400 303.600 293.200 304.400 ;
        RECT 302.000 304.200 302.800 317.800 ;
        RECT 303.600 304.200 304.400 317.800 ;
        RECT 305.200 304.200 306.000 317.800 ;
        RECT 306.800 304.200 307.600 315.800 ;
        RECT 308.500 306.400 309.100 337.600 ;
        RECT 310.100 332.400 310.700 345.600 ;
        RECT 311.700 332.400 312.300 353.600 ;
        RECT 314.900 352.400 315.500 371.600 ;
        RECT 319.700 358.400 320.300 371.600 ;
        RECT 326.000 369.600 326.800 370.400 ;
        RECT 327.600 369.600 328.400 370.400 ;
        RECT 329.200 369.600 330.000 370.400 ;
        RECT 321.200 365.600 322.000 366.400 ;
        RECT 319.600 357.600 320.400 358.400 ;
        RECT 321.300 354.400 321.900 365.600 ;
        RECT 326.100 358.400 326.700 369.600 ;
        RECT 327.700 366.400 328.300 369.600 ;
        RECT 329.300 368.400 329.900 369.600 ;
        RECT 329.200 367.600 330.000 368.400 ;
        RECT 327.600 365.600 328.400 366.400 ;
        RECT 324.400 357.600 325.200 358.400 ;
        RECT 326.000 357.600 326.800 358.400 ;
        RECT 324.500 354.400 325.100 357.600 ;
        RECT 321.200 353.600 322.000 354.400 ;
        RECT 322.800 353.600 323.600 354.400 ;
        RECT 324.400 353.600 325.200 354.400 ;
        RECT 314.800 351.600 315.600 352.400 ;
        RECT 321.200 351.600 322.000 352.400 ;
        RECT 321.300 350.400 321.900 351.600 ;
        RECT 314.800 349.600 315.600 350.400 ;
        RECT 321.200 349.600 322.000 350.400 ;
        RECT 322.900 348.400 323.500 353.600 ;
        RECT 327.600 351.600 328.400 352.400 ;
        RECT 326.000 349.600 326.800 350.400 ;
        RECT 318.000 347.600 318.800 348.400 ;
        RECT 322.800 347.600 323.600 348.400 ;
        RECT 318.100 346.400 318.700 347.600 ;
        RECT 318.000 345.600 318.800 346.400 ;
        RECT 326.100 344.400 326.700 349.600 ;
        RECT 326.000 343.600 326.800 344.400 ;
        RECT 327.700 340.400 328.300 351.600 ;
        RECT 330.900 350.400 331.500 375.600 ;
        RECT 335.700 374.400 336.300 375.600 ;
        RECT 335.600 373.600 336.400 374.400 ;
        RECT 337.200 373.600 338.000 374.400 ;
        RECT 340.400 373.600 341.200 374.400 ;
        RECT 346.800 373.600 347.600 374.400 ;
        RECT 337.200 371.600 338.000 372.400 ;
        RECT 345.200 371.600 346.000 372.400 ;
        RECT 337.300 370.400 337.900 371.600 ;
        RECT 332.400 369.600 333.200 370.400 ;
        RECT 334.000 369.600 334.800 370.400 ;
        RECT 337.200 369.600 338.000 370.400 ;
        RECT 332.500 368.400 333.100 369.600 ;
        RECT 332.400 367.600 333.200 368.400 ;
        RECT 346.900 358.400 347.500 373.600 ;
        RECT 351.600 369.600 352.400 370.400 ;
        RECT 351.700 366.400 352.300 369.600 ;
        RECT 351.600 365.600 352.400 366.400 ;
        RECT 356.400 364.200 357.200 377.800 ;
        RECT 358.000 364.200 358.800 377.800 ;
        RECT 359.600 366.200 360.400 377.800 ;
        RECT 361.200 373.600 362.000 374.400 ;
        RECT 362.800 366.200 363.600 377.800 ;
        RECT 364.400 375.600 365.200 376.400 ;
        RECT 364.500 364.400 365.100 375.600 ;
        RECT 366.000 366.200 366.800 377.800 ;
        RECT 364.400 363.600 365.200 364.400 ;
        RECT 367.600 364.200 368.400 377.800 ;
        RECT 369.200 364.200 370.000 377.800 ;
        RECT 370.800 364.200 371.600 377.800 ;
        RECT 388.400 377.600 389.200 378.400 ;
        RECT 386.800 373.600 387.600 374.400 ;
        RECT 393.200 373.600 394.000 374.400 ;
        RECT 386.900 372.400 387.500 373.600 ;
        RECT 382.000 371.600 382.800 372.400 ;
        RECT 386.800 371.600 387.600 372.400 ;
        RECT 391.600 371.600 392.400 372.400 ;
        RECT 399.600 371.600 400.400 372.400 ;
        RECT 380.400 363.600 381.200 364.400 ;
        RECT 361.200 361.600 362.000 362.400 ;
        RECT 369.200 361.600 370.000 362.400 ;
        RECT 361.300 358.400 361.900 361.600 ;
        RECT 369.300 358.400 369.900 361.600 ;
        RECT 346.800 357.600 347.600 358.400 ;
        RECT 361.200 357.600 362.000 358.400 ;
        RECT 369.200 357.600 370.000 358.400 ;
        RECT 372.400 357.600 373.200 358.400 ;
        RECT 337.200 353.600 338.000 354.400 ;
        RECT 338.800 353.600 339.600 354.400 ;
        RECT 337.300 352.400 337.900 353.600 ;
        RECT 372.500 352.400 373.100 357.600 ;
        RECT 378.800 355.600 379.600 356.400 ;
        RECT 375.600 353.600 376.400 354.400 ;
        RECT 378.800 353.600 379.600 354.400 ;
        RECT 337.200 351.600 338.000 352.400 ;
        RECT 340.400 351.600 341.200 352.400 ;
        RECT 356.400 351.600 357.200 352.400 ;
        RECT 372.400 351.600 373.200 352.400 ;
        RECT 330.800 349.600 331.600 350.400 ;
        RECT 334.000 349.600 334.800 350.400 ;
        RECT 337.200 349.600 338.000 350.400 ;
        RECT 338.800 349.600 339.600 350.400 ;
        RECT 332.400 347.600 333.200 348.400 ;
        RECT 329.200 345.600 330.000 346.400 ;
        RECT 329.300 344.400 329.900 345.600 ;
        RECT 329.200 343.600 330.000 344.400 ;
        RECT 332.500 344.300 333.100 347.600 ;
        RECT 334.100 346.400 334.700 349.600 ;
        RECT 337.300 348.400 337.900 349.600 ;
        RECT 338.900 348.400 339.500 349.600 ;
        RECT 337.200 347.600 338.000 348.400 ;
        RECT 338.800 347.600 339.600 348.400 ;
        RECT 340.500 346.400 341.100 351.600 ;
        RECT 342.000 349.600 342.800 350.400 ;
        RECT 346.800 349.600 347.600 350.400 ;
        RECT 353.200 349.600 354.000 350.400 ;
        RECT 334.000 345.600 334.800 346.400 ;
        RECT 340.400 345.600 341.200 346.400 ;
        RECT 332.500 343.700 334.700 344.300 ;
        RECT 327.600 339.600 328.400 340.400 ;
        RECT 310.000 331.600 310.800 332.400 ;
        RECT 311.600 331.600 312.400 332.400 ;
        RECT 314.800 331.600 315.600 332.400 ;
        RECT 314.900 322.400 315.500 331.600 ;
        RECT 318.000 324.200 318.800 337.800 ;
        RECT 319.600 324.200 320.400 337.800 ;
        RECT 321.200 326.200 322.000 337.800 ;
        RECT 322.800 333.600 323.600 334.400 ;
        RECT 314.800 321.600 315.600 322.400 ;
        RECT 318.000 321.600 318.800 322.400 ;
        RECT 308.400 305.600 309.200 306.400 ;
        RECT 292.500 298.400 293.100 303.600 ;
        RECT 305.200 301.600 306.000 302.400 ;
        RECT 286.000 284.200 286.800 297.800 ;
        RECT 287.600 284.200 288.400 297.800 ;
        RECT 289.200 284.200 290.000 297.800 ;
        RECT 290.800 286.200 291.600 297.800 ;
        RECT 292.400 297.600 293.200 298.400 ;
        RECT 292.400 295.600 293.200 296.400 ;
        RECT 294.000 286.200 294.800 297.800 ;
        RECT 295.600 295.600 296.400 296.400 ;
        RECT 295.700 294.400 296.300 295.600 ;
        RECT 295.600 293.600 296.400 294.400 ;
        RECT 297.200 286.200 298.000 297.800 ;
        RECT 298.800 284.200 299.600 297.800 ;
        RECT 300.400 284.200 301.200 297.800 ;
        RECT 305.300 292.400 305.900 301.600 ;
        RECT 305.200 291.600 306.000 292.400 ;
        RECT 281.200 279.600 282.000 280.400 ;
        RECT 295.600 279.600 296.400 280.400 ;
        RECT 257.200 277.600 258.000 278.400 ;
        RECT 252.400 271.600 253.200 272.400 ;
        RECT 255.600 271.600 256.400 272.400 ;
        RECT 255.700 270.400 256.300 271.600 ;
        RECT 249.200 269.600 250.000 270.400 ;
        RECT 250.800 269.600 251.600 270.400 ;
        RECT 254.000 269.600 254.800 270.400 ;
        RECT 255.600 269.600 256.400 270.400 ;
        RECT 258.800 269.600 259.600 270.400 ;
        RECT 249.300 266.400 249.900 269.600 ;
        RECT 254.100 268.400 254.700 269.600 ;
        RECT 254.000 267.600 254.800 268.400 ;
        RECT 247.600 265.600 248.400 266.400 ;
        RECT 249.200 265.600 250.000 266.400 ;
        RECT 246.000 261.600 246.800 262.400 ;
        RECT 247.600 243.600 248.400 244.400 ;
        RECT 239.600 226.300 240.400 226.400 ;
        RECT 238.100 225.700 240.400 226.300 ;
        RECT 238.100 220.400 238.700 225.700 ;
        RECT 239.600 225.600 240.400 225.700 ;
        RECT 244.400 225.600 245.200 226.400 ;
        RECT 226.800 219.600 227.600 220.400 ;
        RECT 238.000 219.600 238.800 220.400 ;
        RECT 222.000 215.600 222.800 216.400 ;
        RECT 223.600 215.600 224.400 216.400 ;
        RECT 209.200 213.600 210.000 214.400 ;
        RECT 212.400 213.600 213.200 214.400 ;
        RECT 215.600 213.600 216.400 214.400 ;
        RECT 218.800 213.600 219.600 214.400 ;
        RECT 220.400 213.600 221.200 214.400 ;
        RECT 207.600 212.300 208.400 212.400 ;
        RECT 206.100 211.700 208.400 212.300 ;
        RECT 207.600 211.600 208.400 211.700 ;
        RECT 214.000 211.600 214.800 212.400 ;
        RECT 206.000 209.600 206.800 210.400 ;
        RECT 202.800 207.600 203.600 208.400 ;
        RECT 199.700 205.700 201.900 206.300 ;
        RECT 175.600 197.700 177.900 198.300 ;
        RECT 175.600 197.600 176.400 197.700 ;
        RECT 180.400 197.600 181.200 198.400 ;
        RECT 183.600 197.600 184.400 198.400 ;
        RECT 175.600 189.600 176.400 190.400 ;
        RECT 191.600 189.600 192.400 190.400 ;
        RECT 174.000 181.600 174.800 182.400 ;
        RECT 167.600 175.600 168.400 176.400 ;
        RECT 167.700 172.400 168.300 175.600 ;
        RECT 167.600 171.600 168.400 172.400 ;
        RECT 169.200 166.200 170.000 177.800 ;
        RECT 170.800 164.200 171.600 177.800 ;
        RECT 172.400 164.200 173.200 177.800 ;
        RECT 174.000 164.200 174.800 177.800 ;
        RECT 175.700 172.400 176.300 189.600 ;
        RECT 182.000 187.600 182.800 188.400 ;
        RECT 178.800 183.600 179.600 184.400 ;
        RECT 178.900 174.400 179.500 183.600 ;
        RECT 178.800 173.600 179.600 174.400 ;
        RECT 175.600 171.600 176.400 172.400 ;
        RECT 175.700 162.300 176.300 171.600 ;
        RECT 174.100 161.700 176.300 162.300 ;
        RECT 164.400 145.600 165.200 146.400 ;
        RECT 154.800 137.600 155.600 138.400 ;
        RECT 161.300 134.400 161.900 143.600 ;
        RECT 151.600 133.600 152.400 134.400 ;
        RECT 161.200 133.600 162.000 134.400 ;
        RECT 151.600 131.600 152.400 132.400 ;
        RECT 159.600 131.600 160.400 132.400 ;
        RECT 162.800 131.600 163.600 132.400 ;
        RECT 150.000 129.600 150.800 130.400 ;
        RECT 151.700 128.300 152.300 131.600 ;
        RECT 156.400 129.600 157.200 130.400 ;
        RECT 150.100 127.700 152.300 128.300 ;
        RECT 150.100 110.400 150.700 127.700 ;
        RECT 159.600 127.600 160.400 128.400 ;
        RECT 159.700 118.400 160.300 127.600 ;
        RECT 164.500 122.400 165.100 145.600 ;
        RECT 166.000 144.200 166.800 155.800 ;
        RECT 167.600 144.200 168.400 157.800 ;
        RECT 169.200 144.200 170.000 157.800 ;
        RECT 170.800 144.200 171.600 157.800 ;
        RECT 172.400 150.300 173.200 150.400 ;
        RECT 174.100 150.300 174.700 161.700 ;
        RECT 172.400 149.700 174.700 150.300 ;
        RECT 172.400 149.600 173.200 149.700 ;
        RECT 172.400 145.600 173.200 146.400 ;
        RECT 172.500 138.400 173.100 145.600 ;
        RECT 172.400 137.600 173.200 138.400 ;
        RECT 166.000 135.600 166.800 136.400 ;
        RECT 166.100 134.400 166.700 135.600 ;
        RECT 166.000 133.600 166.800 134.400 ;
        RECT 167.600 133.600 168.400 134.400 ;
        RECT 172.400 133.600 173.200 134.400 ;
        RECT 172.500 132.400 173.100 133.600 ;
        RECT 169.200 131.600 170.000 132.400 ;
        RECT 172.400 131.600 173.200 132.400 ;
        RECT 169.300 130.400 169.900 131.600 ;
        RECT 169.200 129.600 170.000 130.400 ;
        RECT 172.400 130.300 173.200 130.400 ;
        RECT 170.900 129.700 173.200 130.300 ;
        RECT 164.400 121.600 165.200 122.400 ;
        RECT 159.600 117.600 160.400 118.400 ;
        RECT 159.600 115.600 160.400 116.400 ;
        RECT 153.200 111.600 154.000 112.400 ;
        RECT 138.800 109.600 139.600 110.400 ;
        RECT 143.600 109.600 144.400 110.400 ;
        RECT 148.400 109.600 149.200 110.400 ;
        RECT 150.000 109.600 150.800 110.400 ;
        RECT 137.200 107.600 138.000 108.400 ;
        RECT 114.800 105.600 115.600 106.400 ;
        RECT 129.200 105.600 130.000 106.400 ;
        RECT 132.400 105.600 133.200 106.400 ;
        RECT 134.000 105.600 134.800 106.400 ;
        RECT 103.600 99.600 104.400 100.400 ;
        RECT 108.400 99.600 109.200 100.400 ;
        RECT 87.600 95.600 88.400 96.400 ;
        RECT 87.600 93.600 88.400 94.400 ;
        RECT 90.800 93.600 91.600 94.400 ;
        RECT 95.600 93.600 96.400 94.400 ;
        RECT 87.700 78.400 88.300 93.600 ;
        RECT 95.700 92.400 96.300 93.600 ;
        RECT 103.700 92.400 104.300 99.600 ;
        RECT 90.800 91.600 91.600 92.400 ;
        RECT 95.600 91.600 96.400 92.400 ;
        RECT 97.200 91.600 98.000 92.400 ;
        RECT 103.600 91.600 104.400 92.400 ;
        RECT 106.800 84.200 107.600 97.800 ;
        RECT 108.400 84.200 109.200 97.800 ;
        RECT 110.000 86.200 110.800 97.800 ;
        RECT 111.600 93.600 112.400 94.400 ;
        RECT 113.200 86.200 114.000 97.800 ;
        RECT 114.900 96.400 115.500 105.600 ;
        RECT 114.800 95.600 115.600 96.400 ;
        RECT 116.400 86.200 117.200 97.800 ;
        RECT 118.000 84.200 118.800 97.800 ;
        RECT 119.600 84.200 120.400 97.800 ;
        RECT 121.200 84.200 122.000 97.800 ;
        RECT 87.600 77.600 88.400 78.400 ;
        RECT 81.200 73.600 82.000 74.400 ;
        RECT 84.400 73.600 85.200 74.400 ;
        RECT 86.000 73.600 86.800 74.400 ;
        RECT 54.000 69.600 54.800 70.400 ;
        RECT 76.400 70.300 77.200 70.400 ;
        RECT 74.900 69.700 77.200 70.300 ;
        RECT 74.900 68.400 75.500 69.700 ;
        RECT 76.400 69.600 77.200 69.700 ;
        RECT 78.000 69.600 78.800 70.400 ;
        RECT 79.600 69.600 80.400 70.400 ;
        RECT 46.100 67.700 48.300 68.300 ;
        RECT 30.000 65.600 30.800 66.400 ;
        RECT 30.100 62.400 30.700 65.600 ;
        RECT 30.000 61.600 30.800 62.400 ;
        RECT 30.000 55.600 30.800 56.400 ;
        RECT 31.700 56.300 32.300 67.600 ;
        RECT 39.700 66.400 40.300 67.600 ;
        RECT 42.900 66.400 43.500 67.600 ;
        RECT 34.800 65.600 35.600 66.400 ;
        RECT 39.600 65.600 40.400 66.400 ;
        RECT 42.800 65.600 43.600 66.400 ;
        RECT 36.400 63.600 37.200 64.400 ;
        RECT 38.000 63.600 38.800 64.400 ;
        RECT 34.800 61.600 35.600 62.400 ;
        RECT 34.900 58.400 35.500 61.600 ;
        RECT 38.100 58.400 38.700 63.600 ;
        RECT 34.800 57.600 35.600 58.400 ;
        RECT 38.000 57.600 38.800 58.400 ;
        RECT 39.700 56.400 40.300 65.600 ;
        RECT 44.500 64.400 45.100 67.600 ;
        RECT 44.400 63.600 45.200 64.400 ;
        RECT 31.700 55.700 33.900 56.300 ;
        RECT 30.100 52.400 30.700 55.600 ;
        RECT 33.300 54.400 33.900 55.700 ;
        RECT 39.600 55.600 40.400 56.400 ;
        RECT 31.600 53.600 32.400 54.400 ;
        RECT 33.200 53.600 34.000 54.400 ;
        RECT 26.800 51.700 29.100 52.300 ;
        RECT 26.800 51.600 27.600 51.700 ;
        RECT 30.000 51.600 30.800 52.400 ;
        RECT 15.600 49.600 16.400 50.400 ;
        RECT 25.200 49.600 26.000 50.400 ;
        RECT 20.400 43.600 21.200 44.400 ;
        RECT 26.800 43.600 27.600 44.400 ;
        RECT 20.500 38.400 21.100 43.600 ;
        RECT 26.900 40.400 27.500 43.600 ;
        RECT 22.000 39.600 22.800 40.400 ;
        RECT 26.800 39.600 27.600 40.400 ;
        RECT 12.400 24.200 13.200 37.800 ;
        RECT 14.000 24.200 14.800 37.800 ;
        RECT 15.600 24.200 16.400 37.800 ;
        RECT 20.400 37.600 21.200 38.400 ;
        RECT 17.200 24.200 18.000 35.800 ;
        RECT 18.800 25.600 19.600 26.400 ;
        RECT 2.800 19.600 3.600 20.400 ;
        RECT 9.200 19.600 10.000 20.400 ;
        RECT 2.900 18.400 3.500 19.600 ;
        RECT 2.800 17.600 3.600 18.400 ;
        RECT 12.400 4.200 13.200 17.800 ;
        RECT 14.000 4.200 14.800 17.800 ;
        RECT 15.600 4.200 16.400 17.800 ;
        RECT 17.200 6.200 18.000 17.800 ;
        RECT 18.900 16.400 19.500 25.600 ;
        RECT 20.400 24.200 21.200 35.800 ;
        RECT 22.100 28.400 22.700 39.600 ;
        RECT 38.000 38.300 38.800 38.400 ;
        RECT 39.700 38.300 40.300 55.600 ;
        RECT 46.100 52.400 46.700 67.700 ;
        RECT 50.800 67.600 51.600 68.400 ;
        RECT 52.400 67.600 53.200 68.400 ;
        RECT 55.600 67.600 56.400 68.400 ;
        RECT 62.000 67.600 62.800 68.400 ;
        RECT 74.800 67.600 75.600 68.400 ;
        RECT 49.200 63.600 50.000 64.400 ;
        RECT 49.300 60.400 49.900 63.600 ;
        RECT 49.200 59.600 50.000 60.400 ;
        RECT 55.700 60.300 56.300 67.600 ;
        RECT 54.100 59.700 56.300 60.300 ;
        RECT 46.000 51.600 46.800 52.400 ;
        RECT 22.000 27.600 22.800 28.400 ;
        RECT 23.600 24.200 24.400 35.800 ;
        RECT 25.200 24.200 26.000 37.800 ;
        RECT 26.800 24.200 27.600 37.800 ;
        RECT 38.000 37.700 40.300 38.300 ;
        RECT 38.000 37.600 38.800 37.700 ;
        RECT 46.100 30.400 46.700 51.600 ;
        RECT 49.200 44.200 50.000 57.800 ;
        RECT 50.800 44.200 51.600 57.800 ;
        RECT 52.400 46.200 53.200 57.800 ;
        RECT 54.100 54.400 54.700 59.700 ;
        RECT 54.000 53.600 54.800 54.400 ;
        RECT 55.600 46.200 56.400 57.800 ;
        RECT 57.200 55.600 58.000 56.400 ;
        RECT 57.300 44.400 57.900 55.600 ;
        RECT 58.800 46.200 59.600 57.800 ;
        RECT 54.000 43.600 54.800 44.400 ;
        RECT 57.200 43.600 58.000 44.400 ;
        RECT 60.400 44.200 61.200 57.800 ;
        RECT 62.000 44.200 62.800 57.800 ;
        RECT 63.600 44.200 64.400 57.800 ;
        RECT 74.900 56.400 75.500 67.600 ;
        RECT 74.800 55.600 75.600 56.400 ;
        RECT 31.600 29.600 32.400 30.400 ;
        RECT 46.000 29.600 46.800 30.400 ;
        RECT 18.800 15.600 19.600 16.400 ;
        RECT 20.400 6.200 21.200 17.800 ;
        RECT 22.000 13.600 22.800 14.400 ;
        RECT 23.600 6.200 24.400 17.800 ;
        RECT 25.200 4.200 26.000 17.800 ;
        RECT 26.800 4.200 27.600 17.800 ;
        RECT 31.700 12.400 32.300 29.600 ;
        RECT 47.600 24.200 48.400 37.800 ;
        RECT 49.200 24.200 50.000 37.800 ;
        RECT 50.800 24.200 51.600 37.800 ;
        RECT 52.400 24.200 53.200 35.800 ;
        RECT 54.100 26.400 54.700 43.600 ;
        RECT 54.000 25.600 54.800 26.400 ;
        RECT 54.100 22.300 54.700 25.600 ;
        RECT 55.600 24.200 56.400 35.800 ;
        RECT 57.200 27.600 58.000 28.400 ;
        RECT 58.800 24.200 59.600 35.800 ;
        RECT 60.400 24.200 61.200 37.800 ;
        RECT 62.000 24.200 62.800 37.800 ;
        RECT 66.800 29.600 67.600 30.400 ;
        RECT 74.800 29.600 75.600 30.400 ;
        RECT 66.900 22.400 67.500 29.600 ;
        RECT 52.500 21.700 54.700 22.300 ;
        RECT 31.600 11.600 32.400 12.400 ;
        RECT 44.400 4.200 45.200 17.800 ;
        RECT 46.000 4.200 46.800 17.800 ;
        RECT 47.600 6.200 48.400 17.800 ;
        RECT 49.200 13.600 50.000 14.400 ;
        RECT 50.800 6.200 51.600 17.800 ;
        RECT 52.500 16.400 53.100 21.700 ;
        RECT 60.400 21.600 61.200 22.400 ;
        RECT 66.800 21.600 67.600 22.400 ;
        RECT 52.400 15.600 53.200 16.400 ;
        RECT 54.000 6.200 54.800 17.800 ;
        RECT 55.600 4.200 56.400 17.800 ;
        RECT 57.200 4.200 58.000 17.800 ;
        RECT 58.800 4.200 59.600 17.800 ;
        RECT 60.500 12.400 61.100 21.600 ;
        RECT 78.100 14.400 78.700 69.600 ;
        RECT 79.700 30.400 80.300 69.600 ;
        RECT 81.300 58.400 81.900 73.600 ;
        RECT 87.600 69.600 88.400 70.400 ;
        RECT 87.600 65.600 88.400 66.400 ;
        RECT 87.700 58.400 88.300 65.600 ;
        RECT 92.400 63.600 93.200 64.400 ;
        RECT 102.000 64.200 102.800 77.800 ;
        RECT 103.600 64.200 104.400 77.800 ;
        RECT 105.200 64.200 106.000 77.800 ;
        RECT 106.800 64.200 107.600 75.800 ;
        RECT 108.400 65.600 109.200 66.400 ;
        RECT 110.000 64.200 110.800 75.800 ;
        RECT 111.600 67.600 112.400 68.400 ;
        RECT 113.200 64.200 114.000 75.800 ;
        RECT 114.800 64.200 115.600 77.800 ;
        RECT 116.400 64.200 117.200 77.800 ;
        RECT 119.600 69.600 120.400 70.400 ;
        RECT 130.800 69.600 131.600 70.400 ;
        RECT 81.200 57.600 82.000 58.400 ;
        RECT 87.600 57.600 88.400 58.400 ;
        RECT 79.600 29.600 80.400 30.400 ;
        RECT 92.500 24.400 93.100 63.600 ;
        RECT 94.000 49.600 94.800 50.400 ;
        RECT 94.100 30.400 94.700 49.600 ;
        RECT 98.800 44.200 99.600 57.800 ;
        RECT 100.400 44.200 101.200 57.800 ;
        RECT 102.000 46.200 102.800 57.800 ;
        RECT 103.600 55.600 104.400 56.400 ;
        RECT 103.700 54.400 104.300 55.600 ;
        RECT 103.600 53.600 104.400 54.400 ;
        RECT 105.200 46.200 106.000 57.800 ;
        RECT 106.800 55.600 107.600 56.400 ;
        RECT 94.000 29.600 94.800 30.400 ;
        RECT 87.600 23.600 88.400 24.400 ;
        RECT 92.400 23.600 93.200 24.400 ;
        RECT 87.700 16.400 88.300 23.600 ;
        RECT 94.100 22.400 94.700 29.600 ;
        RECT 98.800 24.200 99.600 37.800 ;
        RECT 100.400 24.200 101.200 37.800 ;
        RECT 102.000 24.200 102.800 35.800 ;
        RECT 103.600 27.600 104.400 28.400 ;
        RECT 90.800 21.600 91.600 22.400 ;
        RECT 94.000 21.600 94.800 22.400 ;
        RECT 100.400 21.600 101.200 22.400 ;
        RECT 87.600 15.600 88.400 16.400 ;
        RECT 70.000 13.600 70.800 14.400 ;
        RECT 78.000 13.600 78.800 14.400 ;
        RECT 82.800 13.600 83.600 14.400 ;
        RECT 70.100 12.400 70.700 13.600 ;
        RECT 82.900 12.400 83.500 13.600 ;
        RECT 90.900 12.400 91.500 21.600 ;
        RECT 60.400 11.600 61.200 12.400 ;
        RECT 68.400 11.600 69.400 12.400 ;
        RECT 70.000 11.600 70.800 12.400 ;
        RECT 79.600 11.600 80.400 12.400 ;
        RECT 82.800 11.600 83.600 12.400 ;
        RECT 90.800 11.600 91.600 12.400 ;
        RECT 92.400 4.200 93.200 17.800 ;
        RECT 94.000 4.200 94.800 17.800 ;
        RECT 95.600 6.200 96.400 17.800 ;
        RECT 97.200 13.600 98.000 14.400 ;
        RECT 98.800 6.200 99.600 17.800 ;
        RECT 100.500 16.400 101.100 21.600 ;
        RECT 103.700 20.400 104.300 27.600 ;
        RECT 105.200 24.200 106.000 35.800 ;
        RECT 106.900 26.400 107.500 55.600 ;
        RECT 108.400 46.200 109.200 57.800 ;
        RECT 110.000 44.200 110.800 57.800 ;
        RECT 111.600 44.200 112.400 57.800 ;
        RECT 113.200 44.200 114.000 57.800 ;
        RECT 106.800 25.600 107.600 26.400 ;
        RECT 106.900 22.400 107.500 25.600 ;
        RECT 108.400 24.200 109.200 35.800 ;
        RECT 110.000 24.200 110.800 37.800 ;
        RECT 111.600 24.200 112.400 37.800 ;
        RECT 113.200 24.200 114.000 37.800 ;
        RECT 119.700 30.400 120.300 69.600 ;
        RECT 130.900 54.400 131.500 69.600 ;
        RECT 132.500 60.400 133.100 105.600 ;
        RECT 135.600 103.600 136.400 104.400 ;
        RECT 135.700 94.400 136.300 103.600 ;
        RECT 138.900 100.400 139.500 109.600 ;
        RECT 145.200 107.600 146.000 108.400 ;
        RECT 148.400 107.600 149.200 108.400 ;
        RECT 140.400 105.600 141.200 106.400 ;
        RECT 143.600 105.600 144.400 106.400 ;
        RECT 140.400 103.600 141.200 104.400 ;
        RECT 138.800 99.600 139.600 100.400 ;
        RECT 140.500 98.400 141.100 103.600 ;
        RECT 143.700 102.400 144.300 105.600 ;
        RECT 143.600 101.600 144.400 102.400 ;
        RECT 140.400 97.600 141.200 98.400 ;
        RECT 143.700 96.400 144.300 101.600 ;
        RECT 137.200 95.600 138.000 96.400 ;
        RECT 142.000 95.600 142.800 96.400 ;
        RECT 143.600 95.600 144.400 96.400 ;
        RECT 145.300 94.400 145.900 107.600 ;
        RECT 146.800 105.600 147.600 106.400 ;
        RECT 150.100 102.400 150.700 109.600 ;
        RECT 151.600 107.600 152.400 108.400 ;
        RECT 150.000 101.600 150.800 102.400 ;
        RECT 135.600 93.600 136.400 94.400 ;
        RECT 145.200 93.600 146.000 94.400 ;
        RECT 145.300 80.400 145.900 93.600 ;
        RECT 150.000 91.600 150.800 92.400 ;
        RECT 150.000 90.300 150.800 90.400 ;
        RECT 151.700 90.300 152.300 107.600 ;
        RECT 153.300 98.400 153.900 111.600 ;
        RECT 154.800 109.600 155.600 110.400 ;
        RECT 154.800 107.600 155.600 108.400 ;
        RECT 159.700 106.400 160.300 115.600 ;
        RECT 164.400 113.600 165.200 114.400 ;
        RECT 164.500 110.400 165.100 113.600 ;
        RECT 170.900 112.400 171.500 129.700 ;
        RECT 172.400 129.600 173.200 129.700 ;
        RECT 167.600 111.600 168.400 112.400 ;
        RECT 170.800 111.600 171.600 112.400 ;
        RECT 164.400 109.600 165.200 110.400 ;
        RECT 167.600 109.600 168.400 110.400 ;
        RECT 170.800 109.600 171.600 110.400 ;
        RECT 174.100 108.400 174.700 149.700 ;
        RECT 175.600 149.600 176.400 150.400 ;
        RECT 175.700 138.400 176.300 149.600 ;
        RECT 175.600 137.600 176.400 138.400 ;
        RECT 178.900 130.400 179.500 173.600 ;
        RECT 180.400 143.600 181.200 144.400 ;
        RECT 182.100 142.300 182.700 187.600 ;
        RECT 193.200 184.200 194.000 197.800 ;
        RECT 194.800 184.200 195.600 197.800 ;
        RECT 196.400 184.200 197.200 197.800 ;
        RECT 198.000 184.200 198.800 195.800 ;
        RECT 199.700 186.400 200.300 205.700 ;
        RECT 214.100 204.400 214.700 211.600 ;
        RECT 215.700 210.400 216.300 213.600 ;
        RECT 215.600 209.600 216.400 210.400 ;
        RECT 217.200 209.600 218.000 210.400 ;
        RECT 201.200 203.600 202.000 204.400 ;
        RECT 214.000 203.600 214.800 204.400 ;
        RECT 201.300 198.300 201.900 203.600 ;
        RECT 201.300 197.700 203.500 198.300 ;
        RECT 199.600 185.600 200.400 186.400 ;
        RECT 201.200 184.200 202.000 195.800 ;
        RECT 202.900 188.400 203.500 197.700 ;
        RECT 202.800 187.600 203.600 188.400 ;
        RECT 204.400 184.200 205.200 195.800 ;
        RECT 206.000 184.200 206.800 197.800 ;
        RECT 207.600 184.200 208.400 197.800 ;
        RECT 218.900 194.400 219.500 213.600 ;
        RECT 222.000 211.600 222.800 212.400 ;
        RECT 223.700 198.400 224.300 215.600 ;
        RECT 226.900 214.400 227.500 219.600 ;
        RECT 233.200 215.600 234.000 216.400 ;
        RECT 226.800 213.600 227.600 214.400 ;
        RECT 233.300 212.400 233.900 215.600 ;
        RECT 226.800 211.600 227.600 212.400 ;
        RECT 228.400 211.600 229.200 212.400 ;
        RECT 233.200 211.600 234.000 212.400 ;
        RECT 225.200 209.600 226.000 210.400 ;
        RECT 223.600 197.600 224.400 198.400 ;
        RECT 218.800 193.600 219.600 194.400 ;
        RECT 222.000 193.600 222.800 194.400 ;
        RECT 210.800 189.600 211.600 190.400 ;
        RECT 218.800 189.600 219.600 190.400 ;
        RECT 193.200 175.600 194.000 176.400 ;
        RECT 199.600 175.600 200.400 176.400 ;
        RECT 186.800 173.600 187.600 174.400 ;
        RECT 210.900 172.400 211.500 189.600 ;
        RECT 218.800 187.600 219.600 188.400 ;
        RECT 218.900 186.400 219.500 187.600 ;
        RECT 222.100 186.400 222.700 193.600 ;
        RECT 223.600 189.600 224.400 190.400 ;
        RECT 218.800 185.600 219.600 186.400 ;
        RECT 222.000 185.600 222.800 186.400 ;
        RECT 223.700 184.400 224.300 189.600 ;
        RECT 223.600 183.600 224.400 184.400 ;
        RECT 226.900 182.400 227.500 211.600 ;
        RECT 228.500 208.400 229.100 211.600 ;
        RECT 231.600 209.600 232.400 210.400 ;
        RECT 228.400 207.600 229.200 208.400 ;
        RECT 228.400 205.600 229.200 206.400 ;
        RECT 228.500 194.400 229.100 205.600 ;
        RECT 228.400 193.600 229.200 194.400 ;
        RECT 231.700 192.400 232.300 209.600 ;
        RECT 233.200 207.600 234.000 208.400 ;
        RECT 233.300 192.400 233.900 207.600 ;
        RECT 228.400 191.600 229.200 192.400 ;
        RECT 231.600 191.600 232.400 192.400 ;
        RECT 233.200 191.600 234.000 192.400 ;
        RECT 228.500 186.400 229.100 191.600 ;
        RECT 230.000 187.600 230.800 188.400 ;
        RECT 233.300 188.300 233.900 191.600 ;
        RECT 234.800 189.600 235.600 190.400 ;
        RECT 238.100 188.400 238.700 219.600 ;
        RECT 244.500 214.400 245.100 225.600 ;
        RECT 244.400 213.600 245.200 214.400 ;
        RECT 239.600 212.300 240.400 212.400 ;
        RECT 239.600 211.700 241.900 212.300 ;
        RECT 239.600 211.600 240.400 211.700 ;
        RECT 241.300 210.400 241.900 211.700 ;
        RECT 246.000 211.600 246.800 212.400 ;
        RECT 239.600 209.600 240.400 210.400 ;
        RECT 241.200 209.600 242.000 210.400 ;
        RECT 239.700 208.400 240.300 209.600 ;
        RECT 239.600 207.600 240.400 208.400 ;
        RECT 242.800 207.600 243.600 208.400 ;
        RECT 233.300 187.700 235.500 188.300 ;
        RECT 228.400 185.600 229.200 186.400 ;
        RECT 230.000 185.600 230.800 186.400 ;
        RECT 226.800 181.600 227.600 182.400 ;
        RECT 196.400 171.600 197.200 172.400 ;
        RECT 210.800 171.600 211.600 172.400 ;
        RECT 196.500 170.400 197.100 171.600 ;
        RECT 190.000 169.600 190.800 170.400 ;
        RECT 196.400 169.600 197.200 170.400 ;
        RECT 199.600 169.600 200.400 170.400 ;
        RECT 183.600 163.600 184.400 164.400 ;
        RECT 183.700 152.400 184.300 163.600 ;
        RECT 190.100 154.400 190.700 169.600 ;
        RECT 190.000 153.600 190.800 154.400 ;
        RECT 183.600 151.600 184.400 152.400 ;
        RECT 188.400 151.600 189.200 152.400 ;
        RECT 193.200 151.600 194.000 152.400 ;
        RECT 180.500 141.700 182.700 142.300 ;
        RECT 178.800 129.600 179.600 130.400 ;
        RECT 180.500 116.400 181.100 141.700 ;
        RECT 183.700 140.300 184.300 151.600 ;
        RECT 193.300 150.400 193.900 151.600 ;
        RECT 199.700 150.400 200.300 169.600 ;
        RECT 202.800 163.600 203.600 164.400 ;
        RECT 212.400 164.200 213.200 177.800 ;
        RECT 214.000 164.200 214.800 177.800 ;
        RECT 215.600 164.200 216.400 177.800 ;
        RECT 217.200 166.200 218.000 177.800 ;
        RECT 218.800 175.600 219.600 176.400 ;
        RECT 218.900 172.400 219.500 175.600 ;
        RECT 218.800 171.600 219.600 172.400 ;
        RECT 220.400 166.200 221.200 177.800 ;
        RECT 222.000 173.600 222.800 174.400 ;
        RECT 222.000 171.600 222.800 172.400 ;
        RECT 218.800 163.600 219.600 164.400 ;
        RECT 201.200 151.600 202.000 152.400 ;
        RECT 185.200 149.600 186.000 150.400 ;
        RECT 193.200 149.600 194.000 150.400 ;
        RECT 199.600 149.600 200.400 150.400 ;
        RECT 182.100 139.700 184.300 140.300 ;
        RECT 182.100 136.400 182.700 139.700 ;
        RECT 182.000 135.600 182.800 136.400 ;
        RECT 183.400 132.300 184.400 132.400 ;
        RECT 185.300 132.300 185.900 149.600 ;
        RECT 193.200 147.600 194.000 148.400 ;
        RECT 201.300 146.400 201.900 151.600 ;
        RECT 202.900 146.400 203.500 163.600 ;
        RECT 218.900 150.400 219.500 163.600 ;
        RECT 220.400 161.600 221.200 162.400 ;
        RECT 220.500 152.400 221.100 161.600 ;
        RECT 220.400 151.600 221.200 152.400 ;
        RECT 204.400 149.600 205.200 150.400 ;
        RECT 207.600 149.600 208.400 150.400 ;
        RECT 210.800 149.600 211.600 150.400 ;
        RECT 218.800 149.600 219.600 150.400 ;
        RECT 207.700 148.400 208.300 149.600 ;
        RECT 206.000 147.600 206.800 148.400 ;
        RECT 207.600 147.600 208.400 148.400 ;
        RECT 210.900 146.400 211.500 149.600 ;
        RECT 215.600 147.600 216.400 148.400 ;
        RECT 194.800 145.600 195.600 146.400 ;
        RECT 201.200 145.600 202.000 146.400 ;
        RECT 202.800 145.600 203.600 146.400 ;
        RECT 207.600 145.600 208.400 146.400 ;
        RECT 210.800 145.600 211.600 146.400 ;
        RECT 183.400 131.700 185.900 132.300 ;
        RECT 183.400 131.600 184.400 131.700 ;
        RECT 185.200 127.600 186.000 128.400 ;
        RECT 180.400 115.600 181.200 116.400 ;
        RECT 178.800 113.600 179.600 114.400 ;
        RECT 178.900 112.400 179.500 113.600 ;
        RECT 178.800 111.600 179.600 112.400 ;
        RECT 183.600 109.600 184.400 110.400 ;
        RECT 183.700 108.400 184.300 109.600 ;
        RECT 174.000 107.600 174.800 108.400 ;
        RECT 175.600 107.600 176.400 108.400 ;
        RECT 183.600 107.600 184.400 108.400 ;
        RECT 159.600 105.600 160.400 106.400 ;
        RECT 161.200 105.600 162.000 106.400 ;
        RECT 174.000 105.600 174.800 106.400 ;
        RECT 161.300 104.400 161.900 105.600 ;
        RECT 175.700 104.400 176.300 107.600 ;
        RECT 177.200 105.600 178.000 106.400 ;
        RECT 161.200 103.600 162.000 104.400 ;
        RECT 175.600 103.600 176.400 104.400 ;
        RECT 183.700 98.400 184.300 107.600 ;
        RECT 153.200 97.600 154.000 98.400 ;
        RECT 154.800 93.600 155.600 94.400 ;
        RECT 153.200 91.600 154.000 92.400 ;
        RECT 150.000 89.700 152.300 90.300 ;
        RECT 150.000 89.600 150.800 89.700 ;
        RECT 153.200 89.600 154.000 90.400 ;
        RECT 154.900 88.400 155.500 93.600 ;
        RECT 156.400 90.200 157.200 95.800 ;
        RECT 154.800 87.600 155.600 88.400 ;
        RECT 159.600 86.200 160.400 97.800 ;
        RECT 164.400 93.600 165.200 94.400 ;
        RECT 161.200 91.800 162.000 92.600 ;
        RECT 161.300 90.400 161.900 91.800 ;
        RECT 161.200 89.600 162.000 90.400 ;
        RECT 134.000 79.600 134.800 80.400 ;
        RECT 145.200 79.600 146.000 80.400 ;
        RECT 134.100 78.400 134.700 79.600 ;
        RECT 134.000 77.600 134.800 78.400 ;
        RECT 134.000 67.600 134.800 68.400 ;
        RECT 132.400 59.600 133.200 60.400 ;
        RECT 132.500 56.400 133.100 59.600 ;
        RECT 134.100 58.400 134.700 67.600 ;
        RECT 143.600 64.200 144.400 77.800 ;
        RECT 145.200 64.200 146.000 77.800 ;
        RECT 146.800 64.200 147.600 77.800 ;
        RECT 148.400 64.200 149.200 75.800 ;
        RECT 150.000 65.600 150.800 66.400 ;
        RECT 151.600 64.200 152.400 75.800 ;
        RECT 153.200 67.600 154.000 68.400 ;
        RECT 154.800 64.200 155.600 75.800 ;
        RECT 156.400 64.200 157.200 77.800 ;
        RECT 158.000 64.200 158.800 77.800 ;
        RECT 162.800 71.600 163.600 72.400 ;
        RECT 159.600 67.600 160.400 68.400 ;
        RECT 148.400 61.600 149.200 62.400 ;
        RECT 134.000 57.600 134.800 58.400 ;
        RECT 138.800 57.600 139.600 58.400 ;
        RECT 138.900 56.400 139.500 57.600 ;
        RECT 132.400 55.600 133.200 56.400 ;
        RECT 135.600 55.600 136.400 56.400 ;
        RECT 137.200 55.600 138.000 56.400 ;
        RECT 138.800 55.600 139.600 56.400 ;
        RECT 143.600 56.300 144.400 56.400 ;
        RECT 143.600 55.700 147.500 56.300 ;
        RECT 143.600 55.600 144.400 55.700 ;
        RECT 130.800 53.600 131.600 54.400 ;
        RECT 122.800 51.600 123.800 52.400 ;
        RECT 114.800 29.600 115.600 30.400 ;
        RECT 119.600 29.600 120.400 30.400 ;
        RECT 119.600 23.600 120.400 24.400 ;
        RECT 122.800 23.600 123.600 24.400 ;
        RECT 106.800 21.600 107.600 22.400 ;
        RECT 103.600 19.600 104.400 20.400 ;
        RECT 100.400 15.600 101.200 16.400 ;
        RECT 102.000 6.200 102.800 17.800 ;
        RECT 103.600 4.200 104.400 17.800 ;
        RECT 105.200 4.200 106.000 17.800 ;
        RECT 106.800 4.200 107.600 17.800 ;
        RECT 119.700 16.400 120.300 23.600 ;
        RECT 121.200 19.600 122.000 20.400 ;
        RECT 121.300 18.400 121.900 19.600 ;
        RECT 121.200 17.600 122.000 18.400 ;
        RECT 119.600 15.600 120.400 16.400 ;
        RECT 116.400 11.600 117.400 12.400 ;
        RECT 130.900 10.400 131.500 53.600 ;
        RECT 135.600 52.300 136.400 52.400 ;
        RECT 137.300 52.300 137.900 55.600 ;
        RECT 135.600 51.700 137.900 52.300 ;
        RECT 135.600 51.600 136.400 51.700 ;
        RECT 145.200 51.600 146.000 52.400 ;
        RECT 146.900 52.300 147.500 55.700 ;
        RECT 148.500 54.400 149.100 61.600 ;
        RECT 159.700 58.400 160.300 67.600 ;
        RECT 164.500 66.400 165.100 93.600 ;
        RECT 169.200 86.200 170.000 97.800 ;
        RECT 174.000 97.600 174.800 98.400 ;
        RECT 183.600 97.600 184.400 98.400 ;
        RECT 185.300 96.400 185.900 127.600 ;
        RECT 193.200 124.200 194.000 137.800 ;
        RECT 194.800 124.200 195.600 137.800 ;
        RECT 196.400 124.200 197.200 137.800 ;
        RECT 198.000 126.200 198.800 137.800 ;
        RECT 199.600 135.600 200.400 136.400 ;
        RECT 199.700 122.400 200.300 135.600 ;
        RECT 201.200 126.200 202.000 137.800 ;
        RECT 202.800 133.600 203.600 134.400 ;
        RECT 204.400 126.200 205.200 137.800 ;
        RECT 206.000 124.200 206.800 137.800 ;
        RECT 207.600 124.200 208.400 137.800 ;
        RECT 217.200 135.600 218.000 136.400 ;
        RECT 217.300 132.400 217.900 135.600 ;
        RECT 218.800 133.600 219.600 134.400 ;
        RECT 210.800 131.600 211.600 132.400 ;
        RECT 217.200 131.600 218.000 132.400 ;
        RECT 196.400 121.600 197.200 122.400 ;
        RECT 199.600 121.600 200.400 122.400 ;
        RECT 188.400 104.200 189.200 117.800 ;
        RECT 190.000 104.200 190.800 117.800 ;
        RECT 191.600 104.200 192.400 115.800 ;
        RECT 193.200 107.600 194.000 108.400 ;
        RECT 194.800 104.200 195.600 115.800 ;
        RECT 196.500 106.400 197.100 121.600 ;
        RECT 196.400 105.600 197.200 106.400 ;
        RECT 196.500 102.300 197.100 105.600 ;
        RECT 198.000 104.200 198.800 115.800 ;
        RECT 199.600 104.200 200.400 117.800 ;
        RECT 201.200 104.200 202.000 117.800 ;
        RECT 202.800 104.200 203.600 117.800 ;
        RECT 207.600 105.600 208.400 106.400 ;
        RECT 196.500 101.700 198.700 102.300 ;
        RECT 188.400 99.600 189.200 100.400 ;
        RECT 185.200 95.600 186.000 96.400 ;
        RECT 185.300 86.400 185.900 95.600 ;
        RECT 188.500 92.400 189.100 99.600 ;
        RECT 193.200 96.300 194.000 96.400 ;
        RECT 196.400 96.300 197.200 96.400 ;
        RECT 193.200 95.700 197.200 96.300 ;
        RECT 193.200 95.600 194.000 95.700 ;
        RECT 196.400 95.600 197.200 95.700 ;
        RECT 193.200 93.600 194.000 94.400 ;
        RECT 188.400 91.600 189.200 92.400 ;
        RECT 185.200 85.600 186.000 86.400 ;
        RECT 178.800 83.600 179.600 84.400 ;
        RECT 193.200 83.600 194.000 84.400 ;
        RECT 167.600 73.600 168.400 74.400 ;
        RECT 167.700 72.400 168.300 73.600 ;
        RECT 167.600 71.600 168.400 72.400 ;
        RECT 177.200 71.600 178.000 72.400 ;
        RECT 177.300 70.400 177.900 71.600 ;
        RECT 177.200 69.600 178.000 70.400 ;
        RECT 164.400 65.600 165.200 66.400 ;
        RECT 159.600 57.600 160.400 58.400 ;
        RECT 169.200 57.600 170.000 58.400 ;
        RECT 170.800 57.600 171.600 58.400 ;
        RECT 170.900 56.400 171.500 57.600 ;
        RECT 154.800 55.600 155.600 56.400 ;
        RECT 159.600 55.600 160.400 56.400 ;
        RECT 166.000 55.600 166.800 56.400 ;
        RECT 170.800 55.600 171.600 56.400 ;
        RECT 148.400 53.600 149.200 54.400 ;
        RECT 154.900 52.400 155.500 55.600 ;
        RECT 148.400 52.300 149.200 52.400 ;
        RECT 146.900 51.700 149.200 52.300 ;
        RECT 148.400 51.600 149.200 51.700 ;
        RECT 154.800 51.600 155.600 52.400 ;
        RECT 158.000 51.600 158.800 52.400 ;
        RECT 145.300 50.400 145.900 51.600 ;
        RECT 159.700 50.400 160.300 55.600 ;
        RECT 162.800 53.600 163.600 54.400 ;
        RECT 166.100 52.400 166.700 55.600 ;
        RECT 174.000 53.600 174.800 54.400 ;
        RECT 162.800 51.600 163.600 52.400 ;
        RECT 166.000 51.600 166.800 52.400 ;
        RECT 134.000 49.600 134.800 50.400 ;
        RECT 145.200 49.600 146.000 50.400 ;
        RECT 159.600 49.600 160.400 50.400 ;
        RECT 134.100 38.400 134.700 49.600 ;
        RECT 142.000 43.600 142.800 44.400 ;
        RECT 134.000 37.600 134.800 38.400 ;
        RECT 135.600 33.600 136.400 34.400 ;
        RECT 135.700 24.400 136.300 33.600 ;
        RECT 135.600 23.600 136.400 24.400 ;
        RECT 135.700 14.400 136.300 23.600 ;
        RECT 142.100 14.400 142.700 43.600 ;
        RECT 166.100 42.400 166.700 51.600 ;
        RECT 177.300 50.400 177.900 69.600 ;
        RECT 177.200 49.600 178.000 50.400 ;
        RECT 166.000 41.600 166.800 42.400 ;
        RECT 169.200 41.600 170.000 42.400 ;
        RECT 162.800 39.600 163.600 40.400 ;
        RECT 166.000 39.600 166.800 40.400 ;
        RECT 143.600 24.200 144.400 37.800 ;
        RECT 145.200 24.200 146.000 37.800 ;
        RECT 146.800 24.200 147.600 37.800 ;
        RECT 148.400 24.200 149.200 35.800 ;
        RECT 150.000 25.600 150.800 26.400 ;
        RECT 150.100 22.400 150.700 25.600 ;
        RECT 151.600 24.200 152.400 35.800 ;
        RECT 153.200 27.600 154.000 28.400 ;
        RECT 153.300 24.400 153.900 27.600 ;
        RECT 153.200 23.600 154.000 24.400 ;
        RECT 154.800 24.200 155.600 35.800 ;
        RECT 156.400 24.200 157.200 37.800 ;
        RECT 158.000 24.200 158.800 37.800 ;
        RECT 162.900 32.400 163.500 39.600 ;
        RECT 162.800 31.600 163.600 32.400 ;
        RECT 162.900 30.400 163.500 31.600 ;
        RECT 162.800 29.600 163.600 30.400 ;
        RECT 150.000 21.600 150.800 22.400 ;
        RECT 154.800 21.600 155.600 22.400 ;
        RECT 135.600 13.600 136.400 14.400 ;
        RECT 142.000 13.600 142.800 14.400 ;
        RECT 130.800 9.600 131.600 10.400 ;
        RECT 148.400 4.200 149.200 17.800 ;
        RECT 150.000 4.200 150.800 17.800 ;
        RECT 151.600 4.200 152.400 17.800 ;
        RECT 153.200 6.200 154.000 17.800 ;
        RECT 154.900 16.400 155.500 21.600 ;
        RECT 154.800 15.600 155.600 16.400 ;
        RECT 156.400 6.200 157.200 17.800 ;
        RECT 158.000 13.600 158.800 14.400 ;
        RECT 159.600 6.200 160.400 17.800 ;
        RECT 161.200 4.200 162.000 17.800 ;
        RECT 162.800 4.200 163.600 17.800 ;
        RECT 166.100 12.400 166.700 39.600 ;
        RECT 169.300 38.400 169.900 41.600 ;
        RECT 178.900 40.400 179.500 83.600 ;
        RECT 193.300 80.400 193.900 83.600 ;
        RECT 185.200 79.600 186.000 80.400 ;
        RECT 193.200 79.600 194.000 80.400 ;
        RECT 180.400 64.200 181.200 77.800 ;
        RECT 182.000 64.200 182.800 77.800 ;
        RECT 183.600 64.200 184.400 75.800 ;
        RECT 185.300 68.400 185.900 79.600 ;
        RECT 185.200 67.600 186.000 68.400 ;
        RECT 186.800 64.200 187.600 75.800 ;
        RECT 188.400 65.600 189.200 66.400 ;
        RECT 190.000 64.200 190.800 75.800 ;
        RECT 191.600 64.200 192.400 77.800 ;
        RECT 193.200 64.200 194.000 77.800 ;
        RECT 194.800 64.200 195.600 77.800 ;
        RECT 196.400 69.600 197.200 70.400 ;
        RECT 198.100 66.400 198.700 101.700 ;
        RECT 207.700 96.400 208.300 105.600 ;
        RECT 209.200 97.600 210.000 98.400 ;
        RECT 207.600 95.600 208.400 96.400 ;
        RECT 204.400 93.600 205.200 94.400 ;
        RECT 204.500 90.400 205.100 93.600 ;
        RECT 207.700 92.400 208.300 95.600 ;
        RECT 209.300 94.400 209.900 97.600 ;
        RECT 209.200 93.600 210.000 94.400 ;
        RECT 207.600 91.600 208.400 92.400 ;
        RECT 199.600 89.600 200.400 90.400 ;
        RECT 204.400 89.600 205.200 90.400 ;
        RECT 204.500 88.400 205.100 89.600 ;
        RECT 204.400 87.600 205.200 88.400 ;
        RECT 204.500 78.400 205.100 87.600 ;
        RECT 209.300 78.400 209.900 93.600 ;
        RECT 204.400 77.600 205.200 78.400 ;
        RECT 209.200 77.600 210.000 78.400 ;
        RECT 210.900 70.400 211.500 131.600 ;
        RECT 220.500 130.400 221.100 151.600 ;
        RECT 222.100 150.400 222.700 171.600 ;
        RECT 223.600 166.200 224.400 177.800 ;
        RECT 225.200 164.200 226.000 177.800 ;
        RECT 226.800 164.200 227.600 177.800 ;
        RECT 230.100 168.400 230.700 185.600 ;
        RECT 233.200 183.600 234.000 184.400 ;
        RECT 233.300 180.400 233.900 183.600 ;
        RECT 233.200 179.600 234.000 180.400 ;
        RECT 230.000 167.600 230.800 168.400 ;
        RECT 234.900 166.400 235.500 187.700 ;
        RECT 238.000 187.600 238.800 188.400 ;
        RECT 238.100 186.400 238.700 187.600 ;
        RECT 238.000 185.600 238.800 186.400 ;
        RECT 239.600 183.600 240.400 184.400 ;
        RECT 236.400 175.600 237.200 176.400 ;
        RECT 234.800 165.600 235.600 166.400 ;
        RECT 236.500 164.400 237.100 175.600 ;
        RECT 238.000 173.600 238.800 174.400 ;
        RECT 238.000 171.600 238.800 172.400 ;
        RECT 238.100 164.400 238.700 171.600 ;
        RECT 236.400 163.600 237.200 164.400 ;
        RECT 238.000 163.600 238.800 164.400 ;
        RECT 222.000 149.600 222.800 150.400 ;
        RECT 225.200 149.600 226.000 150.400 ;
        RECT 230.000 144.200 230.800 157.800 ;
        RECT 231.600 144.200 232.400 157.800 ;
        RECT 233.200 144.200 234.000 155.800 ;
        RECT 234.800 147.600 235.600 148.400 ;
        RECT 236.400 144.200 237.200 155.800 ;
        RECT 238.100 146.400 238.700 163.600 ;
        RECT 239.700 158.400 240.300 183.600 ;
        RECT 241.200 171.600 242.000 172.400 ;
        RECT 242.900 162.400 243.500 207.600 ;
        RECT 246.100 190.300 246.700 211.600 ;
        RECT 247.700 206.400 248.300 243.600 ;
        RECT 249.300 234.400 249.900 265.600 ;
        RECT 255.700 264.400 256.300 269.600 ;
        RECT 258.900 266.400 259.500 269.600 ;
        RECT 260.400 267.600 261.200 268.400 ;
        RECT 269.800 267.600 270.800 268.400 ;
        RECT 260.500 266.400 261.100 267.600 ;
        RECT 258.800 265.600 259.600 266.400 ;
        RECT 260.400 265.600 261.200 266.400 ;
        RECT 252.400 263.600 253.200 264.400 ;
        RECT 255.600 263.600 256.400 264.400 ;
        RECT 279.600 264.200 280.400 277.800 ;
        RECT 281.200 264.200 282.000 277.800 ;
        RECT 282.800 264.200 283.600 277.800 ;
        RECT 284.400 264.200 285.200 275.800 ;
        RECT 286.000 265.600 286.800 266.400 ;
        RECT 252.500 260.400 253.100 263.600 ;
        RECT 286.100 260.400 286.700 265.600 ;
        RECT 287.600 264.200 288.400 275.800 ;
        RECT 289.200 267.600 290.000 268.400 ;
        RECT 289.200 265.600 290.000 266.400 ;
        RECT 252.400 259.600 253.200 260.400 ;
        RECT 286.000 259.600 286.800 260.400 ;
        RECT 257.200 244.200 258.000 257.800 ;
        RECT 258.800 244.200 259.600 257.800 ;
        RECT 260.400 244.200 261.200 257.800 ;
        RECT 262.000 246.200 262.800 257.800 ;
        RECT 263.600 255.600 264.400 256.400 ;
        RECT 263.700 242.400 264.300 255.600 ;
        RECT 265.200 246.200 266.000 257.800 ;
        RECT 266.800 253.600 267.600 254.400 ;
        RECT 266.900 242.400 267.500 253.600 ;
        RECT 268.400 246.200 269.200 257.800 ;
        RECT 270.000 244.200 270.800 257.800 ;
        RECT 271.600 244.200 272.400 257.800 ;
        RECT 286.100 256.400 286.700 259.600 ;
        RECT 289.300 258.400 289.900 265.600 ;
        RECT 290.800 264.200 291.600 275.800 ;
        RECT 292.400 264.200 293.200 277.800 ;
        RECT 294.000 264.200 294.800 277.800 ;
        RECT 295.700 272.000 296.300 279.600 ;
        RECT 295.600 271.200 296.400 272.000 ;
        RECT 305.300 262.400 305.900 291.600 ;
        RECT 306.800 279.600 307.600 280.400 ;
        RECT 306.900 272.400 307.500 279.600 ;
        RECT 306.800 271.600 307.600 272.400 ;
        RECT 308.500 266.400 309.100 305.600 ;
        RECT 310.000 304.200 310.800 315.800 ;
        RECT 311.600 307.600 312.400 308.400 ;
        RECT 311.700 294.400 312.300 307.600 ;
        RECT 313.200 304.200 314.000 315.800 ;
        RECT 314.800 304.200 315.600 317.800 ;
        RECT 316.400 304.200 317.200 317.800 ;
        RECT 318.100 312.000 318.700 321.600 ;
        RECT 322.900 312.400 323.500 333.600 ;
        RECT 324.400 326.200 325.200 337.800 ;
        RECT 326.000 337.600 326.800 338.400 ;
        RECT 326.100 336.400 326.700 337.600 ;
        RECT 326.000 335.600 326.800 336.400 ;
        RECT 327.600 326.200 328.400 337.800 ;
        RECT 329.200 324.200 330.000 337.800 ;
        RECT 330.800 324.200 331.600 337.800 ;
        RECT 332.400 324.200 333.200 337.800 ;
        RECT 332.400 319.600 333.200 320.400 ;
        RECT 330.800 317.600 331.600 318.400 ;
        RECT 332.500 314.400 333.100 319.600 ;
        RECT 326.000 313.600 326.800 314.400 ;
        RECT 332.400 313.600 333.200 314.400 ;
        RECT 318.000 311.200 318.800 312.000 ;
        RECT 322.800 311.600 323.600 312.400 ;
        RECT 318.100 302.400 318.700 311.200 ;
        RECT 326.100 310.400 326.700 313.600 ;
        RECT 326.000 309.600 326.800 310.400 ;
        RECT 327.600 307.600 328.400 308.400 ;
        RECT 330.800 307.600 331.600 308.400 ;
        RECT 318.000 301.600 318.800 302.400 ;
        RECT 327.700 298.400 328.300 307.600 ;
        RECT 330.900 306.400 331.500 307.600 ;
        RECT 330.800 305.600 331.600 306.400 ;
        RECT 327.600 297.600 328.400 298.400 ;
        RECT 330.800 297.600 331.600 298.400 ;
        RECT 330.900 296.400 331.500 297.600 ;
        RECT 330.800 295.600 331.600 296.400 ;
        RECT 311.600 293.600 312.400 294.400 ;
        RECT 310.000 291.600 310.800 292.400 ;
        RECT 327.600 291.600 328.400 292.400 ;
        RECT 308.400 265.600 309.200 266.400 ;
        RECT 305.200 261.600 306.000 262.400 ;
        RECT 310.100 260.400 310.700 291.600 ;
        RECT 329.200 289.600 330.000 290.400 ;
        RECT 329.300 288.400 329.900 289.600 ;
        RECT 329.200 287.600 330.000 288.400 ;
        RECT 330.800 287.600 331.600 288.400 ;
        RECT 311.600 264.200 312.400 277.800 ;
        RECT 313.200 264.200 314.000 277.800 ;
        RECT 314.800 264.200 315.600 275.800 ;
        RECT 316.400 267.600 317.200 268.400 ;
        RECT 316.500 260.400 317.100 267.600 ;
        RECT 318.000 264.200 318.800 275.800 ;
        RECT 319.600 265.600 320.400 266.400 ;
        RECT 321.200 264.200 322.000 275.800 ;
        RECT 322.800 264.200 323.600 277.800 ;
        RECT 324.400 264.200 325.200 277.800 ;
        RECT 326.000 264.200 326.800 277.800 ;
        RECT 318.000 261.600 318.800 262.400 ;
        RECT 327.600 261.600 328.400 262.400 ;
        RECT 305.200 259.600 306.000 260.400 ;
        RECT 310.000 259.600 310.800 260.400 ;
        RECT 316.400 259.600 317.200 260.400 ;
        RECT 289.200 257.600 290.000 258.400 ;
        RECT 286.000 255.600 286.800 256.400 ;
        RECT 276.400 249.600 277.200 250.400 ;
        RECT 257.200 241.600 258.000 242.400 ;
        RECT 263.600 241.600 264.400 242.400 ;
        RECT 266.800 241.600 267.600 242.400 ;
        RECT 249.200 233.600 250.000 234.400 ;
        RECT 249.200 229.600 250.000 230.400 ;
        RECT 250.800 224.200 251.600 237.800 ;
        RECT 252.400 224.200 253.200 237.800 ;
        RECT 254.000 224.200 254.800 237.800 ;
        RECT 255.600 224.200 256.400 235.800 ;
        RECT 257.300 226.400 257.900 241.600 ;
        RECT 257.200 225.600 258.000 226.400 ;
        RECT 257.300 220.400 257.900 225.600 ;
        RECT 258.800 224.200 259.600 235.800 ;
        RECT 260.400 227.600 261.200 228.400 ;
        RECT 262.000 224.200 262.800 235.800 ;
        RECT 263.600 224.200 264.400 237.800 ;
        RECT 265.200 224.200 266.000 237.800 ;
        RECT 276.500 232.400 277.100 249.600 ;
        RECT 298.800 244.200 299.600 257.800 ;
        RECT 300.400 244.200 301.200 257.800 ;
        RECT 302.000 244.200 302.800 257.800 ;
        RECT 303.600 246.200 304.400 257.800 ;
        RECT 305.300 256.400 305.900 259.600 ;
        RECT 305.200 255.600 306.000 256.400 ;
        RECT 305.300 238.400 305.900 255.600 ;
        RECT 306.800 246.200 307.600 257.800 ;
        RECT 308.400 253.600 309.200 254.400 ;
        RECT 308.500 240.400 309.100 253.600 ;
        RECT 310.000 246.200 310.800 257.800 ;
        RECT 311.600 244.200 312.400 257.800 ;
        RECT 313.200 244.200 314.000 257.800 ;
        RECT 318.100 250.400 318.700 261.600 ;
        RECT 322.800 259.600 323.600 260.400 ;
        RECT 322.900 258.400 323.500 259.600 ;
        RECT 322.800 257.600 323.600 258.400 ;
        RECT 321.200 255.600 322.000 256.400 ;
        RECT 318.000 249.600 318.800 250.400 ;
        RECT 308.400 239.600 309.200 240.400 ;
        RECT 276.400 231.600 277.200 232.400 ;
        RECT 276.500 230.400 277.100 231.600 ;
        RECT 270.000 229.600 270.800 230.400 ;
        RECT 276.400 229.600 277.200 230.400 ;
        RECT 282.800 227.600 283.600 228.400 ;
        RECT 276.400 225.600 277.200 226.400 ;
        RECT 286.000 223.600 286.800 224.400 ;
        RECT 295.600 224.200 296.400 237.800 ;
        RECT 297.200 224.200 298.000 237.800 ;
        RECT 298.800 224.200 299.600 237.800 ;
        RECT 302.000 237.600 302.800 238.400 ;
        RECT 305.200 237.600 306.000 238.400 ;
        RECT 300.400 224.200 301.200 235.800 ;
        RECT 302.100 226.400 302.700 237.600 ;
        RECT 302.000 225.600 302.800 226.400 ;
        RECT 284.400 221.600 285.200 222.400 ;
        RECT 257.200 219.600 258.000 220.400 ;
        RECT 263.600 219.600 264.400 220.400 ;
        RECT 250.800 217.600 251.600 218.400 ;
        RECT 255.600 217.600 256.400 218.400 ;
        RECT 247.600 205.600 248.400 206.400 ;
        RECT 247.600 203.600 248.400 204.400 ;
        RECT 247.700 192.400 248.300 203.600 ;
        RECT 247.600 191.600 248.400 192.400 ;
        RECT 246.100 189.700 248.300 190.300 ;
        RECT 244.400 185.600 245.200 186.400 ;
        RECT 244.500 178.400 245.100 185.600 ;
        RECT 244.400 177.600 245.200 178.400 ;
        RECT 244.400 175.600 245.200 176.400 ;
        RECT 246.000 173.600 246.800 174.400 ;
        RECT 247.700 174.300 248.300 189.700 ;
        RECT 249.200 189.600 250.000 190.400 ;
        RECT 249.300 186.400 249.900 189.600 ;
        RECT 249.200 185.600 250.000 186.400 ;
        RECT 250.900 174.400 251.500 217.600 ;
        RECT 255.700 206.400 256.300 217.600 ;
        RECT 255.600 205.600 256.400 206.400 ;
        RECT 252.400 191.600 253.200 192.400 ;
        RECT 252.500 190.400 253.100 191.600 ;
        RECT 252.400 189.600 253.200 190.400 ;
        RECT 254.000 189.600 254.800 190.400 ;
        RECT 254.100 178.400 254.700 189.600 ;
        RECT 254.000 177.600 254.800 178.400 ;
        RECT 255.700 174.400 256.300 205.600 ;
        RECT 257.200 204.200 258.000 217.800 ;
        RECT 258.800 204.200 259.600 217.800 ;
        RECT 260.400 204.200 261.200 217.800 ;
        RECT 262.000 206.200 262.800 217.800 ;
        RECT 263.700 216.400 264.300 219.600 ;
        RECT 263.600 215.600 264.400 216.400 ;
        RECT 265.200 206.200 266.000 217.800 ;
        RECT 266.800 213.600 267.600 214.400 ;
        RECT 266.900 210.400 267.500 213.600 ;
        RECT 266.800 209.600 267.600 210.400 ;
        RECT 268.400 206.200 269.200 217.800 ;
        RECT 270.000 204.200 270.800 217.800 ;
        RECT 271.600 204.200 272.400 217.800 ;
        RECT 276.400 211.600 277.200 212.400 ;
        RECT 258.800 201.600 259.600 202.400 ;
        RECT 258.900 178.400 259.500 201.600 ;
        RECT 268.200 189.600 269.200 190.400 ;
        RECT 266.800 187.600 267.600 188.400 ;
        RECT 262.000 185.600 262.800 186.400 ;
        RECT 263.600 185.600 264.400 186.400 ;
        RECT 260.400 179.600 261.200 180.400 ;
        RECT 258.800 177.600 259.600 178.400 ;
        RECT 257.200 175.600 258.000 176.400 ;
        RECT 257.300 174.400 257.900 175.600 ;
        RECT 260.500 174.400 261.100 179.600 ;
        RECT 247.700 173.700 249.900 174.300 ;
        RECT 249.300 172.400 249.900 173.700 ;
        RECT 250.800 173.600 251.600 174.400 ;
        RECT 255.600 173.600 256.400 174.400 ;
        RECT 257.200 173.600 258.000 174.400 ;
        RECT 260.400 173.600 261.200 174.400 ;
        RECT 249.200 171.600 250.000 172.400 ;
        RECT 246.000 169.600 246.800 170.400 ;
        RECT 246.100 162.400 246.700 169.600 ;
        RECT 242.800 161.600 243.600 162.400 ;
        RECT 246.000 161.600 246.800 162.400 ;
        RECT 239.600 157.600 240.400 158.400 ;
        RECT 238.000 145.600 238.800 146.400 ;
        RECT 239.600 144.200 240.400 155.800 ;
        RECT 241.200 144.200 242.000 157.800 ;
        RECT 242.800 144.200 243.600 157.800 ;
        RECT 244.400 144.200 245.200 157.800 ;
        RECT 249.300 142.400 249.900 171.600 ;
        RECT 250.900 170.400 251.500 173.600 ;
        RECT 262.100 172.400 262.700 185.600 ;
        RECT 252.400 171.600 253.200 172.400 ;
        RECT 262.000 171.600 262.800 172.400 ;
        RECT 252.500 170.400 253.100 171.600 ;
        RECT 250.800 169.600 251.600 170.400 ;
        RECT 252.400 169.600 253.200 170.400 ;
        RECT 257.200 169.600 258.000 170.400 ;
        RECT 252.500 166.300 253.100 169.600 ;
        RECT 250.900 165.700 253.100 166.300 ;
        RECT 233.200 141.600 234.000 142.400 ;
        RECT 249.200 141.600 250.000 142.400 ;
        RECT 228.400 139.600 229.200 140.400 ;
        RECT 228.500 134.400 229.100 139.600 ;
        RECT 226.800 133.600 227.600 134.400 ;
        RECT 228.400 133.600 229.200 134.400 ;
        RECT 233.300 132.400 233.900 141.600 ;
        RECT 250.900 138.400 251.500 165.700 ;
        RECT 255.600 153.600 256.400 154.400 ;
        RECT 255.700 152.400 256.300 153.600 ;
        RECT 255.600 151.600 256.400 152.400 ;
        RECT 254.000 143.600 254.800 144.400 ;
        RECT 250.800 137.600 251.600 138.400 ;
        RECT 254.100 136.400 254.700 143.600 ;
        RECT 242.800 135.600 243.600 136.400 ;
        RECT 246.000 135.600 246.800 136.400 ;
        RECT 252.400 135.600 253.200 136.400 ;
        RECT 254.000 135.600 254.800 136.400 ;
        RECT 238.000 133.600 238.800 134.400 ;
        RECT 249.200 133.600 250.000 134.400 ;
        RECT 252.400 133.600 253.200 134.400 ;
        RECT 238.100 132.400 238.700 133.600 ;
        RECT 254.100 132.400 254.700 135.600 ;
        RECT 226.800 131.600 227.600 132.400 ;
        RECT 230.000 131.600 230.800 132.400 ;
        RECT 231.600 131.600 232.400 132.400 ;
        RECT 233.200 131.600 234.000 132.400 ;
        RECT 238.000 131.600 238.800 132.400 ;
        RECT 249.200 131.600 250.000 132.400 ;
        RECT 254.000 131.600 254.800 132.400 ;
        RECT 220.400 129.600 221.200 130.400 ;
        RECT 222.000 129.600 222.800 130.400 ;
        RECT 214.000 119.600 214.800 120.400 ;
        RECT 214.100 116.400 214.700 119.600 ;
        RECT 222.000 117.600 222.800 118.400 ;
        RECT 214.000 115.600 214.800 116.400 ;
        RECT 212.400 113.600 213.200 114.400 ;
        RECT 212.500 112.400 213.100 113.600 ;
        RECT 212.400 111.600 213.200 112.400 ;
        RECT 214.100 106.400 214.700 115.600 ;
        RECT 222.100 112.400 222.700 117.600 ;
        RECT 226.900 112.400 227.500 131.600 ;
        RECT 222.000 111.600 222.800 112.400 ;
        RECT 226.800 111.600 227.600 112.400 ;
        RECT 220.400 109.600 221.200 110.400 ;
        RECT 215.600 107.600 216.400 108.400 ;
        RECT 214.000 105.600 214.800 106.400 ;
        RECT 222.100 100.400 222.700 111.600 ;
        RECT 225.200 109.600 226.000 110.400 ;
        RECT 225.200 107.600 226.000 108.400 ;
        RECT 225.300 106.400 225.900 107.600 ;
        RECT 225.200 105.600 226.000 106.400 ;
        RECT 222.000 99.600 222.800 100.400 ;
        RECT 225.300 98.400 225.900 105.600 ;
        RECT 218.800 97.600 219.600 98.400 ;
        RECT 225.200 97.600 226.000 98.400 ;
        RECT 218.900 96.400 219.500 97.600 ;
        RECT 231.700 96.400 232.300 131.600 ;
        RECT 249.300 130.400 249.900 131.600 ;
        RECT 233.200 129.600 234.000 130.400 ;
        RECT 249.200 129.600 250.000 130.400 ;
        RECT 236.400 127.600 237.200 128.400 ;
        RECT 236.500 110.400 237.100 127.600 ;
        RECT 246.000 123.600 246.800 124.400 ;
        RECT 246.100 114.400 246.700 123.600 ;
        RECT 246.000 113.600 246.800 114.400 ;
        RECT 239.600 111.600 240.400 112.400 ;
        RECT 247.600 111.600 248.400 112.400 ;
        RECT 236.400 109.600 237.200 110.400 ;
        RECT 233.200 108.300 234.000 108.400 ;
        RECT 233.200 107.700 235.500 108.300 ;
        RECT 233.200 107.600 234.000 107.700 ;
        RECT 233.200 105.600 234.000 106.400 ;
        RECT 234.900 102.400 235.500 107.700 ;
        RECT 239.700 106.400 240.300 111.600 ;
        RECT 249.300 108.400 249.900 129.600 ;
        RECT 250.800 123.600 251.600 124.400 ;
        RECT 250.900 118.400 251.500 123.600 ;
        RECT 250.800 117.600 251.600 118.400 ;
        RECT 252.400 113.600 253.200 114.400 ;
        RECT 252.500 110.400 253.100 113.600 ;
        RECT 255.700 110.400 256.300 151.600 ;
        RECT 257.300 136.400 257.900 169.600 ;
        RECT 258.800 165.600 259.600 166.400 ;
        RECT 258.900 158.400 259.500 165.600 ;
        RECT 258.800 157.600 259.600 158.400 ;
        RECT 260.400 149.600 261.200 150.400 ;
        RECT 260.500 148.400 261.100 149.600 ;
        RECT 260.400 147.600 261.200 148.400 ;
        RECT 262.000 147.600 262.800 148.400 ;
        RECT 257.200 135.600 258.000 136.400 ;
        RECT 260.500 134.400 261.100 147.600 ;
        RECT 263.700 146.400 264.300 185.600 ;
        RECT 268.400 183.600 269.200 184.400 ;
        RECT 278.000 184.200 278.800 197.800 ;
        RECT 279.600 184.200 280.400 197.800 ;
        RECT 281.200 184.200 282.000 197.800 ;
        RECT 282.800 184.200 283.600 195.800 ;
        RECT 284.500 186.400 285.100 221.600 ;
        RECT 286.100 216.400 286.700 223.600 ;
        RECT 302.100 222.400 302.700 225.600 ;
        RECT 303.600 224.200 304.400 235.800 ;
        RECT 305.200 227.600 306.000 228.400 ;
        RECT 305.300 226.400 305.900 227.600 ;
        RECT 305.200 225.600 306.000 226.400 ;
        RECT 306.800 224.200 307.600 235.800 ;
        RECT 308.400 224.200 309.200 237.800 ;
        RECT 310.000 224.200 310.800 237.800 ;
        RECT 311.600 231.200 312.400 232.400 ;
        RECT 302.000 221.600 302.800 222.400 ;
        RECT 308.400 221.600 309.200 222.400 ;
        RECT 289.200 219.600 290.000 220.400 ;
        RECT 289.300 218.400 289.900 219.600 ;
        RECT 289.200 217.600 290.000 218.400 ;
        RECT 286.000 215.600 286.800 216.400 ;
        RECT 292.400 215.600 293.200 216.400 ;
        RECT 286.100 214.400 286.700 215.600 ;
        RECT 286.000 213.600 286.800 214.400 ;
        RECT 292.400 203.600 293.200 204.400 ;
        RECT 302.000 204.200 302.800 217.800 ;
        RECT 303.600 204.200 304.400 217.800 ;
        RECT 305.200 204.200 306.000 217.800 ;
        RECT 306.800 206.200 307.600 217.800 ;
        RECT 308.500 216.400 309.100 221.600 ;
        RECT 308.400 215.600 309.200 216.400 ;
        RECT 310.000 206.200 310.800 217.800 ;
        RECT 311.600 213.600 312.400 214.400 ;
        RECT 313.200 206.200 314.000 217.800 ;
        RECT 314.800 204.200 315.600 217.800 ;
        RECT 316.400 204.200 317.200 217.800 ;
        RECT 318.100 212.400 318.700 249.600 ;
        RECT 321.300 238.400 321.900 255.600 ;
        RECT 327.700 254.400 328.300 261.600 ;
        RECT 322.800 253.600 323.600 254.400 ;
        RECT 327.600 253.600 328.400 254.400 ;
        RECT 329.200 253.600 330.000 254.400 ;
        RECT 322.900 250.400 323.500 253.600 ;
        RECT 329.200 251.600 330.000 252.400 ;
        RECT 329.300 250.400 329.900 251.600 ;
        RECT 322.800 249.600 323.600 250.400 ;
        RECT 329.200 249.600 330.000 250.400 ;
        RECT 321.200 237.600 322.000 238.400 ;
        RECT 324.400 231.600 325.200 232.400 ;
        RECT 321.200 229.600 322.000 230.400 ;
        RECT 324.500 228.400 325.100 231.600 ;
        RECT 327.600 229.600 328.400 230.400 ;
        RECT 329.300 230.300 329.900 249.600 ;
        RECT 330.900 236.400 331.500 287.600 ;
        RECT 332.500 270.400 333.100 313.600 ;
        RECT 334.100 310.300 334.700 343.700 ;
        RECT 342.100 340.400 342.700 349.600 ;
        RECT 345.200 347.600 346.000 348.400 ;
        RECT 351.600 347.600 352.400 348.400 ;
        RECT 345.200 345.600 346.000 346.400 ;
        RECT 345.300 342.400 345.900 345.600 ;
        RECT 351.600 343.600 352.400 344.400 ;
        RECT 345.200 341.600 346.000 342.400 ;
        RECT 337.200 339.600 338.000 340.400 ;
        RECT 342.000 339.600 342.800 340.400 ;
        RECT 337.300 314.400 337.900 339.600 ;
        RECT 351.700 338.400 352.300 343.600 ;
        RECT 351.600 337.600 352.400 338.400 ;
        RECT 353.300 334.400 353.900 349.600 ;
        RECT 356.500 340.400 357.100 351.600 ;
        RECT 372.500 350.400 373.100 351.600 ;
        RECT 361.200 349.600 362.000 350.400 ;
        RECT 366.000 349.600 366.800 350.400 ;
        RECT 369.200 349.600 370.000 350.400 ;
        RECT 372.400 349.600 373.200 350.400 ;
        RECT 374.000 349.600 374.800 350.400 ;
        RECT 375.600 349.600 376.400 350.400 ;
        RECT 354.800 339.600 355.600 340.400 ;
        RECT 356.400 339.600 357.200 340.400 ;
        RECT 354.900 334.400 355.500 339.600 ;
        RECT 356.400 335.600 357.200 336.400 ;
        RECT 343.600 333.600 344.400 334.400 ;
        RECT 348.400 333.600 349.200 334.400 ;
        RECT 353.200 333.600 354.000 334.400 ;
        RECT 354.800 333.600 355.600 334.400 ;
        RECT 343.700 332.400 344.300 333.600 ;
        RECT 343.600 331.600 344.400 332.400 ;
        RECT 343.600 327.600 344.400 328.400 ;
        RECT 335.600 313.600 336.400 314.400 ;
        RECT 337.200 313.600 338.000 314.400 ;
        RECT 335.600 310.300 336.400 310.400 ;
        RECT 334.100 309.700 336.400 310.300 ;
        RECT 335.600 309.600 336.400 309.700 ;
        RECT 337.300 308.400 337.900 313.600 ;
        RECT 337.200 307.600 338.000 308.400 ;
        RECT 340.400 307.600 341.200 308.400 ;
        RECT 340.400 305.600 341.200 306.400 ;
        RECT 343.700 300.400 344.300 327.600 ;
        RECT 346.800 323.600 347.600 324.400 ;
        RECT 346.900 318.400 347.500 323.600 ;
        RECT 346.800 317.600 347.600 318.400 ;
        RECT 346.900 310.400 347.500 317.600 ;
        RECT 348.500 314.400 349.100 333.600 ;
        RECT 354.900 332.400 355.500 333.600 ;
        RECT 353.200 331.600 354.000 332.400 ;
        RECT 354.800 331.600 355.600 332.400 ;
        RECT 351.600 329.600 352.400 330.400 ;
        RECT 348.400 313.600 349.200 314.400 ;
        RECT 348.400 311.600 349.200 312.400 ;
        RECT 345.200 309.600 346.000 310.400 ;
        RECT 346.800 309.600 347.600 310.400 ;
        RECT 348.400 309.600 349.200 310.400 ;
        RECT 343.600 299.600 344.400 300.400 ;
        RECT 345.300 298.400 345.900 309.600 ;
        RECT 346.800 307.600 347.600 308.400 ;
        RECT 346.900 304.400 347.500 307.600 ;
        RECT 351.700 306.400 352.300 329.600 ;
        RECT 353.300 322.400 353.900 331.600 ;
        RECT 358.000 329.600 358.800 330.400 ;
        RECT 359.600 329.600 360.400 330.400 ;
        RECT 356.400 325.600 357.200 326.400 ;
        RECT 353.200 321.600 354.000 322.400 ;
        RECT 353.200 311.600 354.000 312.400 ;
        RECT 353.300 308.400 353.900 311.600 ;
        RECT 356.500 308.400 357.100 325.600 ;
        RECT 358.100 312.400 358.700 329.600 ;
        RECT 361.300 328.400 361.900 349.600 ;
        RECT 362.800 347.600 363.600 348.400 ;
        RECT 364.400 347.600 365.200 348.400 ;
        RECT 362.900 338.400 363.500 347.600 ;
        RECT 364.500 346.400 365.100 347.600 ;
        RECT 364.400 345.600 365.200 346.400 ;
        RECT 366.100 344.400 366.700 349.600 ;
        RECT 366.000 343.600 366.800 344.400 ;
        RECT 367.600 343.600 368.400 344.400 ;
        RECT 364.400 341.600 365.200 342.400 ;
        RECT 364.500 340.300 365.100 341.600 ;
        RECT 367.700 340.300 368.300 343.600 ;
        RECT 369.300 342.300 369.900 349.600 ;
        RECT 370.800 347.600 371.600 348.400 ;
        RECT 370.900 344.400 371.500 347.600 ;
        RECT 370.800 343.600 371.600 344.400 ;
        RECT 369.300 341.700 373.100 342.300 ;
        RECT 364.500 339.700 368.300 340.300 ;
        RECT 362.800 337.600 363.600 338.400 ;
        RECT 364.400 335.600 365.200 336.400 ;
        RECT 364.500 334.400 365.100 335.600 ;
        RECT 364.400 333.600 365.200 334.400 ;
        RECT 372.500 334.300 373.100 341.700 ;
        RECT 374.100 336.400 374.700 349.600 ;
        RECT 375.700 336.400 376.300 349.600 ;
        RECT 377.200 347.600 378.000 348.400 ;
        RECT 374.000 335.600 374.800 336.400 ;
        RECT 375.600 335.600 376.400 336.400 ;
        RECT 374.000 334.300 374.800 334.400 ;
        RECT 372.500 333.700 374.800 334.300 ;
        RECT 374.000 333.600 374.800 333.700 ;
        RECT 375.700 332.400 376.300 335.600 ;
        RECT 362.800 331.600 363.600 332.400 ;
        RECT 370.800 331.600 371.600 332.400 ;
        RECT 375.600 331.600 376.400 332.400 ;
        RECT 366.000 329.600 366.800 330.400 ;
        RECT 359.600 327.600 360.400 328.400 ;
        RECT 361.200 327.600 362.000 328.400 ;
        RECT 359.700 318.400 360.300 327.600 ;
        RECT 366.100 322.400 366.700 329.600 ;
        RECT 370.900 324.400 371.500 331.600 ;
        RECT 375.600 329.600 376.400 330.400 ;
        RECT 375.700 328.400 376.300 329.600 ;
        RECT 375.600 327.600 376.400 328.400 ;
        RECT 369.200 323.600 370.000 324.400 ;
        RECT 370.800 323.600 371.600 324.400 ;
        RECT 364.400 321.600 365.200 322.400 ;
        RECT 366.000 321.600 366.800 322.400 ;
        RECT 369.200 321.600 370.000 322.400 ;
        RECT 359.600 317.600 360.400 318.400 ;
        RECT 361.200 313.600 362.000 314.400 ;
        RECT 361.300 312.400 361.900 313.600 ;
        RECT 358.000 311.600 358.800 312.400 ;
        RECT 361.200 311.600 362.000 312.400 ;
        RECT 359.600 309.600 360.400 310.400 ;
        RECT 353.200 307.600 354.000 308.400 ;
        RECT 356.400 307.600 357.200 308.400 ;
        RECT 351.600 305.600 352.400 306.400 ;
        RECT 346.800 303.600 347.600 304.400 ;
        RECT 345.200 297.600 346.000 298.400 ;
        RECT 351.700 294.400 352.300 305.600 ;
        RECT 359.700 298.400 360.300 309.600 ;
        RECT 364.500 306.400 365.100 321.600 ;
        RECT 369.300 318.400 369.900 321.600 ;
        RECT 375.700 320.400 376.300 327.600 ;
        RECT 375.600 319.600 376.400 320.400 ;
        RECT 369.200 317.600 370.000 318.400 ;
        RECT 370.800 313.600 371.600 314.400 ;
        RECT 375.600 313.600 376.400 314.400 ;
        RECT 369.200 307.600 370.000 308.400 ;
        RECT 364.400 305.600 365.200 306.400 ;
        RECT 361.200 303.600 362.000 304.400 ;
        RECT 362.800 303.600 363.600 304.400 ;
        RECT 359.600 297.600 360.400 298.400 ;
        RECT 361.300 296.400 361.900 303.600 ;
        RECT 362.900 298.400 363.500 303.600 ;
        RECT 370.900 298.400 371.500 313.600 ;
        RECT 375.700 312.400 376.300 313.600 ;
        RECT 375.600 311.600 376.400 312.400 ;
        RECT 375.600 309.600 376.400 310.400 ;
        RECT 372.400 307.600 373.200 308.400 ;
        RECT 372.500 304.400 373.100 307.600 ;
        RECT 377.300 306.400 377.900 347.600 ;
        RECT 378.900 346.400 379.500 353.600 ;
        RECT 378.800 345.600 379.600 346.400 ;
        RECT 380.500 334.400 381.100 363.600 ;
        RECT 382.000 357.600 382.800 358.400 ;
        RECT 382.100 348.400 382.700 357.600 ;
        RECT 386.900 356.400 387.500 371.600 ;
        RECT 388.400 369.600 389.200 370.400 ;
        RECT 388.500 368.400 389.100 369.600 ;
        RECT 388.400 367.600 389.200 368.400 ;
        RECT 390.000 367.600 390.800 368.400 ;
        RECT 390.100 362.400 390.700 367.600 ;
        RECT 399.700 366.400 400.300 371.600 ;
        RECT 399.600 365.600 400.400 366.400 ;
        RECT 402.800 364.200 403.600 377.800 ;
        RECT 404.400 364.200 405.200 377.800 ;
        RECT 406.000 366.200 406.800 377.800 ;
        RECT 407.600 373.600 408.400 374.400 ;
        RECT 407.700 368.400 408.300 373.600 ;
        RECT 407.600 367.600 408.400 368.400 ;
        RECT 409.200 366.200 410.000 377.800 ;
        RECT 410.800 375.600 411.600 376.400 ;
        RECT 410.900 364.400 411.500 375.600 ;
        RECT 412.400 366.200 413.200 377.800 ;
        RECT 410.800 363.600 411.600 364.400 ;
        RECT 414.000 364.200 414.800 377.800 ;
        RECT 415.600 364.200 416.400 377.800 ;
        RECT 417.200 364.200 418.000 377.800 ;
        RECT 426.800 373.600 427.800 374.400 ;
        RECT 446.000 373.600 446.800 374.400 ;
        RECT 437.800 371.600 438.800 372.400 ;
        RECT 390.000 361.600 390.800 362.400 ;
        RECT 391.600 361.600 392.400 362.400 ;
        RECT 394.800 361.600 395.600 362.400 ;
        RECT 412.400 361.600 413.200 362.400 ;
        RECT 388.400 359.600 389.200 360.400 ;
        RECT 388.500 358.400 389.100 359.600 ;
        RECT 388.400 357.600 389.200 358.400 ;
        RECT 386.800 355.600 387.600 356.400 ;
        RECT 383.600 353.600 384.400 354.400 ;
        RECT 383.700 350.400 384.300 353.600 ;
        RECT 383.600 349.600 384.400 350.400 ;
        RECT 386.900 348.400 387.500 355.600 ;
        RECT 391.700 348.400 392.300 361.600 ;
        RECT 393.200 359.600 394.000 360.400 ;
        RECT 393.300 350.400 393.900 359.600 ;
        RECT 394.900 356.300 395.500 361.600 ;
        RECT 398.000 359.600 398.800 360.400 ;
        RECT 406.000 359.600 406.800 360.400 ;
        RECT 396.400 358.300 397.200 358.400 ;
        RECT 398.100 358.300 398.700 359.600 ;
        RECT 406.100 358.400 406.700 359.600 ;
        RECT 396.400 357.700 398.700 358.300 ;
        RECT 396.400 357.600 397.200 357.700 ;
        RECT 406.000 357.600 406.800 358.400 ;
        RECT 394.900 355.700 398.700 356.300 ;
        RECT 396.400 351.600 397.200 352.400 ;
        RECT 393.200 349.600 394.000 350.400 ;
        RECT 394.800 349.600 395.600 350.400 ;
        RECT 382.000 347.600 382.800 348.400 ;
        RECT 386.800 347.600 387.600 348.400 ;
        RECT 391.600 347.600 392.400 348.400 ;
        RECT 385.200 345.600 386.000 346.400 ;
        RECT 388.400 345.600 389.200 346.400 ;
        RECT 394.900 346.300 395.500 349.600 ;
        RECT 396.500 348.400 397.100 351.600 ;
        RECT 398.100 350.400 398.700 355.700 ;
        RECT 399.700 355.700 408.300 356.300 ;
        RECT 399.700 354.400 400.300 355.700 ;
        RECT 407.700 354.400 408.300 355.700 ;
        RECT 409.200 355.600 410.000 356.400 ;
        RECT 399.600 353.600 400.400 354.400 ;
        RECT 401.200 353.600 402.000 354.400 ;
        RECT 406.000 353.600 406.800 354.400 ;
        RECT 407.600 353.600 408.400 354.400 ;
        RECT 401.300 350.400 401.900 353.600 ;
        RECT 402.800 351.600 403.600 352.400 ;
        RECT 398.000 349.600 398.800 350.400 ;
        RECT 401.200 349.600 402.000 350.400 ;
        RECT 396.400 347.600 397.200 348.400 ;
        RECT 394.900 345.700 397.100 346.300 ;
        RECT 388.500 338.400 389.100 345.600 ;
        RECT 396.500 344.400 397.100 345.700 ;
        RECT 399.600 345.600 400.400 346.400 ;
        RECT 394.800 343.600 395.600 344.400 ;
        RECT 396.400 343.600 397.200 344.400 ;
        RECT 394.900 338.400 395.500 343.600 ;
        RECT 399.700 338.400 400.300 345.600 ;
        RECT 401.300 344.400 401.900 349.600 ;
        RECT 402.900 348.400 403.500 351.600 ;
        RECT 406.100 350.400 406.700 353.600 ;
        RECT 407.600 351.600 408.400 352.400 ;
        RECT 404.400 349.600 405.200 350.400 ;
        RECT 406.000 349.600 406.800 350.400 ;
        RECT 402.800 347.600 403.600 348.400 ;
        RECT 401.200 343.600 402.000 344.400 ;
        RECT 382.000 337.600 382.800 338.400 ;
        RECT 388.400 337.600 389.200 338.400 ;
        RECT 394.800 337.600 395.600 338.400 ;
        RECT 399.600 337.600 400.400 338.400 ;
        RECT 391.600 335.600 392.400 336.400 ;
        RECT 398.000 335.600 398.800 336.400 ;
        RECT 380.400 333.600 381.200 334.400 ;
        RECT 391.700 332.400 392.300 335.600 ;
        RECT 398.100 334.400 398.700 335.600 ;
        RECT 393.200 333.600 394.000 334.400 ;
        RECT 398.000 333.600 398.800 334.400 ;
        RECT 402.800 333.600 403.600 334.400 ;
        RECT 382.000 331.600 382.800 332.400 ;
        RECT 391.600 331.600 392.400 332.400 ;
        RECT 378.800 325.600 379.600 326.400 ;
        RECT 378.900 310.400 379.500 325.600 ;
        RECT 378.800 309.600 379.600 310.400 ;
        RECT 382.100 308.400 382.700 331.600 ;
        RECT 383.600 329.600 384.400 330.400 ;
        RECT 388.400 329.600 389.200 330.400 ;
        RECT 393.300 324.400 393.900 333.600 ;
        RECT 394.800 329.600 395.600 330.400 ;
        RECT 398.000 329.600 398.800 330.400 ;
        RECT 386.800 323.600 387.600 324.400 ;
        RECT 393.200 323.600 394.000 324.400 ;
        RECT 386.900 314.400 387.500 323.600 ;
        RECT 398.100 314.400 398.700 329.600 ;
        RECT 399.600 327.600 400.400 328.400 ;
        RECT 399.700 318.400 400.300 327.600 ;
        RECT 401.200 325.600 402.000 326.400 ;
        RECT 402.900 320.400 403.500 333.600 ;
        RECT 404.500 326.400 405.100 349.600 ;
        RECT 407.700 346.400 408.300 351.600 ;
        RECT 409.300 346.400 409.900 355.600 ;
        RECT 412.500 354.400 413.100 361.600 ;
        RECT 446.100 358.400 446.700 373.600 ;
        RECT 447.600 364.200 448.400 377.800 ;
        RECT 449.200 364.200 450.000 377.800 ;
        RECT 450.800 364.200 451.600 377.800 ;
        RECT 452.400 366.200 453.200 377.800 ;
        RECT 454.000 375.600 454.800 376.400 ;
        RECT 441.200 357.600 442.000 358.400 ;
        RECT 446.000 357.600 446.800 358.400 ;
        RECT 412.400 353.600 413.200 354.400 ;
        RECT 420.400 353.600 421.200 354.400 ;
        RECT 420.500 352.400 421.100 353.600 ;
        RECT 441.300 352.400 441.900 357.600 ;
        RECT 454.100 354.400 454.700 375.600 ;
        RECT 455.600 366.200 456.400 377.800 ;
        RECT 457.200 373.600 458.000 374.400 ;
        RECT 457.300 358.400 457.900 373.600 ;
        RECT 458.800 366.200 459.600 377.800 ;
        RECT 460.400 364.200 461.200 377.800 ;
        RECT 462.000 364.200 462.800 377.800 ;
        RECT 463.600 371.600 464.400 372.400 ;
        RECT 474.800 371.600 475.600 372.400 ;
        RECT 457.200 357.600 458.000 358.400 ;
        RECT 444.400 353.600 445.200 354.400 ;
        RECT 449.200 353.600 450.000 354.400 ;
        RECT 454.000 353.600 454.800 354.400 ;
        RECT 420.400 351.600 421.200 352.400 ;
        RECT 434.800 351.600 435.600 352.400 ;
        RECT 439.600 351.600 440.400 352.400 ;
        RECT 441.200 351.600 442.000 352.400 ;
        RECT 450.800 351.600 451.600 352.400 ;
        RECT 452.400 351.600 453.200 352.400 ;
        RECT 462.000 351.600 462.800 352.400 ;
        RECT 412.400 349.600 413.200 350.400 ;
        RECT 420.400 349.600 421.200 350.400 ;
        RECT 422.000 349.600 422.800 350.400 ;
        RECT 410.800 347.600 411.600 348.400 ;
        RECT 420.500 346.400 421.100 349.600 ;
        RECT 407.600 345.600 408.400 346.400 ;
        RECT 409.200 345.600 410.000 346.400 ;
        RECT 420.400 345.600 421.200 346.400 ;
        RECT 409.200 343.600 410.000 344.400 ;
        RECT 410.800 343.600 411.600 344.400 ;
        RECT 409.300 334.400 409.900 343.600 ;
        RECT 412.400 337.600 413.200 338.400 ;
        RECT 422.100 336.400 422.700 349.600 ;
        RECT 423.600 345.600 424.400 346.400 ;
        RECT 423.700 336.400 424.300 345.600 ;
        RECT 428.400 337.600 429.200 338.400 ;
        RECT 417.200 335.600 418.000 336.400 ;
        RECT 418.800 335.600 419.600 336.400 ;
        RECT 422.000 335.600 422.800 336.400 ;
        RECT 423.600 335.600 424.400 336.400 ;
        RECT 417.300 334.400 417.900 335.600 ;
        RECT 409.200 333.600 410.000 334.400 ;
        RECT 417.200 333.600 418.000 334.400 ;
        RECT 407.600 331.600 408.400 332.400 ;
        RECT 414.000 331.600 414.800 332.400 ;
        RECT 407.700 328.400 408.300 331.600 ;
        RECT 409.200 329.600 410.000 330.400 ;
        RECT 407.600 327.600 408.400 328.400 ;
        RECT 404.400 325.600 405.200 326.400 ;
        RECT 407.600 326.300 408.400 326.400 ;
        RECT 409.300 326.300 409.900 329.600 ;
        RECT 407.600 325.700 409.900 326.300 ;
        RECT 407.600 325.600 408.400 325.700 ;
        RECT 412.400 323.600 413.200 324.400 ;
        RECT 407.600 321.600 408.400 322.400 ;
        RECT 402.800 319.600 403.600 320.400 ;
        RECT 407.700 318.400 408.300 321.600 ;
        RECT 409.200 319.600 410.000 320.400 ;
        RECT 399.600 317.600 400.400 318.400 ;
        RECT 407.600 317.600 408.400 318.400 ;
        RECT 386.800 313.600 387.600 314.400 ;
        RECT 398.000 313.600 398.800 314.400 ;
        RECT 401.200 313.600 402.000 314.400 ;
        RECT 406.000 313.600 406.800 314.400 ;
        RECT 407.600 313.600 408.400 314.400 ;
        RECT 383.600 311.600 384.400 312.400 ;
        RECT 383.700 310.400 384.300 311.600 ;
        RECT 386.900 310.400 387.500 313.600 ;
        RECT 407.700 312.400 408.300 313.600 ;
        RECT 409.300 312.400 409.900 319.600 ;
        RECT 391.600 312.300 392.400 312.400 ;
        RECT 398.000 312.300 398.800 312.400 ;
        RECT 391.600 311.700 398.800 312.300 ;
        RECT 391.600 311.600 392.400 311.700 ;
        RECT 398.000 311.600 398.800 311.700 ;
        RECT 407.600 311.600 408.400 312.400 ;
        RECT 409.200 312.300 410.000 312.400 ;
        RECT 409.200 311.700 411.500 312.300 ;
        RECT 409.200 311.600 410.000 311.700 ;
        RECT 383.600 309.600 384.400 310.400 ;
        RECT 386.800 309.600 387.600 310.400 ;
        RECT 394.800 309.600 395.600 310.400 ;
        RECT 399.600 309.600 400.400 310.400 ;
        RECT 407.600 309.600 408.400 310.400 ;
        RECT 378.800 307.600 379.600 308.400 ;
        RECT 382.000 307.600 382.800 308.400 ;
        RECT 385.200 307.600 386.000 308.400 ;
        RECT 390.000 307.600 390.800 308.400 ;
        RECT 396.400 307.600 397.200 308.400 ;
        RECT 375.600 305.600 376.400 306.400 ;
        RECT 377.200 305.600 378.000 306.400 ;
        RECT 372.400 303.600 373.200 304.400 ;
        RECT 378.900 298.400 379.500 307.600 ;
        RECT 390.000 305.600 390.800 306.400 ;
        RECT 390.100 300.400 390.700 305.600 ;
        RECT 390.000 299.600 390.800 300.400 ;
        RECT 396.500 298.400 397.100 307.600 ;
        RECT 399.700 306.400 400.300 309.600 ;
        RECT 407.700 308.400 408.300 309.600 ;
        RECT 406.000 307.600 406.800 308.400 ;
        RECT 407.600 307.600 408.400 308.400 ;
        RECT 399.600 305.600 400.400 306.400 ;
        RECT 406.100 298.400 406.700 307.600 ;
        RECT 409.200 299.600 410.000 300.400 ;
        RECT 362.800 297.600 363.600 298.400 ;
        RECT 370.800 297.600 371.600 298.400 ;
        RECT 374.000 297.600 374.800 298.400 ;
        RECT 378.800 297.600 379.600 298.400 ;
        RECT 383.600 297.600 384.400 298.400 ;
        RECT 396.400 297.600 397.200 298.400 ;
        RECT 398.000 297.600 398.800 298.400 ;
        RECT 406.000 297.600 406.800 298.400 ;
        RECT 354.800 295.600 355.600 296.400 ;
        RECT 361.200 295.600 362.000 296.400 ;
        RECT 366.000 295.600 366.800 296.400 ;
        RECT 369.200 295.600 370.000 296.400 ;
        RECT 375.600 295.600 376.400 296.400 ;
        RECT 337.200 293.600 338.000 294.400 ;
        RECT 346.800 293.600 347.600 294.400 ;
        RECT 351.600 293.600 352.400 294.400 ;
        RECT 353.200 293.600 354.000 294.400 ;
        RECT 346.900 292.400 347.500 293.600 ;
        RECT 335.600 291.600 336.400 292.400 ;
        RECT 346.800 291.600 347.600 292.400 ;
        RECT 335.700 290.400 336.300 291.600 ;
        RECT 335.600 289.600 336.400 290.400 ;
        RECT 340.400 289.600 341.200 290.400 ;
        RECT 345.200 289.600 346.000 290.400 ;
        RECT 335.600 273.600 336.400 274.400 ;
        RECT 338.800 271.600 339.600 272.400 ;
        RECT 332.400 269.600 333.200 270.400 ;
        RECT 337.200 259.600 338.000 260.400 ;
        RECT 337.300 258.400 337.900 259.600 ;
        RECT 337.200 257.600 338.000 258.400 ;
        RECT 338.900 254.400 339.500 271.600 ;
        RECT 343.600 269.600 344.400 270.400 ;
        RECT 342.000 267.600 342.800 268.400 ;
        RECT 340.400 263.600 341.200 264.400 ;
        RECT 340.500 262.400 341.100 263.600 ;
        RECT 340.400 261.600 341.200 262.400 ;
        RECT 342.100 260.400 342.700 267.600 ;
        RECT 342.000 259.600 342.800 260.400 ;
        RECT 340.400 257.600 341.200 258.400 ;
        RECT 340.500 256.400 341.100 257.600 ;
        RECT 340.400 255.600 341.200 256.400 ;
        RECT 334.000 253.600 334.800 254.400 ;
        RECT 338.800 253.600 339.600 254.400 ;
        RECT 330.800 235.600 331.600 236.400 ;
        RECT 330.800 231.600 331.600 232.400 ;
        RECT 332.400 231.600 333.200 232.400 ;
        RECT 332.500 230.400 333.100 231.600 ;
        RECT 329.300 229.700 331.500 230.300 ;
        RECT 319.600 227.600 320.400 228.400 ;
        RECT 322.800 227.600 323.600 228.400 ;
        RECT 324.400 227.600 325.200 228.400 ;
        RECT 326.000 227.600 326.800 228.400 ;
        RECT 329.200 227.600 330.000 228.400 ;
        RECT 322.900 222.400 323.500 227.600 ;
        RECT 319.600 221.600 320.400 222.400 ;
        RECT 322.800 221.600 323.600 222.400 ;
        RECT 318.000 211.600 318.800 212.400 ;
        RECT 318.100 210.800 318.700 211.600 ;
        RECT 318.000 210.000 318.800 210.800 ;
        RECT 284.400 185.600 285.200 186.400 ;
        RECT 286.000 184.200 286.800 195.800 ;
        RECT 287.600 187.600 288.400 188.400 ;
        RECT 289.200 184.200 290.000 195.800 ;
        RECT 290.800 184.200 291.600 197.800 ;
        RECT 292.400 184.200 293.200 197.800 ;
        RECT 295.600 195.600 296.400 196.400 ;
        RECT 266.800 175.600 267.600 176.400 ;
        RECT 265.200 173.600 266.000 174.400 ;
        RECT 266.900 172.400 267.500 175.600 ;
        RECT 266.800 171.600 267.600 172.400 ;
        RECT 268.500 170.400 269.100 183.600 ;
        RECT 270.000 181.600 270.800 182.400 ;
        RECT 270.100 176.400 270.700 181.600 ;
        RECT 271.600 177.600 272.400 178.400 ;
        RECT 270.000 175.600 270.800 176.400 ;
        RECT 281.300 175.700 286.700 176.300 ;
        RECT 273.200 173.600 274.000 174.400 ;
        RECT 281.300 172.400 281.900 175.700 ;
        RECT 286.100 174.400 286.700 175.700 ;
        RECT 289.200 175.600 290.000 176.400 ;
        RECT 290.800 175.600 291.600 176.400 ;
        RECT 289.300 174.400 289.900 175.600 ;
        RECT 282.800 173.600 283.600 174.400 ;
        RECT 286.000 173.600 286.800 174.400 ;
        RECT 289.200 173.600 290.000 174.400 ;
        RECT 270.000 171.600 270.800 172.400 ;
        RECT 281.200 171.600 282.000 172.400 ;
        RECT 284.400 171.600 285.200 172.400 ;
        RECT 292.400 171.600 293.200 172.400 ;
        RECT 268.400 169.600 269.200 170.400 ;
        RECT 265.200 167.600 266.000 168.400 ;
        RECT 268.500 152.400 269.100 169.600 ;
        RECT 270.100 158.400 270.700 171.600 ;
        RECT 292.500 170.400 293.100 171.600 ;
        RECT 287.600 169.600 288.400 170.400 ;
        RECT 292.400 169.600 293.200 170.400 ;
        RECT 286.000 167.600 286.800 168.400 ;
        RECT 286.100 158.400 286.700 167.600 ;
        RECT 270.000 157.600 270.800 158.400 ;
        RECT 286.000 157.600 286.800 158.400 ;
        RECT 290.800 157.600 291.600 158.400 ;
        RECT 271.600 153.600 272.400 154.400 ;
        RECT 279.600 153.600 280.400 154.400 ;
        RECT 268.400 151.600 269.200 152.400 ;
        RECT 266.800 149.600 267.600 150.400 ;
        RECT 270.000 149.600 270.800 150.400 ;
        RECT 266.900 148.400 267.500 149.600 ;
        RECT 279.700 148.400 280.300 153.600 ;
        RECT 290.900 150.400 291.500 157.600 ;
        RECT 295.700 150.400 296.300 195.600 ;
        RECT 297.200 189.600 298.000 190.400 ;
        RECT 297.300 182.400 297.900 189.600 ;
        RECT 303.600 183.600 304.400 184.400 ;
        RECT 313.200 184.200 314.000 197.800 ;
        RECT 314.800 184.200 315.600 197.800 ;
        RECT 316.400 184.200 317.200 197.800 ;
        RECT 318.000 184.200 318.800 195.800 ;
        RECT 319.700 186.400 320.300 221.600 ;
        RECT 326.100 220.400 326.700 227.600 ;
        RECT 329.300 226.400 329.900 227.600 ;
        RECT 329.200 225.600 330.000 226.400 ;
        RECT 326.000 219.600 326.800 220.400 ;
        RECT 326.000 215.600 326.800 216.400 ;
        RECT 330.900 212.400 331.500 229.700 ;
        RECT 332.400 229.600 333.200 230.400 ;
        RECT 334.100 228.400 334.700 253.600 ;
        RECT 345.300 252.400 345.900 289.600 ;
        RECT 346.900 272.400 347.500 291.600 ;
        RECT 354.900 276.400 355.500 295.600 ;
        RECT 367.600 293.600 368.400 294.400 ;
        RECT 369.300 292.400 369.900 295.600 ;
        RECT 372.400 293.600 373.200 294.400 ;
        RECT 356.400 291.600 357.200 292.400 ;
        RECT 369.200 291.600 370.000 292.400 ;
        RECT 356.500 288.400 357.100 291.600 ;
        RECT 372.500 288.400 373.100 293.600 ;
        RECT 375.700 292.400 376.300 295.600 ;
        RECT 377.200 293.600 378.000 294.400 ;
        RECT 375.600 291.600 376.400 292.400 ;
        RECT 377.200 289.600 378.000 290.400 ;
        RECT 356.400 287.600 357.200 288.400 ;
        RECT 372.400 287.600 373.200 288.400 ;
        RECT 354.800 275.600 355.600 276.400 ;
        RECT 346.800 271.600 347.600 272.400 ;
        RECT 354.800 271.200 355.600 272.000 ;
        RECT 354.900 270.400 355.500 271.200 ;
        RECT 354.800 269.600 355.600 270.400 ;
        RECT 346.800 263.600 347.600 264.400 ;
        RECT 346.900 256.400 347.500 263.600 ;
        RECT 348.400 261.600 349.200 262.400 ;
        RECT 348.500 258.400 349.100 261.600 ;
        RECT 348.400 257.600 349.200 258.400 ;
        RECT 346.800 255.600 347.600 256.400 ;
        RECT 354.900 252.400 355.500 269.600 ;
        RECT 356.400 264.200 357.200 277.800 ;
        RECT 358.000 264.200 358.800 277.800 ;
        RECT 359.600 264.200 360.400 275.800 ;
        RECT 361.200 267.600 362.000 268.400 ;
        RECT 361.300 262.400 361.900 267.600 ;
        RECT 362.800 264.200 363.600 275.800 ;
        RECT 364.400 265.600 365.200 266.400 ;
        RECT 366.000 264.200 366.800 275.800 ;
        RECT 367.600 264.200 368.400 277.800 ;
        RECT 369.200 264.200 370.000 277.800 ;
        RECT 370.800 264.200 371.600 277.800 ;
        RECT 361.200 261.600 362.000 262.400 ;
        RECT 375.600 259.600 376.400 260.400 ;
        RECT 345.200 251.600 346.000 252.400 ;
        RECT 354.800 251.600 355.600 252.400 ;
        RECT 354.900 250.400 355.500 251.600 ;
        RECT 348.400 250.300 349.200 250.400 ;
        RECT 346.900 249.700 349.200 250.300 ;
        RECT 345.200 247.600 346.000 248.400 ;
        RECT 337.200 231.600 338.000 232.400 ;
        RECT 338.800 232.300 339.600 232.400 ;
        RECT 338.800 231.700 341.100 232.300 ;
        RECT 338.800 231.600 339.600 231.700 ;
        RECT 337.300 230.400 337.900 231.600 ;
        RECT 338.900 230.400 339.500 231.600 ;
        RECT 337.200 229.600 338.000 230.400 ;
        RECT 338.800 229.600 339.600 230.400 ;
        RECT 332.400 227.600 333.200 228.400 ;
        RECT 334.000 227.600 334.800 228.400 ;
        RECT 337.200 227.600 338.000 228.400 ;
        RECT 334.000 215.600 334.800 216.400 ;
        RECT 332.400 213.600 333.200 214.400 ;
        RECT 330.800 211.600 331.600 212.400 ;
        RECT 319.600 185.600 320.400 186.400 ;
        RECT 321.200 184.200 322.000 195.800 ;
        RECT 322.800 187.600 323.600 188.400 ;
        RECT 297.200 181.600 298.000 182.400 ;
        RECT 303.700 176.400 304.300 183.600 ;
        RECT 322.900 178.400 323.500 187.600 ;
        RECT 324.400 184.200 325.200 195.800 ;
        RECT 326.000 184.200 326.800 197.800 ;
        RECT 327.600 184.200 328.400 197.800 ;
        RECT 334.100 196.400 334.700 215.600 ;
        RECT 335.600 211.600 336.400 212.400 ;
        RECT 335.700 210.400 336.300 211.600 ;
        RECT 335.600 209.600 336.400 210.400 ;
        RECT 334.000 195.600 334.800 196.400 ;
        RECT 332.400 191.600 333.200 192.400 ;
        RECT 332.500 182.400 333.100 191.600 ;
        RECT 335.700 186.400 336.300 209.600 ;
        RECT 337.200 193.600 338.000 194.400 ;
        RECT 337.300 190.400 337.900 193.600 ;
        RECT 337.200 189.600 338.000 190.400 ;
        RECT 337.300 186.400 337.900 189.600 ;
        RECT 335.600 185.600 336.400 186.400 ;
        RECT 337.200 185.600 338.000 186.400 ;
        RECT 338.800 185.600 339.600 186.400 ;
        RECT 324.400 181.600 325.200 182.400 ;
        RECT 332.400 181.600 333.200 182.400 ;
        RECT 303.600 175.600 304.400 176.400 ;
        RECT 303.700 152.400 304.300 175.600 ;
        RECT 305.200 164.200 306.000 177.800 ;
        RECT 306.800 164.200 307.600 177.800 ;
        RECT 308.400 164.200 309.200 177.800 ;
        RECT 310.000 166.200 310.800 177.800 ;
        RECT 311.600 175.600 312.400 176.400 ;
        RECT 311.700 164.400 312.300 175.600 ;
        RECT 313.200 166.200 314.000 177.800 ;
        RECT 314.800 177.600 315.600 178.400 ;
        RECT 314.900 174.400 315.500 177.600 ;
        RECT 314.800 173.600 315.600 174.400 ;
        RECT 316.400 166.200 317.200 177.800 ;
        RECT 311.600 163.600 312.400 164.400 ;
        RECT 318.000 164.200 318.800 177.800 ;
        RECT 319.600 164.200 320.400 177.800 ;
        RECT 322.800 177.600 323.600 178.400 ;
        RECT 324.500 172.400 325.100 181.600 ;
        RECT 332.400 179.600 333.200 180.400 ;
        RECT 332.500 174.400 333.100 179.600 ;
        RECT 334.000 175.600 334.800 176.400 ;
        RECT 332.400 173.600 333.200 174.400 ;
        RECT 321.200 171.600 322.000 172.400 ;
        RECT 324.400 171.600 325.200 172.400 ;
        RECT 303.600 151.600 304.400 152.400 ;
        RECT 281.200 149.600 282.000 150.400 ;
        RECT 290.800 149.600 291.600 150.400 ;
        RECT 295.400 149.600 296.400 150.400 ;
        RECT 265.200 147.600 266.000 148.400 ;
        RECT 266.800 147.600 267.600 148.400 ;
        RECT 279.600 147.600 280.400 148.400 ;
        RECT 281.300 148.300 281.900 149.600 ;
        RECT 282.800 148.300 283.600 148.800 ;
        RECT 281.300 148.000 283.600 148.300 ;
        RECT 281.300 147.700 283.500 148.000 ;
        RECT 287.600 147.600 288.400 148.400 ;
        RECT 262.000 145.600 262.800 146.400 ;
        RECT 263.600 145.600 264.400 146.400 ;
        RECT 265.300 138.400 265.900 147.600 ;
        RECT 266.800 145.600 267.600 146.400 ;
        RECT 265.200 137.600 266.000 138.400 ;
        RECT 260.400 133.600 261.200 134.400 ;
        RECT 257.200 131.600 258.000 132.400 ;
        RECT 260.400 131.600 261.200 132.400 ;
        RECT 263.600 131.600 264.400 132.400 ;
        RECT 250.800 109.600 251.600 110.400 ;
        RECT 252.400 109.600 253.200 110.400 ;
        RECT 255.600 109.600 256.400 110.400 ;
        RECT 250.900 108.400 251.500 109.600 ;
        RECT 252.500 108.400 253.100 109.600 ;
        RECT 242.800 107.600 243.600 108.400 ;
        RECT 246.000 107.600 246.800 108.400 ;
        RECT 249.200 107.600 250.000 108.400 ;
        RECT 250.800 107.600 251.600 108.400 ;
        RECT 252.400 107.600 253.200 108.400 ;
        RECT 254.000 107.600 254.800 108.400 ;
        RECT 236.400 105.600 237.200 106.400 ;
        RECT 239.600 105.600 240.400 106.400 ;
        RECT 241.200 105.600 242.000 106.400 ;
        RECT 234.800 101.600 235.600 102.400 ;
        RECT 212.400 95.600 213.200 96.400 ;
        RECT 218.800 95.600 219.600 96.400 ;
        RECT 222.000 95.600 222.800 96.400 ;
        RECT 226.800 95.600 227.600 96.400 ;
        RECT 228.400 95.600 229.200 96.400 ;
        RECT 231.600 95.600 232.400 96.400 ;
        RECT 234.800 95.600 235.600 96.400 ;
        RECT 212.500 94.400 213.100 95.600 ;
        RECT 218.900 94.400 219.500 95.600 ;
        RECT 212.400 93.600 213.200 94.400 ;
        RECT 218.800 93.600 219.600 94.400 ;
        RECT 222.100 92.400 222.700 95.600 ;
        RECT 228.500 94.400 229.100 95.600 ;
        RECT 234.900 94.400 235.500 95.600 ;
        RECT 223.600 93.600 224.400 94.400 ;
        RECT 225.200 93.600 226.000 94.400 ;
        RECT 228.400 93.600 229.200 94.400 ;
        RECT 231.600 93.600 232.400 94.400 ;
        RECT 234.800 93.600 235.600 94.400 ;
        RECT 236.400 93.600 237.200 94.400 ;
        RECT 238.000 93.600 238.800 94.400 ;
        RECT 222.000 91.600 222.800 92.400 ;
        RECT 225.300 92.300 225.900 93.600 ;
        RECT 236.500 92.400 237.100 93.600 ;
        RECT 223.700 91.700 225.900 92.300 ;
        RECT 222.100 90.400 222.700 91.600 ;
        RECT 212.400 89.600 213.200 90.400 ;
        RECT 222.000 89.600 222.800 90.400 ;
        RECT 223.700 88.400 224.300 91.700 ;
        RECT 236.400 91.600 237.200 92.400 ;
        RECT 226.800 89.600 227.600 90.400 ;
        RECT 238.100 88.400 238.700 93.600 ;
        RECT 241.300 92.400 241.900 105.600 ;
        RECT 242.900 96.400 243.500 107.600 ;
        RECT 244.400 105.600 245.200 106.400 ;
        RECT 242.800 95.600 243.600 96.400 ;
        RECT 241.200 91.600 242.000 92.400 ;
        RECT 242.900 90.400 243.500 95.600 ;
        RECT 244.500 94.400 245.100 105.600 ;
        RECT 254.100 104.400 254.700 107.600 ;
        RECT 257.300 106.400 257.900 131.600 ;
        RECT 260.500 130.400 261.100 131.600 ;
        RECT 263.700 130.400 264.300 131.600 ;
        RECT 260.400 129.600 261.200 130.400 ;
        RECT 263.600 129.600 264.400 130.400 ;
        RECT 266.900 120.400 267.500 145.600 ;
        RECT 305.200 144.200 306.000 157.800 ;
        RECT 306.800 144.200 307.600 157.800 ;
        RECT 308.400 144.200 309.200 157.800 ;
        RECT 310.000 144.200 310.800 155.800 ;
        RECT 311.600 145.600 312.400 146.400 ;
        RECT 310.000 141.600 310.800 142.400 ;
        RECT 273.200 135.600 274.000 136.400 ;
        RECT 274.800 127.600 275.600 128.400 ;
        RECT 266.800 119.600 267.600 120.400 ;
        RECT 258.800 111.600 259.600 112.400 ;
        RECT 258.900 110.400 259.500 111.600 ;
        RECT 258.800 109.600 259.600 110.400 ;
        RECT 257.200 105.600 258.000 106.400 ;
        RECT 247.600 103.600 248.400 104.400 ;
        RECT 254.000 103.600 254.800 104.400 ;
        RECT 246.000 99.600 246.800 100.400 ;
        RECT 244.400 93.600 245.200 94.400 ;
        RECT 246.100 92.400 246.700 99.600 ;
        RECT 247.700 94.300 248.300 103.600 ;
        RECT 250.800 101.600 251.600 102.400 ;
        RECT 250.900 98.400 251.500 101.600 ;
        RECT 258.900 98.400 259.500 109.600 ;
        RECT 262.000 107.600 262.800 108.400 ;
        RECT 262.100 100.400 262.700 107.600 ;
        RECT 266.900 106.400 267.500 119.600 ;
        RECT 274.900 110.400 275.500 127.600 ;
        RECT 282.800 124.200 283.600 137.800 ;
        RECT 284.400 124.200 285.200 137.800 ;
        RECT 286.000 124.200 286.800 137.800 ;
        RECT 287.600 126.200 288.400 137.800 ;
        RECT 289.200 135.600 290.000 136.400 ;
        RECT 289.300 124.300 289.900 135.600 ;
        RECT 290.800 126.200 291.600 137.800 ;
        RECT 292.400 133.600 293.200 134.400 ;
        RECT 294.000 126.200 294.800 137.800 ;
        RECT 289.300 123.700 291.500 124.300 ;
        RECT 295.600 124.200 296.400 137.800 ;
        RECT 297.200 124.200 298.000 137.800 ;
        RECT 306.800 133.600 307.600 134.400 ;
        RECT 310.100 132.400 310.700 141.600 ;
        RECT 310.000 131.600 310.800 132.400 ;
        RECT 303.600 129.600 304.400 130.400 ;
        RECT 306.800 129.600 307.600 130.400 ;
        RECT 274.600 109.600 275.600 110.400 ;
        RECT 266.800 105.600 267.600 106.400 ;
        RECT 263.600 103.600 264.400 104.400 ;
        RECT 284.400 104.200 285.200 117.800 ;
        RECT 286.000 104.200 286.800 117.800 ;
        RECT 287.600 104.200 288.400 117.800 ;
        RECT 289.200 104.200 290.000 115.800 ;
        RECT 290.900 106.400 291.500 123.700 ;
        RECT 290.800 105.600 291.600 106.400 ;
        RECT 262.000 99.600 262.800 100.400 ;
        RECT 250.800 97.600 251.600 98.400 ;
        RECT 258.800 97.600 259.600 98.400 ;
        RECT 262.000 97.600 262.800 98.400 ;
        RECT 249.200 95.600 250.000 96.400 ;
        RECT 260.400 95.600 261.200 96.400 ;
        RECT 247.700 93.700 249.900 94.300 ;
        RECT 246.000 91.600 246.800 92.400 ;
        RECT 247.600 91.600 248.400 92.400 ;
        RECT 242.800 89.600 243.600 90.400 ;
        RECT 223.600 87.600 224.400 88.400 ;
        RECT 238.000 87.600 238.800 88.400 ;
        RECT 231.600 83.600 232.400 84.400 ;
        RECT 231.700 80.400 232.300 83.600 ;
        RECT 228.400 79.600 229.200 80.400 ;
        RECT 231.600 79.600 232.400 80.400 ;
        RECT 210.800 69.600 211.600 70.400 ;
        RECT 217.200 69.600 218.000 70.400 ;
        RECT 198.000 65.600 198.800 66.400 ;
        RECT 218.800 64.200 219.600 77.800 ;
        RECT 220.400 64.200 221.200 77.800 ;
        RECT 222.000 64.200 222.800 77.800 ;
        RECT 223.600 64.200 224.400 75.800 ;
        RECT 225.200 65.600 226.000 66.400 ;
        RECT 226.800 64.200 227.600 75.800 ;
        RECT 228.500 68.400 229.100 79.600 ;
        RECT 228.400 67.600 229.200 68.400 ;
        RECT 230.000 64.200 230.800 75.800 ;
        RECT 231.600 64.200 232.400 77.800 ;
        RECT 233.200 64.200 234.000 77.800 ;
        RECT 247.600 73.600 248.400 74.400 ;
        RECT 239.600 69.600 240.400 70.400 ;
        RECT 214.000 59.600 214.800 60.400 ;
        RECT 218.800 59.600 219.600 60.400 ;
        RECT 230.000 59.600 230.800 60.400 ;
        RECT 180.400 49.600 181.200 50.400 ;
        RECT 180.500 40.400 181.100 49.600 ;
        RECT 185.200 44.200 186.000 57.800 ;
        RECT 186.800 44.200 187.600 57.800 ;
        RECT 188.400 46.200 189.200 57.800 ;
        RECT 190.000 53.600 190.800 54.400 ;
        RECT 190.100 52.400 190.700 53.600 ;
        RECT 190.000 51.600 190.800 52.400 ;
        RECT 191.600 46.200 192.400 57.800 ;
        RECT 193.200 55.600 194.000 56.400 ;
        RECT 193.300 42.400 193.900 55.600 ;
        RECT 194.800 46.200 195.600 57.800 ;
        RECT 196.400 44.200 197.200 57.800 ;
        RECT 198.000 44.200 198.800 57.800 ;
        RECT 199.600 44.200 200.400 57.800 ;
        RECT 202.800 53.600 203.600 54.400 ;
        RECT 212.400 53.600 213.200 54.400 ;
        RECT 185.200 41.600 186.000 42.400 ;
        RECT 193.200 41.600 194.000 42.400 ;
        RECT 178.800 39.600 179.600 40.400 ;
        RECT 180.400 39.600 181.200 40.400 ;
        RECT 169.200 37.600 170.000 38.400 ;
        RECT 178.800 24.200 179.600 37.800 ;
        RECT 180.400 24.200 181.200 37.800 ;
        RECT 182.000 24.200 182.800 37.800 ;
        RECT 183.600 24.200 184.400 35.800 ;
        RECT 185.300 26.400 185.900 41.600 ;
        RECT 194.800 39.600 195.600 40.400 ;
        RECT 185.200 25.600 186.000 26.400 ;
        RECT 185.300 22.400 185.900 25.600 ;
        RECT 186.800 24.200 187.600 35.800 ;
        RECT 188.400 27.600 189.200 28.400 ;
        RECT 190.000 24.200 190.800 35.800 ;
        RECT 191.600 24.200 192.400 37.800 ;
        RECT 193.200 24.200 194.000 37.800 ;
        RECT 194.900 32.000 195.500 39.600 ;
        RECT 194.800 31.200 195.600 32.000 ;
        RECT 202.900 28.400 203.500 53.600 ;
        RECT 212.500 50.300 213.100 53.600 ;
        RECT 214.100 52.400 214.700 59.600 ;
        RECT 214.000 51.600 214.800 52.400 ;
        RECT 215.600 51.600 216.400 52.400 ;
        RECT 218.900 50.400 219.500 59.600 ;
        RECT 226.800 55.600 227.600 56.400 ;
        RECT 223.600 53.600 224.400 54.400 ;
        RECT 222.000 51.600 222.800 52.400 ;
        RECT 212.500 49.700 214.700 50.300 ;
        RECT 210.800 47.600 211.600 48.400 ;
        RECT 207.600 31.600 208.400 32.400 ;
        RECT 210.900 30.400 211.500 47.600 ;
        RECT 214.100 34.400 214.700 49.700 ;
        RECT 218.800 49.600 219.600 50.400 ;
        RECT 214.000 33.600 214.800 34.400 ;
        RECT 218.800 31.600 219.600 32.400 ;
        RECT 222.000 31.600 222.800 32.400 ;
        RECT 210.800 29.600 211.600 30.400 ;
        RECT 212.400 29.600 213.200 30.400 ;
        RECT 214.000 29.600 214.800 30.400 ;
        RECT 222.000 29.600 222.800 30.400 ;
        RECT 212.500 28.400 213.100 29.600 ;
        RECT 202.800 27.600 203.600 28.400 ;
        RECT 204.400 27.600 205.200 28.400 ;
        RECT 212.400 27.600 213.200 28.400 ;
        RECT 202.900 22.400 203.500 27.600 ;
        RECT 212.500 24.300 213.100 27.600 ;
        RECT 214.100 26.400 214.700 29.600 ;
        RECT 223.700 28.400 224.300 53.600 ;
        RECT 226.900 52.400 227.500 55.600 ;
        RECT 230.100 52.400 230.700 59.600 ;
        RECT 234.800 55.600 235.600 56.400 ;
        RECT 226.800 51.600 227.600 52.400 ;
        RECT 230.000 51.600 230.800 52.400 ;
        RECT 236.200 51.600 237.200 52.400 ;
        RECT 225.200 49.600 226.000 50.400 ;
        RECT 225.300 38.400 225.900 49.600 ;
        RECT 226.800 47.600 227.600 48.400 ;
        RECT 225.200 37.600 226.000 38.400 ;
        RECT 226.900 32.400 227.500 47.600 ;
        RECT 230.100 32.400 230.700 51.600 ;
        RECT 239.700 50.400 240.300 69.600 ;
        RECT 247.700 66.400 248.300 73.600 ;
        RECT 242.800 65.600 243.600 66.400 ;
        RECT 247.600 65.600 248.400 66.400 ;
        RECT 242.900 58.400 243.500 65.600 ;
        RECT 249.300 60.400 249.900 93.700 ;
        RECT 257.200 91.600 258.000 92.400 ;
        RECT 252.400 71.600 253.200 72.400 ;
        RECT 257.200 71.600 258.000 72.400 ;
        RECT 252.500 70.400 253.100 71.600 ;
        RECT 252.400 69.600 253.200 70.400 ;
        RECT 262.100 68.400 262.700 97.600 ;
        RECT 263.700 94.400 264.300 103.600 ;
        RECT 290.900 100.400 291.500 105.600 ;
        RECT 292.400 104.200 293.200 115.800 ;
        RECT 294.000 107.600 294.800 108.400 ;
        RECT 295.600 104.200 296.400 115.800 ;
        RECT 297.200 104.200 298.000 117.800 ;
        RECT 298.800 104.200 299.600 117.800 ;
        RECT 303.700 112.400 304.300 129.600 ;
        RECT 300.400 111.200 301.200 112.000 ;
        RECT 303.600 111.600 304.400 112.400 ;
        RECT 286.000 99.600 286.800 100.400 ;
        RECT 290.800 99.600 291.600 100.400 ;
        RECT 263.600 93.600 264.400 94.400 ;
        RECT 278.000 91.600 278.800 92.400 ;
        RECT 263.600 85.600 264.400 86.400 ;
        RECT 262.000 67.600 262.800 68.400 ;
        RECT 262.100 66.400 262.700 67.600 ;
        RECT 263.700 66.400 264.300 85.600 ;
        RECT 273.200 69.600 274.000 70.400 ;
        RECT 278.100 70.300 278.700 91.600 ;
        RECT 279.600 84.200 280.400 97.800 ;
        RECT 281.200 84.200 282.000 97.800 ;
        RECT 282.800 84.200 283.600 97.800 ;
        RECT 284.400 86.200 285.200 97.800 ;
        RECT 286.100 96.400 286.700 99.600 ;
        RECT 286.000 95.600 286.800 96.400 ;
        RECT 286.100 80.400 286.700 95.600 ;
        RECT 287.600 86.200 288.400 97.800 ;
        RECT 289.200 93.600 290.000 94.400 ;
        RECT 290.800 86.200 291.600 97.800 ;
        RECT 292.400 84.200 293.200 97.800 ;
        RECT 294.000 84.200 294.800 97.800 ;
        RECT 300.500 92.400 301.100 111.200 ;
        RECT 308.400 107.600 309.200 108.400 ;
        RECT 303.600 103.600 304.400 104.400 ;
        RECT 303.700 96.400 304.300 103.600 ;
        RECT 308.500 98.400 309.100 107.600 ;
        RECT 311.700 106.400 312.300 145.600 ;
        RECT 313.200 144.200 314.000 155.800 ;
        RECT 314.800 147.600 315.600 148.400 ;
        RECT 316.400 144.200 317.200 155.800 ;
        RECT 318.000 144.200 318.800 157.800 ;
        RECT 319.600 144.200 320.400 157.800 ;
        RECT 321.300 152.000 321.900 171.600 ;
        RECT 329.200 169.600 330.000 170.400 ;
        RECT 330.800 163.600 331.600 164.400 ;
        RECT 321.200 151.200 322.000 152.000 ;
        RECT 326.000 151.600 326.800 152.400 ;
        RECT 329.200 151.600 330.000 152.400 ;
        RECT 321.200 143.600 322.000 144.400 ;
        RECT 318.000 139.600 318.800 140.400 ;
        RECT 314.800 135.600 315.600 136.400 ;
        RECT 316.400 133.600 317.200 134.400 ;
        RECT 314.800 131.600 315.600 132.400 ;
        RECT 314.900 130.400 315.500 131.600 ;
        RECT 316.500 130.400 317.100 133.600 ;
        RECT 314.800 129.600 315.600 130.400 ;
        RECT 316.400 129.600 317.200 130.400 ;
        RECT 313.200 111.600 314.000 112.400 ;
        RECT 311.600 105.600 312.400 106.400 ;
        RECT 313.200 103.600 314.000 104.400 ;
        RECT 308.400 97.600 309.200 98.400 ;
        RECT 303.600 95.600 304.400 96.400 ;
        RECT 306.800 95.600 307.600 96.400 ;
        RECT 300.400 91.600 301.200 92.400 ;
        RECT 305.200 83.600 306.000 84.400 ;
        RECT 286.000 79.600 286.800 80.400 ;
        RECT 290.800 79.600 291.600 80.400 ;
        RECT 278.100 69.700 280.300 70.300 ;
        RECT 262.000 65.600 262.800 66.400 ;
        RECT 263.600 65.600 264.400 66.400 ;
        RECT 266.800 65.600 267.600 66.400 ;
        RECT 255.600 63.600 256.400 64.400 ;
        RECT 249.200 59.600 250.000 60.400 ;
        RECT 242.800 57.600 243.600 58.400 ;
        RECT 233.200 49.600 234.000 50.400 ;
        RECT 239.600 49.600 240.400 50.400 ;
        RECT 246.000 44.200 246.800 57.800 ;
        RECT 247.600 44.200 248.400 57.800 ;
        RECT 249.200 44.200 250.000 57.800 ;
        RECT 250.800 46.200 251.600 57.800 ;
        RECT 252.400 55.600 253.200 56.400 ;
        RECT 252.500 42.400 253.100 55.600 ;
        RECT 254.000 46.200 254.800 57.800 ;
        RECT 255.600 55.600 256.400 56.400 ;
        RECT 255.700 54.400 256.300 55.600 ;
        RECT 255.600 53.600 256.400 54.400 ;
        RECT 257.200 46.200 258.000 57.800 ;
        RECT 258.800 44.200 259.600 57.800 ;
        RECT 260.400 44.200 261.200 57.800 ;
        RECT 262.000 49.600 262.800 50.800 ;
        RECT 279.700 50.400 280.300 69.700 ;
        RECT 284.400 64.200 285.200 77.800 ;
        RECT 286.000 64.200 286.800 77.800 ;
        RECT 287.600 64.200 288.400 77.800 ;
        RECT 289.200 64.200 290.000 75.800 ;
        RECT 290.900 66.400 291.500 79.600 ;
        RECT 290.800 65.600 291.600 66.400 ;
        RECT 290.900 60.400 291.500 65.600 ;
        RECT 292.400 64.200 293.200 75.800 ;
        RECT 294.000 67.600 294.800 68.400 ;
        RECT 294.100 66.400 294.700 67.600 ;
        RECT 294.000 65.600 294.800 66.400 ;
        RECT 294.000 63.600 294.800 64.400 ;
        RECT 295.600 64.200 296.400 75.800 ;
        RECT 297.200 64.200 298.000 77.800 ;
        RECT 298.800 64.200 299.600 77.800 ;
        RECT 305.300 76.400 305.900 83.600 ;
        RECT 308.400 79.600 309.200 80.400 ;
        RECT 305.200 75.600 306.000 76.400 ;
        RECT 303.600 71.600 304.400 72.400 ;
        RECT 303.700 64.400 304.300 71.600 ;
        RECT 308.500 70.400 309.100 79.600 ;
        RECT 313.300 74.400 313.900 103.600 ;
        RECT 314.900 92.400 315.500 129.600 ;
        RECT 318.100 112.400 318.700 139.600 ;
        RECT 321.300 134.400 321.900 143.600 ;
        RECT 321.200 133.600 322.000 134.400 ;
        RECT 326.100 132.400 326.700 151.600 ;
        RECT 329.200 147.600 330.000 148.400 ;
        RECT 330.900 146.400 331.500 163.600 ;
        RECT 334.100 154.400 334.700 175.600 ;
        RECT 338.900 172.400 339.500 185.600 ;
        RECT 338.800 171.600 339.600 172.400 ;
        RECT 340.500 170.300 341.100 231.700 ;
        RECT 343.600 227.600 344.400 228.400 ;
        RECT 345.300 218.400 345.900 247.600 ;
        RECT 342.000 217.600 342.800 218.400 ;
        RECT 343.600 217.600 344.400 218.400 ;
        RECT 345.200 217.600 346.000 218.400 ;
        RECT 342.100 216.400 342.700 217.600 ;
        RECT 342.000 215.600 342.800 216.400 ;
        RECT 342.000 213.600 342.800 214.400 ;
        RECT 342.100 200.400 342.700 213.600 ;
        RECT 346.900 210.400 347.500 249.700 ;
        RECT 348.400 249.600 349.200 249.700 ;
        RECT 354.800 249.600 355.600 250.400 ;
        RECT 358.000 244.200 358.800 257.800 ;
        RECT 359.600 244.200 360.400 257.800 ;
        RECT 361.200 246.200 362.000 257.800 ;
        RECT 362.800 255.600 363.600 256.400 ;
        RECT 362.900 254.400 363.500 255.600 ;
        RECT 362.800 253.600 363.600 254.400 ;
        RECT 362.800 251.600 363.600 252.400 ;
        RECT 362.900 244.300 363.500 251.600 ;
        RECT 364.400 246.200 365.200 257.800 ;
        RECT 366.000 255.600 366.800 256.400 ;
        RECT 361.300 243.700 363.500 244.300 ;
        RECT 356.400 241.600 357.200 242.400 ;
        RECT 356.500 238.400 357.100 241.600 ;
        RECT 361.300 238.400 361.900 243.700 ;
        RECT 356.400 237.600 357.200 238.400 ;
        RECT 361.200 237.600 362.000 238.400 ;
        RECT 366.100 236.400 366.700 255.600 ;
        RECT 367.600 246.200 368.400 257.800 ;
        RECT 369.200 244.200 370.000 257.800 ;
        RECT 370.800 244.200 371.600 257.800 ;
        RECT 372.400 244.200 373.200 257.800 ;
        RECT 351.600 235.600 352.400 236.400 ;
        RECT 361.200 235.600 362.000 236.400 ;
        RECT 366.000 235.600 366.800 236.400 ;
        RECT 346.800 209.600 347.600 210.400 ;
        RECT 350.000 206.200 350.800 217.800 ;
        RECT 342.000 199.600 342.800 200.400 ;
        RECT 348.400 199.600 349.200 200.400 ;
        RECT 345.200 192.300 346.000 192.400 ;
        RECT 345.200 191.700 347.500 192.300 ;
        RECT 345.200 191.600 346.000 191.700 ;
        RECT 342.000 189.600 342.800 190.400 ;
        RECT 342.100 186.400 342.700 189.600 ;
        RECT 345.200 187.600 346.000 188.400 ;
        RECT 342.000 185.600 342.800 186.400 ;
        RECT 343.600 185.600 344.400 186.400 ;
        RECT 342.000 177.600 342.800 178.400 ;
        RECT 343.700 170.400 344.300 185.600 ;
        RECT 338.900 169.700 341.100 170.300 ;
        RECT 337.200 155.600 338.000 156.400 ;
        RECT 334.000 153.600 334.800 154.400 ;
        RECT 337.300 150.400 337.900 155.600 ;
        RECT 338.900 152.400 339.500 169.700 ;
        RECT 343.600 169.600 344.400 170.400 ;
        RECT 338.800 151.600 339.600 152.400 ;
        RECT 340.400 151.600 341.200 152.400 ;
        RECT 343.700 152.300 344.300 169.600 ;
        RECT 345.200 152.300 346.000 152.400 ;
        RECT 343.700 151.700 346.000 152.300 ;
        RECT 345.200 151.600 346.000 151.700 ;
        RECT 332.400 149.600 333.200 150.400 ;
        RECT 337.200 149.600 338.000 150.400 ;
        RECT 330.800 145.600 331.600 146.400 ;
        RECT 332.500 142.400 333.100 149.600 ;
        RECT 337.300 146.400 337.900 149.600 ;
        RECT 337.200 145.600 338.000 146.400 ;
        RECT 338.900 142.400 339.500 151.600 ;
        RECT 340.500 150.400 341.100 151.600 ;
        RECT 340.400 149.600 341.200 150.400 ;
        RECT 343.600 149.600 344.400 150.400 ;
        RECT 343.700 148.400 344.300 149.600 ;
        RECT 343.600 147.600 344.400 148.400 ;
        RECT 343.700 144.400 344.300 147.600 ;
        RECT 343.600 143.600 344.400 144.400 ;
        RECT 332.400 141.600 333.200 142.400 ;
        RECT 338.800 141.600 339.600 142.400 ;
        RECT 345.300 140.400 345.900 151.600 ;
        RECT 346.900 150.400 347.500 191.700 ;
        RECT 348.500 176.400 349.100 199.600 ;
        RECT 348.400 175.600 349.200 176.400 ;
        RECT 348.500 174.400 349.100 175.600 ;
        RECT 348.400 173.600 349.200 174.400 ;
        RECT 351.700 158.400 352.300 235.600 ;
        RECT 359.600 231.600 360.400 232.400 ;
        RECT 356.400 229.600 357.200 230.400 ;
        RECT 353.200 227.600 354.000 228.400 ;
        RECT 354.800 227.600 355.600 228.400 ;
        RECT 354.900 218.400 355.500 227.600 ;
        RECT 354.800 217.600 355.600 218.400 ;
        RECT 358.000 211.800 358.800 212.600 ;
        RECT 358.100 210.400 358.700 211.800 ;
        RECT 358.000 209.600 358.800 210.400 ;
        RECT 359.600 206.200 360.400 217.800 ;
        RECT 361.300 214.400 361.900 235.600 ;
        RECT 375.700 232.400 376.300 259.600 ;
        RECT 378.900 238.400 379.500 297.600 ;
        RECT 383.700 296.400 384.300 297.600 ;
        RECT 383.600 295.600 384.400 296.400 ;
        RECT 382.000 293.600 382.800 294.400 ;
        RECT 391.600 293.600 392.400 294.400 ;
        RECT 393.200 293.600 394.000 294.400 ;
        RECT 394.800 293.600 395.600 294.400 ;
        RECT 380.400 291.600 381.200 292.400 ;
        RECT 380.500 286.400 381.100 291.600 ;
        RECT 382.100 288.400 382.700 293.600 ;
        RECT 383.600 291.600 384.400 292.400 ;
        RECT 388.400 289.600 389.200 290.400 ;
        RECT 391.700 288.400 392.300 293.600 ;
        RECT 382.000 287.600 382.800 288.400 ;
        RECT 391.600 287.600 392.400 288.400 ;
        RECT 393.300 286.400 393.900 293.600 ;
        RECT 394.900 292.400 395.500 293.600 ;
        RECT 394.800 291.600 395.600 292.400 ;
        RECT 396.400 291.600 397.200 292.400 ;
        RECT 398.100 290.400 398.700 297.600 ;
        RECT 409.300 296.400 409.900 299.600 ;
        RECT 410.900 298.400 411.500 311.700 ;
        RECT 412.500 308.400 413.100 323.600 ;
        RECT 414.100 310.400 414.700 331.600 ;
        RECT 414.000 309.600 414.800 310.400 ;
        RECT 412.400 307.600 413.200 308.400 ;
        RECT 417.300 306.400 417.900 333.600 ;
        RECT 418.900 306.400 419.500 335.600 ;
        RECT 428.500 326.400 429.100 337.600 ;
        RECT 434.900 332.400 435.500 351.600 ;
        RECT 436.400 349.600 437.200 350.400 ;
        RECT 442.800 349.600 443.600 350.400 ;
        RECT 449.200 349.600 450.000 350.400 ;
        RECT 436.400 347.600 437.200 348.400 ;
        RECT 447.600 347.600 448.400 348.400 ;
        RECT 436.500 338.400 437.100 347.600 ;
        RECT 442.800 345.600 443.600 346.400 ;
        RECT 439.600 343.600 440.400 344.400 ;
        RECT 436.400 337.600 437.200 338.400 ;
        RECT 439.700 332.400 440.300 343.600 ;
        RECT 430.000 332.300 430.800 332.400 ;
        RECT 430.000 331.700 432.300 332.300 ;
        RECT 430.000 331.600 430.800 331.700 ;
        RECT 428.400 325.600 429.200 326.400 ;
        RECT 430.000 311.600 430.800 312.400 ;
        RECT 430.100 310.400 430.700 311.600 ;
        RECT 430.000 309.600 430.800 310.400 ;
        RECT 414.000 305.600 414.800 306.400 ;
        RECT 417.200 305.600 418.000 306.400 ;
        RECT 418.800 305.600 419.600 306.400 ;
        RECT 428.400 305.600 429.200 306.400 ;
        RECT 430.000 305.600 430.800 306.400 ;
        RECT 410.800 297.600 411.600 298.400 ;
        RECT 409.200 295.600 410.000 296.400 ;
        RECT 399.600 293.600 400.400 294.400 ;
        RECT 402.800 293.600 403.600 294.400 ;
        RECT 398.000 289.600 398.800 290.400 ;
        RECT 399.600 289.600 400.400 290.400 ;
        RECT 402.900 288.400 403.500 293.600 ;
        RECT 407.600 289.600 408.400 290.400 ;
        RECT 402.800 287.600 403.600 288.400 ;
        RECT 380.400 285.600 381.200 286.400 ;
        RECT 388.400 285.600 389.200 286.400 ;
        RECT 393.200 285.600 394.000 286.400 ;
        RECT 386.800 269.600 387.600 270.400 ;
        RECT 380.400 263.600 381.200 264.400 ;
        RECT 380.500 258.400 381.100 263.600 ;
        RECT 380.400 257.600 381.200 258.400 ;
        RECT 383.600 247.600 384.400 248.400 ;
        RECT 378.800 237.600 379.600 238.400 ;
        RECT 366.000 231.600 366.800 232.400 ;
        RECT 367.600 231.600 368.400 232.400 ;
        RECT 370.800 231.600 371.600 232.400 ;
        RECT 375.600 231.600 376.400 232.400 ;
        RECT 366.100 230.400 366.700 231.600 ;
        RECT 367.700 230.400 368.300 231.600 ;
        RECT 366.000 229.600 366.800 230.400 ;
        RECT 367.600 229.600 368.400 230.400 ;
        RECT 361.200 213.600 362.000 214.400 ;
        RECT 361.300 198.300 361.900 213.600 ;
        RECT 362.800 210.200 363.600 215.800 ;
        RECT 366.100 214.400 366.700 229.600 ;
        RECT 370.900 228.400 371.500 231.600 ;
        RECT 370.800 227.600 371.600 228.400 ;
        RECT 374.000 223.600 374.800 224.400 ;
        RECT 370.800 217.600 371.600 218.400 ;
        RECT 370.900 214.400 371.500 217.600 ;
        RECT 374.100 214.400 374.700 223.600 ;
        RECT 366.000 213.600 366.800 214.400 ;
        RECT 369.200 213.600 370.000 214.400 ;
        RECT 370.800 213.600 371.600 214.400 ;
        RECT 374.000 213.600 374.800 214.400 ;
        RECT 367.600 211.600 368.400 212.400 ;
        RECT 364.400 209.600 365.200 210.400 ;
        RECT 364.500 208.400 365.100 209.600 ;
        RECT 364.400 207.600 365.200 208.400 ;
        RECT 369.300 204.400 369.900 213.600 ;
        RECT 372.400 211.600 373.200 212.400 ;
        RECT 375.700 208.400 376.300 231.600 ;
        RECT 377.200 229.600 378.000 230.400 ;
        RECT 378.800 225.600 379.600 226.400 ;
        RECT 378.800 223.600 379.600 224.400 ;
        RECT 378.900 216.400 379.500 223.600 ;
        RECT 378.800 215.600 379.600 216.400 ;
        RECT 378.800 213.600 379.600 214.400 ;
        RECT 380.400 213.600 381.200 214.400 ;
        RECT 382.000 213.600 382.800 214.400 ;
        RECT 377.200 211.600 378.000 212.400 ;
        RECT 370.800 207.600 371.600 208.400 ;
        RECT 375.600 207.600 376.400 208.400 ;
        RECT 369.200 203.600 370.000 204.400 ;
        RECT 353.200 191.200 354.000 192.000 ;
        RECT 353.300 182.400 353.900 191.200 ;
        RECT 354.800 184.200 355.600 197.800 ;
        RECT 356.400 184.200 357.200 197.800 ;
        RECT 361.300 197.700 363.500 198.300 ;
        RECT 358.000 184.200 358.800 195.800 ;
        RECT 359.600 187.600 360.400 188.400 ;
        RECT 359.600 185.600 360.400 186.400 ;
        RECT 353.200 181.600 354.000 182.400 ;
        RECT 354.800 177.600 355.600 178.400 ;
        RECT 353.200 175.600 354.000 176.400 ;
        RECT 353.200 163.600 354.000 164.400 ;
        RECT 351.600 157.600 352.400 158.400 ;
        RECT 351.600 151.600 352.400 152.400 ;
        RECT 353.300 150.400 353.900 163.600 ;
        RECT 354.900 158.400 355.500 177.600 ;
        RECT 356.400 175.600 357.200 176.400 ;
        RECT 356.500 174.400 357.100 175.600 ;
        RECT 356.400 173.600 357.200 174.400 ;
        RECT 356.500 160.400 357.100 173.600 ;
        RECT 359.700 172.400 360.300 185.600 ;
        RECT 361.200 184.200 362.000 195.800 ;
        RECT 362.900 186.400 363.500 197.700 ;
        RECT 362.800 185.600 363.600 186.400 ;
        RECT 362.900 184.400 363.500 185.600 ;
        RECT 362.800 183.600 363.600 184.400 ;
        RECT 364.400 184.200 365.200 195.800 ;
        RECT 366.000 184.200 366.800 197.800 ;
        RECT 367.600 184.200 368.400 197.800 ;
        RECT 369.200 184.200 370.000 197.800 ;
        RECT 370.900 178.400 371.500 207.600 ;
        RECT 377.300 192.400 377.900 211.600 ;
        RECT 378.900 198.400 379.500 213.600 ;
        RECT 382.100 210.400 382.700 213.600 ;
        RECT 383.700 212.400 384.300 247.600 ;
        RECT 385.200 243.600 386.000 244.400 ;
        RECT 385.300 224.400 385.900 243.600 ;
        RECT 386.900 230.400 387.500 269.600 ;
        RECT 388.500 256.400 389.100 285.600 ;
        RECT 391.600 264.200 392.400 277.800 ;
        RECT 393.200 264.200 394.000 277.800 ;
        RECT 394.800 264.200 395.600 275.800 ;
        RECT 396.400 267.600 397.200 268.400 ;
        RECT 398.000 264.200 398.800 275.800 ;
        RECT 399.600 265.600 400.400 266.400 ;
        RECT 401.200 264.200 402.000 275.800 ;
        RECT 402.800 264.200 403.600 277.800 ;
        RECT 404.400 264.200 405.200 277.800 ;
        RECT 406.000 264.200 406.800 277.800 ;
        RECT 409.300 270.400 409.900 295.600 ;
        RECT 414.100 292.400 414.700 305.600 ;
        RECT 415.600 295.600 416.400 296.400 ;
        RECT 414.000 291.600 414.800 292.400 ;
        RECT 417.300 274.400 417.900 305.600 ;
        RECT 418.900 296.400 419.500 305.600 ;
        RECT 418.800 295.600 419.600 296.400 ;
        RECT 418.800 291.600 419.600 292.400 ;
        RECT 422.000 291.600 422.800 292.400 ;
        RECT 428.500 286.400 429.100 305.600 ;
        RECT 430.100 298.400 430.700 305.600 ;
        RECT 431.700 304.400 432.300 331.700 ;
        RECT 434.800 331.600 435.600 332.400 ;
        RECT 439.600 331.600 440.400 332.400 ;
        RECT 438.000 329.600 438.800 330.400 ;
        RECT 441.200 329.600 442.000 330.400 ;
        RECT 438.100 324.400 438.700 329.600 ;
        RECT 441.300 328.400 441.900 329.600 ;
        RECT 441.200 327.600 442.000 328.400 ;
        RECT 438.000 323.600 438.800 324.400 ;
        RECT 439.600 323.600 440.400 324.400 ;
        RECT 434.800 315.600 435.600 316.400 ;
        RECT 433.200 309.600 434.000 310.400 ;
        RECT 431.600 303.600 432.400 304.400 ;
        RECT 430.000 297.600 430.800 298.400 ;
        RECT 431.700 292.400 432.300 303.600 ;
        RECT 434.900 292.400 435.500 315.600 ;
        RECT 436.400 311.600 437.200 312.400 ;
        RECT 439.700 308.400 440.300 323.600 ;
        RECT 441.200 321.600 442.000 322.400 ;
        RECT 439.600 307.600 440.400 308.400 ;
        RECT 439.600 305.600 440.400 306.400 ;
        RECT 439.700 304.400 440.300 305.600 ;
        RECT 439.600 303.600 440.400 304.400 ;
        RECT 438.000 297.600 438.800 298.400 ;
        RECT 436.400 293.600 437.200 294.400 ;
        RECT 441.300 292.400 441.900 321.600 ;
        RECT 442.900 318.400 443.500 345.600 ;
        RECT 447.700 340.400 448.300 347.600 ;
        RECT 447.600 340.300 448.400 340.400 ;
        RECT 447.600 339.700 449.900 340.300 ;
        RECT 447.600 339.600 448.400 339.700 ;
        RECT 444.400 335.600 445.200 336.400 ;
        RECT 444.500 330.400 445.100 335.600 ;
        RECT 449.300 334.400 449.900 339.700 ;
        RECT 450.900 338.400 451.500 351.600 ;
        RECT 452.500 348.400 453.100 351.600 ;
        RECT 455.600 349.600 456.400 350.400 ;
        RECT 458.800 349.600 459.600 350.400 ;
        RECT 462.000 349.600 462.800 350.400 ;
        RECT 452.400 347.600 453.200 348.400 ;
        RECT 454.000 347.600 454.800 348.400 ;
        RECT 454.100 346.400 454.700 347.600 ;
        RECT 454.000 345.600 454.800 346.400 ;
        RECT 455.700 342.400 456.300 349.600 ;
        RECT 460.400 347.600 461.200 348.400 ;
        RECT 460.500 344.400 461.100 347.600 ;
        RECT 460.400 343.600 461.200 344.400 ;
        RECT 455.600 341.600 456.400 342.400 ;
        RECT 457.200 341.600 458.000 342.400 ;
        RECT 450.800 337.600 451.600 338.400 ;
        RECT 457.300 336.400 457.900 341.600 ;
        RECT 457.200 335.600 458.000 336.400 ;
        RECT 449.200 333.600 450.000 334.400 ;
        RECT 463.700 332.400 464.300 371.600 ;
        RECT 479.600 364.200 480.400 377.800 ;
        RECT 481.200 364.200 482.000 377.800 ;
        RECT 482.800 366.200 483.600 377.800 ;
        RECT 484.400 373.600 485.200 374.400 ;
        RECT 486.000 366.200 486.800 377.800 ;
        RECT 487.600 375.600 488.400 376.400 ;
        RECT 489.200 366.200 490.000 377.800 ;
        RECT 490.800 364.200 491.600 377.800 ;
        RECT 492.400 364.200 493.200 377.800 ;
        RECT 494.000 364.200 494.800 377.800 ;
        RECT 502.000 373.600 502.800 374.400 ;
        RECT 506.800 373.600 507.600 374.400 ;
        RECT 508.400 373.600 509.200 374.400 ;
        RECT 495.600 371.600 496.400 372.400 ;
        RECT 487.600 359.600 488.400 360.400 ;
        RECT 479.600 357.600 480.400 358.400 ;
        RECT 473.200 355.600 474.000 356.400 ;
        RECT 476.400 355.600 477.200 356.400 ;
        RECT 474.800 353.600 475.600 354.400 ;
        RECT 465.200 351.600 466.000 352.400 ;
        RECT 465.200 349.600 466.000 350.400 ;
        RECT 473.200 349.600 474.000 350.400 ;
        RECT 465.300 336.400 465.900 349.600 ;
        RECT 466.800 347.600 467.600 348.400 ;
        RECT 471.600 347.600 472.400 348.400 ;
        RECT 473.300 346.400 473.900 349.600 ;
        RECT 468.400 345.600 469.200 346.400 ;
        RECT 470.000 345.600 470.800 346.400 ;
        RECT 473.200 345.600 474.000 346.400 ;
        RECT 470.100 340.400 470.700 345.600 ;
        RECT 473.300 342.400 473.900 345.600 ;
        RECT 473.200 341.600 474.000 342.400 ;
        RECT 470.000 339.600 470.800 340.400 ;
        RECT 465.200 335.600 466.000 336.400 ;
        RECT 446.000 331.600 446.800 332.400 ;
        RECT 447.600 331.600 448.400 332.400 ;
        RECT 452.400 331.600 453.200 332.400 ;
        RECT 455.600 331.600 456.400 332.400 ;
        RECT 463.600 331.600 464.400 332.400 ;
        RECT 465.200 331.600 466.000 332.400 ;
        RECT 446.100 330.400 446.700 331.600 ;
        RECT 444.400 329.600 445.200 330.400 ;
        RECT 446.000 329.600 446.800 330.400 ;
        RECT 452.500 328.400 453.100 331.600 ;
        RECT 452.400 327.600 453.200 328.400 ;
        RECT 442.800 317.600 443.600 318.400 ;
        RECT 431.600 291.600 432.400 292.400 ;
        RECT 434.800 291.600 435.600 292.400 ;
        RECT 441.200 291.600 442.000 292.400 ;
        RECT 428.400 285.600 429.200 286.400 ;
        RECT 422.000 275.600 422.800 276.400 ;
        RECT 417.200 273.600 418.000 274.400 ;
        RECT 409.200 269.600 410.000 270.400 ;
        RECT 417.300 266.400 417.900 273.600 ;
        RECT 418.800 269.600 419.600 270.400 ;
        RECT 422.100 266.400 422.700 275.600 ;
        RECT 417.200 265.600 418.000 266.400 ;
        RECT 422.000 265.600 422.800 266.400 ;
        RECT 430.000 265.600 430.800 266.400 ;
        RECT 420.400 263.600 421.200 264.400 ;
        RECT 388.400 255.600 389.200 256.400 ;
        RECT 394.800 255.600 395.600 256.400 ;
        RECT 386.800 229.600 387.600 230.400 ;
        RECT 385.200 223.600 386.000 224.400 ;
        RECT 388.400 224.200 389.200 237.800 ;
        RECT 390.000 224.200 390.800 237.800 ;
        RECT 391.600 224.200 392.400 237.800 ;
        RECT 393.200 224.200 394.000 235.800 ;
        RECT 394.900 226.400 395.500 255.600 ;
        RECT 399.600 244.200 400.400 257.800 ;
        RECT 401.200 244.200 402.000 257.800 ;
        RECT 402.800 244.200 403.600 257.800 ;
        RECT 404.400 246.200 405.200 257.800 ;
        RECT 406.000 255.600 406.800 256.400 ;
        RECT 407.600 246.200 408.400 257.800 ;
        RECT 409.200 253.600 410.000 254.400 ;
        RECT 394.800 225.600 395.600 226.400 ;
        RECT 396.400 224.200 397.200 235.800 ;
        RECT 398.000 227.600 398.800 228.400 ;
        RECT 399.600 224.200 400.400 235.800 ;
        RECT 401.200 224.200 402.000 237.800 ;
        RECT 402.800 224.200 403.600 237.800 ;
        RECT 390.000 221.600 390.800 222.400 ;
        RECT 402.800 221.600 403.600 222.400 ;
        RECT 388.400 217.600 389.200 218.400 ;
        RECT 390.100 214.400 390.700 221.600 ;
        RECT 399.600 217.600 400.400 218.400 ;
        RECT 396.400 215.600 397.200 216.400 ;
        RECT 396.500 214.400 397.100 215.600 ;
        RECT 385.200 213.600 386.000 214.400 ;
        RECT 390.000 213.600 390.800 214.400 ;
        RECT 394.800 213.600 395.600 214.400 ;
        RECT 396.400 213.600 397.200 214.400 ;
        RECT 383.600 211.600 384.400 212.400 ;
        RECT 391.600 211.600 392.400 212.400 ;
        RECT 398.000 211.600 398.800 212.400 ;
        RECT 382.000 209.600 382.800 210.400 ;
        RECT 388.400 209.600 389.200 210.400 ;
        RECT 394.800 210.300 395.600 210.400 ;
        RECT 393.300 209.700 395.600 210.300 ;
        RECT 380.400 207.600 381.200 208.400 ;
        RECT 380.500 206.400 381.100 207.600 ;
        RECT 380.400 205.600 381.200 206.400 ;
        RECT 378.800 197.600 379.600 198.400 ;
        RECT 380.500 192.400 381.100 205.600 ;
        RECT 388.500 202.400 389.100 209.600 ;
        RECT 388.400 201.600 389.200 202.400 ;
        RECT 393.300 198.400 393.900 209.700 ;
        RECT 394.800 209.600 395.600 209.700 ;
        RECT 399.700 204.400 400.300 217.600 ;
        RECT 402.900 214.400 403.500 221.600 ;
        RECT 401.200 213.600 402.000 214.400 ;
        RECT 402.800 213.600 403.600 214.400 ;
        RECT 404.400 213.600 405.200 214.400 ;
        RECT 407.600 214.300 408.400 214.400 ;
        RECT 409.300 214.300 409.900 253.600 ;
        RECT 410.800 246.200 411.600 257.800 ;
        RECT 412.400 244.200 413.200 257.800 ;
        RECT 414.000 244.200 414.800 257.800 ;
        RECT 418.800 251.600 419.600 252.400 ;
        RECT 418.800 243.600 419.600 244.400 ;
        RECT 418.900 232.400 419.500 243.600 ;
        RECT 420.500 238.400 421.100 263.600 ;
        RECT 422.100 250.400 422.700 265.600 ;
        RECT 430.000 255.600 430.800 256.400 ;
        RECT 430.100 254.400 430.700 255.600 ;
        RECT 431.700 254.400 432.300 291.600 ;
        RECT 442.900 290.400 443.500 317.600 ;
        RECT 444.400 309.600 445.200 310.400 ;
        RECT 444.500 306.400 445.100 309.600 ;
        RECT 444.400 305.600 445.200 306.400 ;
        RECT 449.200 304.200 450.000 317.800 ;
        RECT 450.800 304.200 451.600 317.800 ;
        RECT 452.400 304.200 453.200 315.800 ;
        RECT 454.000 307.600 454.800 308.400 ;
        RECT 455.600 304.200 456.400 315.800 ;
        RECT 457.200 305.600 458.000 306.400 ;
        RECT 458.800 304.200 459.600 315.800 ;
        RECT 460.400 304.200 461.200 317.800 ;
        RECT 462.000 304.200 462.800 317.800 ;
        RECT 463.600 304.200 464.400 317.800 ;
        RECT 465.300 310.400 465.900 331.600 ;
        RECT 466.800 324.200 467.600 337.800 ;
        RECT 468.400 324.200 469.200 337.800 ;
        RECT 470.000 326.200 470.800 337.800 ;
        RECT 471.600 333.600 472.400 334.400 ;
        RECT 473.200 326.200 474.000 337.800 ;
        RECT 474.900 336.400 475.500 353.600 ;
        RECT 476.500 352.400 477.100 355.600 ;
        RECT 482.800 353.600 483.600 354.400 ;
        RECT 482.900 352.400 483.500 353.600 ;
        RECT 476.400 351.600 477.200 352.400 ;
        RECT 482.800 351.600 483.600 352.400 ;
        RECT 478.000 349.600 478.800 350.400 ;
        RECT 479.600 349.600 480.400 350.400 ;
        RECT 484.400 349.600 485.200 350.400 ;
        RECT 478.100 348.400 478.700 349.600 ;
        RECT 478.000 347.600 478.800 348.400 ;
        RECT 479.700 346.400 480.300 349.600 ;
        RECT 484.500 346.400 485.100 349.600 ;
        RECT 487.700 348.400 488.300 359.600 ;
        RECT 492.400 355.600 493.200 356.400 ;
        RECT 498.800 355.600 499.600 356.400 ;
        RECT 492.500 354.400 493.100 355.600 ;
        RECT 492.400 353.600 493.200 354.400 ;
        RECT 494.000 353.600 494.800 354.400 ;
        RECT 500.400 353.600 501.200 354.400 ;
        RECT 497.200 351.600 498.000 352.400 ;
        RECT 497.300 350.400 497.900 351.600 ;
        RECT 492.400 349.600 493.200 350.400 ;
        RECT 497.200 349.600 498.000 350.400 ;
        RECT 498.800 349.600 499.600 350.400 ;
        RECT 487.600 347.600 488.400 348.400 ;
        RECT 487.700 346.400 488.300 347.600 ;
        RECT 479.600 345.600 480.400 346.400 ;
        RECT 484.400 345.600 485.200 346.400 ;
        RECT 487.600 345.600 488.400 346.400 ;
        RECT 474.800 335.600 475.600 336.400 ;
        RECT 473.200 317.600 474.000 318.400 ;
        RECT 465.200 309.600 466.000 310.400 ;
        RECT 465.300 300.400 465.900 309.600 ;
        RECT 474.900 306.400 475.500 335.600 ;
        RECT 476.400 326.200 477.200 337.800 ;
        RECT 478.000 324.200 478.800 337.800 ;
        RECT 479.600 324.200 480.400 337.800 ;
        RECT 481.200 324.200 482.000 337.800 ;
        RECT 478.000 321.600 478.800 322.400 ;
        RECT 478.100 318.400 478.700 321.600 ;
        RECT 484.500 320.400 485.100 345.600 ;
        RECT 486.000 343.600 486.800 344.400 ;
        RECT 487.600 343.600 488.400 344.400 ;
        RECT 486.100 330.400 486.700 343.600 ;
        RECT 486.000 329.600 486.800 330.400 ;
        RECT 484.400 319.600 485.200 320.400 ;
        RECT 478.000 317.600 478.800 318.400 ;
        RECT 468.400 305.600 469.200 306.400 ;
        RECT 474.800 305.600 475.600 306.400 ;
        RECT 460.400 299.600 461.200 300.400 ;
        RECT 465.200 299.600 466.000 300.400 ;
        RECT 446.000 293.600 446.800 294.400 ;
        RECT 449.200 293.600 450.000 294.400 ;
        RECT 442.800 289.600 443.600 290.400 ;
        RECT 446.100 284.400 446.700 293.600 ;
        RECT 460.500 292.400 461.100 299.600 ;
        RECT 460.400 291.600 461.200 292.400 ;
        RECT 454.000 285.600 454.800 286.400 ;
        RECT 446.000 283.600 446.800 284.400 ;
        RECT 452.400 283.600 453.200 284.400 ;
        RECT 438.000 271.600 438.800 272.400 ;
        RECT 444.400 271.600 445.200 272.400 ;
        RECT 434.800 269.600 435.600 270.400 ;
        RECT 433.200 267.600 434.000 268.400 ;
        RECT 436.400 267.600 437.200 268.400 ;
        RECT 433.300 258.400 433.900 267.600 ;
        RECT 433.200 257.600 434.000 258.400 ;
        RECT 430.000 253.600 430.800 254.400 ;
        RECT 431.600 253.600 432.400 254.400 ;
        RECT 434.600 253.600 435.600 254.400 ;
        RECT 422.000 249.600 422.800 250.400 ;
        RECT 431.600 245.600 432.400 246.400 ;
        RECT 433.200 241.600 434.000 242.400 ;
        RECT 420.400 237.600 421.200 238.400 ;
        RECT 430.000 235.600 430.800 236.400 ;
        RECT 422.000 233.600 422.800 234.400 ;
        RECT 430.100 234.300 430.700 235.600 ;
        RECT 426.900 233.700 430.700 234.300 ;
        RECT 415.600 231.600 416.400 232.400 ;
        RECT 418.800 231.600 419.600 232.400 ;
        RECT 412.400 225.600 413.200 226.400 ;
        RECT 410.800 223.600 411.600 224.400 ;
        RECT 412.400 223.600 413.200 224.400 ;
        RECT 414.000 223.600 414.800 224.400 ;
        RECT 410.900 216.400 411.500 223.600 ;
        RECT 412.500 218.400 413.100 223.600 ;
        RECT 414.100 222.400 414.700 223.600 ;
        RECT 414.000 221.600 414.800 222.400 ;
        RECT 412.400 217.600 413.200 218.400 ;
        RECT 410.800 215.600 411.600 216.400 ;
        RECT 410.900 214.400 411.500 215.600 ;
        RECT 407.600 213.700 409.900 214.300 ;
        RECT 407.600 213.600 408.400 213.700 ;
        RECT 410.800 213.600 411.600 214.400 ;
        RECT 401.300 212.400 401.900 213.600 ;
        RECT 401.200 211.600 402.000 212.400 ;
        RECT 404.500 210.300 405.100 213.600 ;
        RECT 412.500 212.400 413.100 217.600 ;
        RECT 415.700 216.400 416.300 231.600 ;
        RECT 417.200 229.600 418.000 230.400 ;
        RECT 417.300 226.400 417.900 229.600 ;
        RECT 418.800 227.600 419.600 228.400 ;
        RECT 417.200 225.600 418.000 226.400 ;
        RECT 422.100 220.300 422.700 233.600 ;
        RECT 426.900 232.400 427.500 233.700 ;
        RECT 431.600 233.600 432.400 234.400 ;
        RECT 426.800 231.600 427.600 232.400 ;
        RECT 428.400 231.600 429.200 232.400 ;
        RECT 430.000 229.600 430.800 230.400 ;
        RECT 431.600 227.600 432.400 228.400 ;
        RECT 423.600 223.600 424.400 224.400 ;
        RECT 420.500 219.700 422.700 220.300 ;
        RECT 415.600 215.600 416.400 216.400 ;
        RECT 415.600 213.600 416.400 214.400 ;
        RECT 415.700 212.400 416.300 213.600 ;
        RECT 406.000 212.300 406.800 212.400 ;
        RECT 406.000 211.700 408.300 212.300 ;
        RECT 406.000 211.600 406.800 211.700 ;
        RECT 404.500 209.700 406.700 210.300 ;
        RECT 402.800 207.600 403.600 208.400 ;
        RECT 399.600 203.600 400.400 204.400 ;
        RECT 401.200 203.600 402.000 204.400 ;
        RECT 393.200 197.600 394.000 198.400 ;
        RECT 390.000 193.600 390.800 194.400 ;
        RECT 391.600 193.600 392.400 194.400 ;
        RECT 394.800 193.600 395.600 194.400 ;
        RECT 377.200 191.600 378.000 192.400 ;
        RECT 380.400 191.600 381.200 192.400 ;
        RECT 388.400 191.600 389.200 192.400 ;
        RECT 388.500 190.400 389.100 191.600 ;
        RECT 390.100 190.400 390.700 193.600 ;
        RECT 378.800 189.600 379.800 190.400 ;
        RECT 385.200 189.600 386.000 190.400 ;
        RECT 388.400 189.600 389.200 190.400 ;
        RECT 390.000 189.600 390.800 190.400 ;
        RECT 385.300 186.400 385.900 189.600 ;
        RECT 386.800 187.600 387.600 188.400 ;
        RECT 380.400 185.600 381.200 186.400 ;
        RECT 385.200 185.600 386.000 186.400 ;
        RECT 380.400 183.600 381.200 184.400 ;
        RECT 362.800 177.600 363.600 178.400 ;
        RECT 367.600 177.600 368.400 178.400 ;
        RECT 370.800 177.600 371.600 178.400 ;
        RECT 359.600 171.600 360.400 172.400 ;
        RECT 362.800 170.300 363.600 170.400 ;
        RECT 361.300 169.700 363.600 170.300 ;
        RECT 356.400 159.600 357.200 160.400 ;
        RECT 354.800 157.600 355.600 158.400 ;
        RECT 361.300 150.400 361.900 169.700 ;
        RECT 362.800 169.600 363.600 169.700 ;
        RECT 367.700 152.400 368.300 177.600 ;
        RECT 372.400 164.200 373.200 177.800 ;
        RECT 374.000 164.200 374.800 177.800 ;
        RECT 375.600 166.200 376.400 177.800 ;
        RECT 377.200 173.600 378.000 174.400 ;
        RECT 375.600 155.600 376.400 156.400 ;
        RECT 369.200 153.600 370.000 154.400 ;
        RECT 362.800 151.600 363.600 152.400 ;
        RECT 367.600 151.600 368.400 152.400 ;
        RECT 369.300 150.400 369.900 153.600 ;
        RECT 370.800 151.600 371.600 152.400 ;
        RECT 346.800 149.600 347.600 150.400 ;
        RECT 350.000 149.600 350.800 150.400 ;
        RECT 353.200 149.600 354.000 150.400 ;
        RECT 356.400 149.600 357.200 150.400 ;
        RECT 361.200 149.600 362.000 150.400 ;
        RECT 367.600 149.600 368.400 150.400 ;
        RECT 369.200 149.600 370.000 150.400 ;
        RECT 350.100 148.400 350.700 149.600 ;
        RECT 356.500 148.400 357.100 149.600 ;
        RECT 370.900 148.400 371.500 151.600 ;
        RECT 375.700 150.400 376.300 155.600 ;
        RECT 375.600 149.600 376.400 150.400 ;
        RECT 377.300 148.400 377.900 173.600 ;
        RECT 378.800 166.200 379.600 177.800 ;
        RECT 380.500 176.400 381.100 183.600 ;
        RECT 388.400 181.600 389.200 182.400 ;
        RECT 380.400 175.600 381.200 176.400 ;
        RECT 382.000 166.200 382.800 177.800 ;
        RECT 383.600 164.200 384.400 177.800 ;
        RECT 385.200 164.200 386.000 177.800 ;
        RECT 386.800 164.200 387.600 177.800 ;
        RECT 388.500 172.400 389.100 181.600 ;
        RECT 391.700 178.400 392.300 193.600 ;
        RECT 394.900 192.400 395.500 193.600 ;
        RECT 394.800 191.600 395.600 192.400 ;
        RECT 398.000 189.600 398.800 190.400 ;
        RECT 398.100 188.400 398.700 189.600 ;
        RECT 399.700 188.400 400.300 203.600 ;
        RECT 401.300 194.400 401.900 203.600 ;
        RECT 401.200 193.600 402.000 194.400 ;
        RECT 401.200 191.600 402.000 192.400 ;
        RECT 401.300 190.400 401.900 191.600 ;
        RECT 401.200 189.600 402.000 190.400 ;
        RECT 401.300 188.400 401.900 189.600 ;
        RECT 398.000 187.600 398.800 188.400 ;
        RECT 399.600 187.600 400.400 188.400 ;
        RECT 401.200 187.600 402.000 188.400 ;
        RECT 394.800 185.600 395.600 186.400 ;
        RECT 391.600 177.600 392.400 178.400 ;
        RECT 388.400 171.600 389.200 172.400 ;
        RECT 398.100 168.400 398.700 187.600 ;
        RECT 401.200 177.600 402.000 178.400 ;
        RECT 401.300 168.400 401.900 177.600 ;
        RECT 402.900 172.400 403.500 207.600 ;
        RECT 404.400 205.600 405.200 206.400 ;
        RECT 406.100 206.300 406.700 209.700 ;
        RECT 407.700 208.400 408.300 211.700 ;
        RECT 409.200 211.600 410.000 212.400 ;
        RECT 412.400 211.600 413.200 212.400 ;
        RECT 415.600 211.600 416.400 212.400 ;
        RECT 412.400 209.600 413.200 210.400 ;
        RECT 417.200 209.600 418.000 210.400 ;
        RECT 407.600 207.600 408.400 208.400 ;
        RECT 410.800 207.600 411.600 208.400 ;
        RECT 406.100 205.700 408.300 206.300 ;
        RECT 404.500 192.400 405.100 205.600 ;
        RECT 407.700 198.400 408.300 205.700 ;
        RECT 410.900 200.400 411.500 207.600 ;
        RECT 410.800 199.600 411.600 200.400 ;
        RECT 410.900 198.400 411.500 199.600 ;
        RECT 407.600 197.600 408.400 198.400 ;
        RECT 410.800 197.600 411.600 198.400 ;
        RECT 412.500 194.400 413.100 209.600 ;
        RECT 417.300 206.400 417.900 209.600 ;
        RECT 417.200 205.600 418.000 206.400 ;
        RECT 414.000 203.600 414.800 204.400 ;
        RECT 407.600 193.600 408.400 194.400 ;
        RECT 412.400 193.600 413.200 194.400 ;
        RECT 404.400 191.600 405.200 192.400 ;
        RECT 404.400 189.600 405.200 190.400 ;
        RECT 404.500 184.400 405.100 189.600 ;
        RECT 404.400 183.600 405.200 184.400 ;
        RECT 404.500 174.400 405.100 183.600 ;
        RECT 407.700 176.300 408.300 193.600 ;
        RECT 414.100 192.400 414.700 203.600 ;
        RECT 420.500 198.400 421.100 219.700 ;
        RECT 423.700 214.400 424.300 223.600 ;
        RECT 423.600 213.600 424.400 214.400 ;
        RECT 428.400 213.600 429.200 214.400 ;
        RECT 428.500 212.400 429.100 213.600 ;
        RECT 428.400 211.600 429.200 212.400 ;
        RECT 430.000 211.600 430.800 212.400 ;
        RECT 428.500 210.400 429.100 211.600 ;
        RECT 428.400 209.600 429.200 210.400 ;
        RECT 418.800 197.600 419.600 198.400 ;
        RECT 420.400 197.600 421.200 198.400 ;
        RECT 418.900 194.400 419.500 197.600 ;
        RECT 415.600 193.600 416.400 194.400 ;
        RECT 418.800 193.600 419.600 194.400 ;
        RECT 409.200 191.600 410.000 192.400 ;
        RECT 410.800 191.600 411.600 192.400 ;
        RECT 414.000 191.600 414.800 192.400 ;
        RECT 409.300 188.300 409.900 191.600 ;
        RECT 410.900 190.400 411.500 191.600 ;
        RECT 410.800 189.600 411.600 190.400 ;
        RECT 417.200 189.600 418.000 190.400 ;
        RECT 410.800 188.300 411.600 188.400 ;
        RECT 409.300 187.700 411.600 188.300 ;
        RECT 410.800 187.600 411.600 187.700 ;
        RECT 410.900 180.400 411.500 187.600 ;
        RECT 417.300 186.400 417.900 189.600 ;
        RECT 418.900 188.400 419.500 193.600 ;
        RECT 418.800 187.600 419.600 188.400 ;
        RECT 412.400 185.600 413.200 186.400 ;
        RECT 417.200 185.600 418.000 186.400 ;
        RECT 410.800 179.600 411.600 180.400 ;
        RECT 410.900 176.400 411.500 179.600 ;
        RECT 409.200 176.300 410.000 176.400 ;
        RECT 407.700 175.700 410.000 176.300 ;
        RECT 409.200 175.600 410.000 175.700 ;
        RECT 410.800 175.600 411.600 176.400 ;
        RECT 404.400 173.600 405.200 174.400 ;
        RECT 402.800 171.600 403.600 172.400 ;
        RECT 406.000 171.600 406.800 172.400 ;
        RECT 410.800 171.600 411.600 172.400 ;
        RECT 402.800 169.600 403.600 170.400 ;
        RECT 402.900 168.400 403.500 169.600 ;
        RECT 398.000 167.600 398.800 168.400 ;
        RECT 401.200 167.600 402.000 168.400 ;
        RECT 402.800 167.600 403.600 168.400 ;
        RECT 404.400 167.600 405.200 168.400 ;
        RECT 402.900 166.300 403.500 167.600 ;
        RECT 401.300 165.700 403.500 166.300 ;
        RECT 396.400 163.600 397.200 164.400 ;
        RECT 399.600 163.600 400.400 164.400 ;
        RECT 396.500 162.400 397.100 163.600 ;
        RECT 390.000 161.600 390.800 162.400 ;
        RECT 396.400 161.600 397.200 162.400 ;
        RECT 380.400 157.600 381.200 158.400 ;
        RECT 378.800 155.600 379.600 156.400 ;
        RECT 378.900 150.400 379.500 155.600 ;
        RECT 378.800 149.600 379.600 150.400 ;
        RECT 350.000 147.600 350.800 148.400 ;
        RECT 356.400 147.600 357.200 148.400 ;
        RECT 370.800 147.600 371.600 148.400 ;
        RECT 374.000 147.600 374.800 148.400 ;
        RECT 377.200 147.600 378.000 148.400 ;
        RECT 372.400 143.600 373.200 144.400 ;
        RECT 370.800 141.600 371.600 142.400 ;
        RECT 345.200 139.600 346.000 140.400 ;
        RECT 326.000 131.600 326.800 132.400 ;
        RECT 330.800 124.200 331.600 137.800 ;
        RECT 332.400 124.200 333.200 137.800 ;
        RECT 334.000 126.200 334.800 137.800 ;
        RECT 335.600 133.600 336.400 134.400 ;
        RECT 335.700 132.400 336.300 133.600 ;
        RECT 335.600 131.600 336.400 132.400 ;
        RECT 337.200 126.200 338.000 137.800 ;
        RECT 338.800 135.600 339.600 136.400 ;
        RECT 318.000 111.600 318.800 112.400 ;
        RECT 318.100 110.400 318.700 111.600 ;
        RECT 318.000 109.600 318.800 110.400 ;
        RECT 321.200 109.600 322.000 110.400 ;
        RECT 316.400 107.600 317.200 108.400 ;
        RECT 321.300 106.400 321.900 109.600 ;
        RECT 324.400 107.600 325.200 108.400 ;
        RECT 324.500 106.400 325.100 107.600 ;
        RECT 338.900 106.400 339.500 135.600 ;
        RECT 340.400 126.200 341.200 137.800 ;
        RECT 342.000 124.200 342.800 137.800 ;
        RECT 343.600 124.200 344.400 137.800 ;
        RECT 345.200 124.200 346.000 137.800 ;
        RECT 370.900 136.400 371.500 141.600 ;
        RECT 372.500 136.400 373.100 143.600 ;
        RECT 374.100 140.400 374.700 147.600 ;
        RECT 374.000 139.600 374.800 140.400 ;
        RECT 356.400 135.600 357.200 136.400 ;
        RECT 361.200 135.600 362.000 136.400 ;
        RECT 362.800 135.600 363.600 136.400 ;
        RECT 370.800 135.600 371.600 136.400 ;
        RECT 372.400 135.600 373.200 136.400 ;
        RECT 370.900 134.400 371.500 135.600 ;
        RECT 374.100 134.400 374.700 139.600 ;
        RECT 378.800 135.600 379.600 136.400 ;
        RECT 361.200 133.600 362.000 134.400 ;
        RECT 364.400 133.600 365.200 134.400 ;
        RECT 366.000 133.600 366.800 134.400 ;
        RECT 370.800 133.600 371.600 134.400 ;
        RECT 374.000 133.600 374.800 134.400 ;
        RECT 375.600 133.600 376.400 134.400 ;
        RECT 342.000 109.600 342.800 110.400 ;
        RECT 321.200 105.600 322.000 106.400 ;
        RECT 324.400 105.600 325.200 106.400 ;
        RECT 338.800 105.600 339.600 106.400 ;
        RECT 314.800 91.600 315.600 92.400 ;
        RECT 313.200 73.600 314.000 74.400 ;
        RECT 308.400 69.600 309.200 70.400 ;
        RECT 310.000 69.600 310.800 70.400 ;
        RECT 308.500 68.400 309.100 69.600 ;
        RECT 308.400 67.600 309.200 68.400 ;
        RECT 311.600 67.600 312.400 68.400 ;
        RECT 311.700 66.400 312.300 67.600 ;
        RECT 311.600 65.600 312.400 66.400 ;
        RECT 303.600 63.600 304.400 64.400 ;
        RECT 290.800 59.600 291.600 60.400 ;
        RECT 279.600 49.600 280.400 50.400 ;
        RECT 284.400 49.600 285.200 50.400 ;
        RECT 247.600 41.600 248.400 42.400 ;
        RECT 252.400 41.600 253.200 42.400 ;
        RECT 226.800 31.600 227.600 32.400 ;
        RECT 230.000 31.600 230.800 32.400 ;
        RECT 217.200 27.600 218.000 28.400 ;
        RECT 223.600 27.600 224.400 28.400 ;
        RECT 214.000 25.600 214.800 26.400 ;
        RECT 212.500 23.700 214.700 24.300 ;
        RECT 185.200 21.600 186.000 22.400 ;
        RECT 198.000 21.600 198.800 22.400 ;
        RECT 202.800 21.600 203.600 22.400 ;
        RECT 166.000 11.600 166.800 12.400 ;
        RECT 166.100 10.400 166.700 11.600 ;
        RECT 166.000 9.600 166.800 10.400 ;
        RECT 185.200 9.600 186.000 10.400 ;
        RECT 190.000 4.200 190.800 17.800 ;
        RECT 191.600 4.200 192.400 17.800 ;
        RECT 193.200 6.200 194.000 17.800 ;
        RECT 194.800 13.600 195.600 14.400 ;
        RECT 196.400 6.200 197.200 17.800 ;
        RECT 198.100 16.400 198.700 21.600 ;
        RECT 214.100 18.400 214.700 23.700 ;
        RECT 198.000 15.600 198.800 16.400 ;
        RECT 199.600 6.200 200.400 17.800 ;
        RECT 201.200 4.200 202.000 17.800 ;
        RECT 202.800 4.200 203.600 17.800 ;
        RECT 204.400 4.200 205.200 17.800 ;
        RECT 214.000 17.600 214.800 18.400 ;
        RECT 217.300 14.400 217.900 27.600 ;
        RECT 223.700 26.400 224.300 27.600 ;
        RECT 223.600 25.600 224.400 26.400 ;
        RECT 226.800 25.600 227.600 26.400 ;
        RECT 226.900 14.400 227.500 25.600 ;
        RECT 217.200 13.600 218.000 14.400 ;
        RECT 223.600 13.600 224.400 14.400 ;
        RECT 226.800 13.600 227.600 14.400 ;
        RECT 222.000 11.600 222.800 12.400 ;
        RECT 225.200 11.600 226.000 12.400 ;
        RECT 222.100 10.400 222.700 11.600 ;
        RECT 230.100 10.400 230.700 31.600 ;
        RECT 231.600 23.600 232.400 24.400 ;
        RECT 234.800 23.600 235.600 24.400 ;
        RECT 241.200 24.200 242.000 37.800 ;
        RECT 242.800 24.200 243.600 37.800 ;
        RECT 244.400 24.200 245.200 37.800 ;
        RECT 246.000 24.200 246.800 35.800 ;
        RECT 247.700 26.400 248.300 41.600 ;
        RECT 247.600 25.600 248.400 26.400 ;
        RECT 249.200 24.200 250.000 35.800 ;
        RECT 250.800 27.600 251.600 28.400 ;
        RECT 250.900 24.400 251.500 27.600 ;
        RECT 250.800 23.600 251.600 24.400 ;
        RECT 252.400 24.200 253.200 35.800 ;
        RECT 254.000 24.200 254.800 37.800 ;
        RECT 255.600 24.200 256.400 37.800 ;
        RECT 262.100 32.400 262.700 49.600 ;
        RECT 279.600 43.600 280.400 44.400 ;
        RECT 289.200 44.200 290.000 57.800 ;
        RECT 290.800 44.200 291.600 57.800 ;
        RECT 292.400 46.200 293.200 57.800 ;
        RECT 294.100 54.400 294.700 63.600 ;
        RECT 297.200 59.600 298.000 60.400 ;
        RECT 294.000 53.600 294.800 54.400 ;
        RECT 295.600 46.200 296.400 57.800 ;
        RECT 297.300 56.400 297.900 59.600 ;
        RECT 313.300 58.400 313.900 73.600 ;
        RECT 314.900 72.400 315.500 91.600 ;
        RECT 318.000 84.200 318.800 97.800 ;
        RECT 319.600 84.200 320.400 97.800 ;
        RECT 321.200 84.200 322.000 97.800 ;
        RECT 322.800 86.200 323.600 97.800 ;
        RECT 324.500 96.400 325.100 105.600 ;
        RECT 342.100 100.400 342.700 109.600 ;
        RECT 346.800 104.200 347.600 117.800 ;
        RECT 348.400 104.200 349.200 117.800 ;
        RECT 350.000 104.200 350.800 115.800 ;
        RECT 351.600 107.600 352.400 108.400 ;
        RECT 353.200 104.200 354.000 115.800 ;
        RECT 354.800 105.600 355.600 106.400 ;
        RECT 337.200 99.600 338.000 100.400 ;
        RECT 342.000 99.600 342.800 100.400 ;
        RECT 324.400 95.600 325.200 96.400 ;
        RECT 326.000 86.200 326.800 97.800 ;
        RECT 327.600 93.600 328.400 94.400 ;
        RECT 329.200 86.200 330.000 97.800 ;
        RECT 326.000 83.600 326.800 84.400 ;
        RECT 330.800 84.200 331.600 97.800 ;
        RECT 332.400 84.200 333.200 97.800 ;
        RECT 337.300 90.400 337.900 99.600 ;
        RECT 354.900 96.400 355.500 105.600 ;
        RECT 356.400 104.200 357.200 115.800 ;
        RECT 358.000 104.200 358.800 117.800 ;
        RECT 359.600 104.200 360.400 117.800 ;
        RECT 361.200 104.200 362.000 117.800 ;
        RECT 364.500 116.400 365.100 133.600 ;
        RECT 366.100 132.400 366.700 133.600 ;
        RECT 366.000 131.600 366.800 132.400 ;
        RECT 367.600 131.600 368.400 132.400 ;
        RECT 369.200 131.600 370.000 132.400 ;
        RECT 372.400 131.600 373.200 132.400 ;
        RECT 364.400 115.600 365.200 116.400 ;
        RECT 369.300 110.400 369.900 131.600 ;
        RECT 369.200 109.600 370.000 110.400 ;
        RECT 372.500 104.400 373.100 131.600 ;
        RECT 375.700 110.400 376.300 133.600 ;
        RECT 377.200 123.600 378.000 124.400 ;
        RECT 377.300 118.400 377.900 123.600 ;
        RECT 378.900 122.400 379.500 135.600 ;
        RECT 378.800 121.600 379.600 122.400 ;
        RECT 377.200 117.600 378.000 118.400 ;
        RECT 375.600 109.600 376.400 110.400 ;
        RECT 378.800 109.600 379.600 110.400 ;
        RECT 374.000 107.600 374.800 108.400 ;
        RECT 377.200 107.600 378.000 108.400 ;
        RECT 370.800 103.600 371.600 104.400 ;
        RECT 372.400 103.600 373.200 104.400 ;
        RECT 370.900 100.400 371.500 103.600 ;
        RECT 374.100 102.400 374.700 107.600 ;
        RECT 374.000 101.600 374.800 102.400 ;
        RECT 370.800 99.600 371.600 100.400 ;
        RECT 354.800 95.600 355.600 96.400 ;
        RECT 342.000 93.600 342.800 94.400 ;
        RECT 345.200 93.600 346.000 94.400 ;
        RECT 353.200 93.600 354.000 94.400 ;
        RECT 337.200 89.600 338.000 90.400 ;
        RECT 326.100 76.400 326.700 83.600 ;
        RECT 326.000 75.600 326.800 76.400 ;
        RECT 334.000 75.600 334.800 76.400 ;
        RECT 314.800 71.600 315.600 72.400 ;
        RECT 314.900 70.400 315.500 71.600 ;
        RECT 314.800 69.600 315.600 70.400 ;
        RECT 326.100 68.400 326.700 75.600 ;
        RECT 330.800 71.600 331.600 72.400 ;
        RECT 330.900 70.400 331.500 71.600 ;
        RECT 327.600 69.600 328.400 70.400 ;
        RECT 330.800 69.600 331.600 70.400 ;
        RECT 327.700 68.400 328.300 69.600 ;
        RECT 319.600 67.600 320.400 68.400 ;
        RECT 326.000 67.600 326.800 68.400 ;
        RECT 327.600 67.600 328.400 68.400 ;
        RECT 319.700 66.400 320.300 67.600 ;
        RECT 319.600 65.600 320.400 66.400 ;
        RECT 324.400 65.600 325.200 66.400 ;
        RECT 321.200 63.600 322.000 64.400 ;
        RECT 297.200 55.600 298.000 56.400 ;
        RECT 298.800 46.200 299.600 57.800 ;
        RECT 300.400 44.200 301.200 57.800 ;
        RECT 302.000 44.200 302.800 57.800 ;
        RECT 303.600 44.200 304.400 57.800 ;
        RECT 313.200 57.600 314.000 58.400 ;
        RECT 318.000 53.600 318.800 54.400 ;
        RECT 321.300 52.400 321.900 63.600 ;
        RECT 324.500 56.400 325.100 65.600 ;
        RECT 327.600 63.600 328.400 64.400 ;
        RECT 335.600 63.600 336.400 64.400 ;
        RECT 327.700 60.400 328.300 63.600 ;
        RECT 327.600 59.600 328.400 60.400 ;
        RECT 324.400 55.600 325.200 56.400 ;
        RECT 321.200 51.600 322.000 52.400 ;
        RECT 314.800 49.600 315.600 50.400 ;
        RECT 262.000 31.600 262.800 32.400 ;
        RECT 270.000 29.600 270.800 30.400 ;
        RECT 279.700 28.400 280.300 43.600 ;
        RECT 281.200 31.600 282.000 32.400 ;
        RECT 281.300 30.400 281.900 31.600 ;
        RECT 281.200 29.600 282.000 30.400 ;
        RECT 287.600 29.600 288.400 30.400 ;
        RECT 270.000 27.600 270.800 28.400 ;
        RECT 271.600 27.600 272.400 28.400 ;
        RECT 279.600 27.600 280.400 28.400 ;
        RECT 265.200 25.600 266.000 26.400 ;
        RECT 231.700 18.400 232.300 23.600 ;
        RECT 233.200 21.600 234.000 22.400 ;
        RECT 231.600 17.600 232.400 18.400 ;
        RECT 233.300 14.400 233.900 21.600 ;
        RECT 234.900 18.400 235.500 23.600 ;
        RECT 244.400 21.600 245.200 22.400 ;
        RECT 234.800 17.600 235.600 18.400 ;
        RECT 238.000 17.600 238.800 18.400 ;
        RECT 238.100 14.400 238.700 17.600 ;
        RECT 239.600 15.600 240.400 16.400 ;
        RECT 233.200 13.600 234.000 14.400 ;
        RECT 238.000 13.600 238.800 14.400 ;
        RECT 239.700 12.400 240.300 15.600 ;
        RECT 244.500 14.400 245.100 21.600 ;
        RECT 262.000 19.600 262.800 20.400 ;
        RECT 246.000 17.600 246.800 18.400 ;
        RECT 244.400 13.600 245.200 14.400 ;
        RECT 246.100 12.400 246.700 17.600 ;
        RECT 262.100 14.400 262.700 19.600 ;
        RECT 265.300 18.400 265.900 25.600 ;
        RECT 266.800 23.600 267.600 24.400 ;
        RECT 266.900 20.400 267.500 23.600 ;
        RECT 270.100 22.400 270.700 27.600 ;
        RECT 271.700 24.400 272.300 27.600 ;
        RECT 271.600 23.600 272.400 24.400 ;
        RECT 270.000 21.600 270.800 22.400 ;
        RECT 266.800 19.600 267.600 20.400 ;
        RECT 265.200 17.600 266.000 18.400 ;
        RECT 266.800 17.600 267.600 18.400 ;
        RECT 266.900 16.400 267.500 17.600 ;
        RECT 265.200 15.600 266.000 16.400 ;
        RECT 266.800 15.600 267.600 16.400 ;
        RECT 255.600 13.600 256.400 14.400 ;
        RECT 257.200 13.600 258.000 14.400 ;
        RECT 262.000 13.600 262.800 14.400 ;
        RECT 263.600 13.600 264.400 14.400 ;
        RECT 239.600 11.600 240.400 12.400 ;
        RECT 242.800 11.600 243.600 12.400 ;
        RECT 246.000 11.600 246.800 12.400 ;
        RECT 254.000 11.600 254.800 12.400 ;
        RECT 255.600 11.600 256.400 12.400 ;
        RECT 242.900 10.400 243.500 11.600 ;
        RECT 254.100 10.400 254.700 11.600 ;
        RECT 257.300 10.400 257.900 13.600 ;
        RECT 265.300 12.400 265.900 15.600 ;
        RECT 270.100 14.400 270.700 21.600 ;
        RECT 268.400 13.600 269.200 14.400 ;
        RECT 270.000 13.600 270.800 14.400 ;
        RECT 278.000 13.600 278.800 14.400 ;
        RECT 279.600 13.600 280.400 14.400 ;
        RECT 262.000 12.300 262.800 12.400 ;
        RECT 262.000 11.700 264.300 12.300 ;
        RECT 262.000 11.600 262.800 11.700 ;
        RECT 222.000 9.600 222.800 10.400 ;
        RECT 225.200 9.600 226.000 10.400 ;
        RECT 230.000 10.300 230.800 10.400 ;
        RECT 231.600 10.300 232.400 10.400 ;
        RECT 230.000 9.700 232.400 10.300 ;
        RECT 230.000 9.600 230.800 9.700 ;
        RECT 231.600 9.600 232.400 9.700 ;
        RECT 236.400 9.600 237.200 10.400 ;
        RECT 242.800 9.600 243.600 10.400 ;
        RECT 249.200 9.600 250.000 10.400 ;
        RECT 254.000 9.600 254.800 10.400 ;
        RECT 257.200 9.600 258.000 10.400 ;
        RECT 263.700 10.300 264.300 11.700 ;
        RECT 265.200 11.600 266.000 12.400 ;
        RECT 271.600 11.600 272.400 12.400 ;
        RECT 278.100 10.400 278.700 13.600 ;
        RECT 281.300 12.400 281.900 29.600 ;
        RECT 286.000 27.600 286.800 28.400 ;
        RECT 287.600 27.600 288.400 28.400 ;
        RECT 287.700 18.400 288.300 27.600 ;
        RECT 289.200 23.600 290.000 24.400 ;
        RECT 298.800 24.200 299.600 37.800 ;
        RECT 300.400 24.200 301.200 37.800 ;
        RECT 302.000 24.200 302.800 37.800 ;
        RECT 303.600 24.200 304.400 35.800 ;
        RECT 305.200 25.600 306.000 26.400 ;
        RECT 289.300 18.400 289.900 23.600 ;
        RECT 305.300 20.300 305.900 25.600 ;
        RECT 306.800 24.200 307.600 35.800 ;
        RECT 308.400 27.600 309.200 28.400 ;
        RECT 310.000 24.200 310.800 35.800 ;
        RECT 311.600 24.200 312.400 37.800 ;
        RECT 313.200 24.200 314.000 37.800 ;
        RECT 314.900 32.000 315.500 49.600 ;
        RECT 314.800 31.200 315.600 32.000 ;
        RECT 306.800 20.300 307.600 20.400 ;
        RECT 305.300 19.700 307.600 20.300 ;
        RECT 306.800 19.600 307.600 19.700 ;
        RECT 287.600 17.600 288.400 18.400 ;
        RECT 289.200 17.600 290.000 18.400 ;
        RECT 281.200 11.600 282.000 12.400 ;
        RECT 290.600 11.600 291.600 12.400 ;
        RECT 265.200 10.300 266.000 10.400 ;
        RECT 263.700 9.700 266.000 10.300 ;
        RECT 265.200 9.600 266.000 9.700 ;
        RECT 274.800 9.600 275.600 10.400 ;
        RECT 278.000 9.600 278.800 10.400 ;
        RECT 287.600 9.600 288.400 10.400 ;
        RECT 225.300 8.400 225.900 9.600 ;
        RECT 236.500 8.400 237.100 9.600 ;
        RECT 225.200 7.600 226.000 8.400 ;
        RECT 228.400 7.600 229.200 8.400 ;
        RECT 236.400 7.600 237.200 8.400 ;
        RECT 239.600 7.600 240.400 8.400 ;
        RECT 254.000 7.600 254.800 8.400 ;
        RECT 300.400 4.200 301.200 17.800 ;
        RECT 302.000 4.200 302.800 17.800 ;
        RECT 303.600 4.200 304.400 17.800 ;
        RECT 305.200 6.200 306.000 17.800 ;
        RECT 306.900 16.400 307.500 19.600 ;
        RECT 306.800 15.600 307.600 16.400 ;
        RECT 308.400 6.200 309.200 17.800 ;
        RECT 310.000 13.600 310.800 14.400 ;
        RECT 310.100 8.400 310.700 13.600 ;
        RECT 310.000 7.600 310.800 8.400 ;
        RECT 311.600 6.200 312.400 17.800 ;
        RECT 313.200 4.200 314.000 17.800 ;
        RECT 314.800 4.200 315.600 17.800 ;
        RECT 321.300 10.400 321.900 51.600 ;
        RECT 327.600 44.200 328.400 57.800 ;
        RECT 329.200 44.200 330.000 57.800 ;
        RECT 330.800 46.200 331.600 57.800 ;
        RECT 332.400 57.600 333.200 58.400 ;
        RECT 332.500 54.400 333.100 57.600 ;
        RECT 332.400 53.600 333.200 54.400 ;
        RECT 334.000 46.200 334.800 57.800 ;
        RECT 335.700 56.400 336.300 63.600 ;
        RECT 337.300 62.400 337.900 89.600 ;
        RECT 342.100 84.400 342.700 93.600 ;
        RECT 343.600 91.600 344.400 92.400 ;
        RECT 348.400 91.600 349.200 92.400 ;
        RECT 348.500 90.400 349.100 91.600 ;
        RECT 348.400 89.600 349.200 90.400 ;
        RECT 342.000 83.600 342.800 84.400 ;
        RECT 353.300 82.400 353.900 93.600 ;
        RECT 353.200 81.600 354.000 82.400 ;
        RECT 348.400 64.200 349.200 77.800 ;
        RECT 350.000 64.200 350.800 77.800 ;
        RECT 351.600 64.200 352.400 77.800 ;
        RECT 353.200 64.200 354.000 75.800 ;
        RECT 354.900 66.400 355.500 95.600 ;
        RECT 362.800 84.200 363.600 97.800 ;
        RECT 364.400 84.200 365.200 97.800 ;
        RECT 366.000 86.200 366.800 97.800 ;
        RECT 367.600 97.600 368.400 98.400 ;
        RECT 367.700 94.400 368.300 97.600 ;
        RECT 367.600 93.600 368.400 94.400 ;
        RECT 367.600 91.600 368.400 92.400 ;
        RECT 354.800 65.600 355.600 66.400 ;
        RECT 354.900 64.400 355.500 65.600 ;
        RECT 354.800 63.600 355.600 64.400 ;
        RECT 356.400 64.200 357.200 75.800 ;
        RECT 358.000 73.600 358.800 74.400 ;
        RECT 358.100 68.400 358.700 73.600 ;
        RECT 358.000 67.600 358.800 68.400 ;
        RECT 359.600 64.200 360.400 75.800 ;
        RECT 361.200 64.200 362.000 77.800 ;
        RECT 362.800 64.200 363.600 77.800 ;
        RECT 367.700 70.400 368.300 91.600 ;
        RECT 369.200 86.200 370.000 97.800 ;
        RECT 370.800 95.600 371.600 96.400 ;
        RECT 372.400 86.200 373.200 97.800 ;
        RECT 374.000 84.200 374.800 97.800 ;
        RECT 375.600 84.200 376.400 97.800 ;
        RECT 377.200 84.200 378.000 97.800 ;
        RECT 378.800 91.600 379.600 92.400 ;
        RECT 378.900 84.400 379.500 91.600 ;
        RECT 378.800 83.600 379.600 84.400 ;
        RECT 378.800 79.600 379.600 80.400 ;
        RECT 372.400 75.600 373.200 76.400 ;
        RECT 367.600 69.600 368.400 70.400 ;
        RECT 369.200 69.600 370.000 70.400 ;
        RECT 367.700 62.400 368.300 69.600 ;
        RECT 337.200 61.600 338.000 62.400 ;
        RECT 343.600 61.600 344.400 62.400 ;
        RECT 367.600 61.600 368.400 62.400 ;
        RECT 335.600 55.600 336.400 56.400 ;
        RECT 337.200 46.200 338.000 57.800 ;
        RECT 338.800 44.200 339.600 57.800 ;
        RECT 340.400 44.200 341.200 57.800 ;
        RECT 342.000 44.200 342.800 57.800 ;
        RECT 343.700 52.400 344.300 61.600 ;
        RECT 367.600 57.600 368.400 58.400 ;
        RECT 354.800 55.600 355.600 56.400 ;
        RECT 358.000 55.600 358.800 56.400 ;
        RECT 359.600 55.600 360.400 56.400 ;
        RECT 358.000 53.600 358.800 54.400 ;
        RECT 358.100 52.400 358.700 53.600 ;
        RECT 359.700 52.400 360.300 55.600 ;
        RECT 369.300 52.400 369.900 69.600 ;
        RECT 372.500 68.400 373.100 75.600 ;
        RECT 375.600 73.600 376.400 74.400 ;
        RECT 377.200 73.600 378.000 74.400 ;
        RECT 375.700 70.400 376.300 73.600 ;
        RECT 377.300 72.400 377.900 73.600 ;
        RECT 377.200 71.600 378.000 72.400 ;
        RECT 374.000 69.600 374.800 70.400 ;
        RECT 375.600 69.600 376.400 70.400 ;
        RECT 378.900 68.400 379.500 79.600 ;
        RECT 380.500 70.400 381.100 157.600 ;
        RECT 382.000 151.600 382.800 152.400 ;
        RECT 388.400 151.600 389.200 152.400 ;
        RECT 382.100 134.400 382.700 151.600 ;
        RECT 383.600 149.600 384.400 150.400 ;
        RECT 385.200 149.600 386.000 150.400 ;
        RECT 386.800 149.600 387.600 150.400 ;
        RECT 385.300 148.300 385.900 149.600 ;
        RECT 386.800 148.300 387.600 148.400 ;
        RECT 385.300 147.700 387.600 148.300 ;
        RECT 386.800 147.600 387.600 147.700 ;
        RECT 383.600 145.600 384.400 146.400 ;
        RECT 382.000 133.600 382.800 134.400 ;
        RECT 383.700 132.400 384.300 145.600 ;
        RECT 385.200 133.600 386.000 134.400 ;
        RECT 382.000 131.600 382.800 132.400 ;
        RECT 383.600 131.600 384.400 132.400 ;
        RECT 382.000 121.600 382.800 122.400 ;
        RECT 382.100 118.400 382.700 121.600 ;
        RECT 382.000 117.600 382.800 118.400 ;
        RECT 385.300 114.300 385.900 133.600 ;
        RECT 383.700 113.700 385.900 114.300 ;
        RECT 383.700 108.400 384.300 113.700 ;
        RECT 385.200 111.600 386.000 112.400 ;
        RECT 385.300 110.400 385.900 111.600 ;
        RECT 385.200 109.600 386.000 110.400 ;
        RECT 383.600 107.600 384.400 108.400 ;
        RECT 383.600 105.600 384.400 106.400 ;
        RECT 383.700 100.400 384.300 105.600 ;
        RECT 385.200 103.600 386.000 104.400 ;
        RECT 383.600 99.600 384.400 100.400 ;
        RECT 385.300 72.400 385.900 103.600 ;
        RECT 386.900 90.400 387.500 147.600 ;
        RECT 388.400 146.300 389.200 146.400 ;
        RECT 390.100 146.300 390.700 161.600 ;
        RECT 394.800 153.600 395.600 154.400 ;
        RECT 398.000 153.600 398.800 154.400 ;
        RECT 393.200 149.600 394.000 150.400 ;
        RECT 394.900 148.400 395.500 153.600 ;
        RECT 396.400 151.600 397.200 152.400 ;
        RECT 399.700 150.400 400.300 163.600 ;
        RECT 401.300 152.400 401.900 165.700 ;
        RECT 402.800 163.600 403.600 164.400 ;
        RECT 401.200 151.600 402.000 152.400 ;
        RECT 401.300 150.400 401.900 151.600 ;
        RECT 399.600 149.600 400.400 150.400 ;
        RECT 401.200 149.600 402.000 150.400 ;
        RECT 394.800 147.600 395.600 148.400 ;
        RECT 388.400 145.700 390.700 146.300 ;
        RECT 388.400 145.600 389.200 145.700 ;
        RECT 390.100 132.400 390.700 145.700 ;
        RECT 393.200 145.600 394.000 146.400 ;
        RECT 393.300 136.400 393.900 145.600 ;
        RECT 396.400 143.600 397.200 144.400 ;
        RECT 401.200 143.600 402.000 144.400 ;
        RECT 396.500 138.400 397.100 143.600 ;
        RECT 396.400 137.600 397.200 138.400 ;
        RECT 393.200 136.300 394.000 136.400 ;
        RECT 393.200 135.700 395.500 136.300 ;
        RECT 393.200 135.600 394.000 135.700 ;
        RECT 390.000 131.600 390.800 132.400 ;
        RECT 388.400 127.600 389.200 128.400 ;
        RECT 391.600 123.600 392.400 124.400 ;
        RECT 390.000 119.600 390.800 120.400 ;
        RECT 390.100 118.400 390.700 119.600 ;
        RECT 390.000 117.600 390.800 118.400 ;
        RECT 391.700 112.300 392.300 123.600 ;
        RECT 393.200 115.600 394.000 116.400 ;
        RECT 390.100 111.700 392.300 112.300 ;
        RECT 390.100 108.400 390.700 111.700 ;
        RECT 393.300 110.400 393.900 115.600 ;
        RECT 391.600 109.600 392.400 110.400 ;
        RECT 393.200 109.600 394.000 110.400 ;
        RECT 390.000 107.600 390.800 108.400 ;
        RECT 390.100 96.400 390.700 107.600 ;
        RECT 391.700 106.400 392.300 109.600 ;
        RECT 391.600 105.600 392.400 106.400 ;
        RECT 393.200 105.600 394.000 106.400 ;
        RECT 393.300 100.400 393.900 105.600 ;
        RECT 394.900 104.400 395.500 135.700 ;
        RECT 399.600 107.600 400.400 108.400 ;
        RECT 396.400 105.600 397.200 106.400 ;
        RECT 394.800 103.600 395.600 104.400 ;
        RECT 394.800 101.600 395.600 102.400 ;
        RECT 393.200 99.600 394.000 100.400 ;
        RECT 390.000 95.600 390.800 96.400 ;
        RECT 393.300 94.400 393.900 99.600 ;
        RECT 393.200 93.600 394.000 94.400 ;
        RECT 390.000 91.600 390.800 92.400 ;
        RECT 386.800 89.600 387.600 90.400 ;
        RECT 390.000 89.600 390.800 90.400 ;
        RECT 393.200 89.600 394.000 90.400 ;
        RECT 388.400 87.600 389.200 88.400 ;
        RECT 385.200 71.600 386.000 72.400 ;
        RECT 385.300 70.400 385.900 71.600 ;
        RECT 388.500 70.400 389.100 87.600 ;
        RECT 391.600 83.600 392.400 84.400 ;
        RECT 391.700 74.400 392.300 83.600 ;
        RECT 391.600 73.600 392.400 74.400 ;
        RECT 394.900 72.400 395.500 101.600 ;
        RECT 396.500 94.400 397.100 105.600 ;
        RECT 396.400 93.600 397.200 94.400 ;
        RECT 398.000 93.600 398.800 94.400 ;
        RECT 399.600 94.300 400.400 94.400 ;
        RECT 401.300 94.300 401.900 143.600 ;
        RECT 402.900 124.400 403.500 163.600 ;
        RECT 404.500 154.400 405.100 167.600 ;
        RECT 407.600 163.600 408.400 164.400 ;
        RECT 406.000 159.600 406.800 160.400 ;
        RECT 404.400 153.600 405.200 154.400 ;
        RECT 406.100 150.400 406.700 159.600 ;
        RECT 407.600 153.600 408.400 154.400 ;
        RECT 407.700 152.400 408.300 153.600 ;
        RECT 407.600 151.600 408.400 152.400 ;
        RECT 409.200 151.600 410.000 152.400 ;
        RECT 407.700 150.400 408.300 151.600 ;
        RECT 410.900 150.400 411.500 171.600 ;
        RECT 412.500 150.400 413.100 185.600 ;
        RECT 417.300 156.400 417.900 185.600 ;
        RECT 417.200 155.600 418.000 156.400 ;
        RECT 414.000 151.600 414.800 152.400 ;
        RECT 420.500 152.300 421.100 197.600 ;
        RECT 430.100 194.400 430.700 211.600 ;
        RECT 430.000 193.600 430.800 194.400 ;
        RECT 423.600 191.600 424.400 192.400 ;
        RECT 431.700 186.400 432.300 227.600 ;
        RECT 433.300 226.400 433.900 241.600 ;
        RECT 438.100 240.400 438.700 271.600 ;
        RECT 441.200 269.600 442.000 270.400 ;
        RECT 442.800 269.600 443.600 270.400 ;
        RECT 439.600 267.600 440.400 268.400 ;
        RECT 441.300 242.400 441.900 269.600 ;
        RECT 444.500 262.400 445.100 271.600 ;
        RECT 446.100 266.400 446.700 283.600 ;
        RECT 454.100 278.400 454.700 285.600 ;
        RECT 462.000 284.200 462.800 297.800 ;
        RECT 463.600 284.200 464.400 297.800 ;
        RECT 465.200 284.200 466.000 297.800 ;
        RECT 466.800 286.200 467.600 297.800 ;
        RECT 468.500 296.400 469.100 305.600 ;
        RECT 481.200 303.600 482.000 304.400 ;
        RECT 468.400 295.600 469.200 296.400 ;
        RECT 470.000 286.200 470.800 297.800 ;
        RECT 471.600 293.600 472.400 294.400 ;
        RECT 471.700 292.400 472.300 293.600 ;
        RECT 471.600 291.600 472.400 292.400 ;
        RECT 473.200 286.200 474.000 297.800 ;
        RECT 474.800 284.200 475.600 297.800 ;
        RECT 476.400 284.200 477.200 297.800 ;
        RECT 479.600 291.600 480.400 292.400 ;
        RECT 454.000 277.600 454.800 278.400 ;
        RECT 462.000 269.600 462.800 270.400 ;
        RECT 449.200 267.600 450.000 268.400 ;
        RECT 446.000 265.600 446.800 266.400 ;
        RECT 450.800 265.600 451.600 266.400 ;
        RECT 447.600 263.600 448.400 264.400 ;
        RECT 444.400 261.600 445.200 262.400 ;
        RECT 447.700 260.400 448.300 263.600 ;
        RECT 447.600 259.600 448.400 260.400 ;
        RECT 442.800 251.600 443.600 252.400 ;
        RECT 444.400 244.200 445.200 257.800 ;
        RECT 446.000 244.200 446.800 257.800 ;
        RECT 447.600 244.200 448.400 257.800 ;
        RECT 449.200 246.200 450.000 257.800 ;
        RECT 450.900 256.400 451.500 265.600 ;
        RECT 450.800 255.600 451.600 256.400 ;
        RECT 450.800 245.600 451.600 246.400 ;
        RECT 452.400 246.200 453.200 257.800 ;
        RECT 454.000 253.600 454.800 254.400 ;
        RECT 441.200 241.600 442.000 242.400 ;
        RECT 438.000 239.600 438.800 240.400 ;
        RECT 441.200 239.600 442.000 240.400 ;
        RECT 441.300 238.400 441.900 239.600 ;
        RECT 441.200 237.600 442.000 238.400 ;
        RECT 444.400 237.600 445.200 238.400 ;
        RECT 439.600 233.600 440.400 234.400 ;
        RECT 441.200 231.600 442.000 232.400 ;
        RECT 434.800 229.600 435.600 230.400 ;
        RECT 436.400 229.600 437.200 230.400 ;
        RECT 441.200 229.600 442.000 230.400 ;
        RECT 434.900 228.400 435.500 229.600 ;
        RECT 434.800 227.600 435.600 228.400 ;
        RECT 433.200 225.600 434.000 226.400 ;
        RECT 438.000 225.600 438.800 226.400 ;
        RECT 433.300 222.400 433.900 225.600 ;
        RECT 438.100 224.400 438.700 225.600 ;
        RECT 438.000 223.600 438.800 224.400 ;
        RECT 433.200 221.600 434.000 222.400 ;
        RECT 433.300 218.400 433.900 221.600 ;
        RECT 433.200 217.600 434.000 218.400 ;
        RECT 434.800 217.600 435.600 218.400 ;
        RECT 434.900 214.400 435.500 217.600 ;
        RECT 438.100 216.400 438.700 223.600 ;
        RECT 441.300 216.400 441.900 229.600 ;
        RECT 444.500 228.300 445.100 237.600 ;
        RECT 446.000 231.600 446.800 232.400 ;
        RECT 449.200 231.600 450.000 232.400 ;
        RECT 446.000 228.300 446.800 228.400 ;
        RECT 444.500 227.700 446.800 228.300 ;
        RECT 444.500 216.400 445.100 227.700 ;
        RECT 446.000 227.600 446.800 227.700 ;
        RECT 449.300 218.400 449.900 231.600 ;
        RECT 450.900 228.400 451.500 245.600 ;
        RECT 454.100 230.400 454.700 253.600 ;
        RECT 455.600 246.200 456.400 257.800 ;
        RECT 457.200 244.200 458.000 257.800 ;
        RECT 458.800 244.200 459.600 257.800 ;
        RECT 462.100 252.400 462.700 269.600 ;
        RECT 463.600 264.200 464.400 277.800 ;
        RECT 465.200 264.200 466.000 277.800 ;
        RECT 466.800 264.200 467.600 277.800 ;
        RECT 468.400 264.200 469.200 275.800 ;
        RECT 470.000 265.600 470.800 266.400 ;
        RECT 471.600 264.200 472.400 275.800 ;
        RECT 473.200 269.600 474.000 270.400 ;
        RECT 473.300 268.400 473.900 269.600 ;
        RECT 473.200 267.600 474.000 268.400 ;
        RECT 474.800 264.200 475.600 275.800 ;
        RECT 476.400 264.200 477.200 277.800 ;
        RECT 478.000 264.200 478.800 277.800 ;
        RECT 479.700 270.400 480.300 291.600 ;
        RECT 479.600 269.600 480.400 270.400 ;
        RECT 479.600 267.600 480.400 268.400 ;
        RECT 465.200 261.600 466.000 262.400 ;
        RECT 466.800 261.600 467.600 262.400 ;
        RECT 462.000 251.600 462.800 252.400 ;
        RECT 465.300 238.400 465.900 261.600 ;
        RECT 466.900 248.300 467.500 261.600 ;
        RECT 473.200 257.600 474.000 258.400 ;
        RECT 468.400 255.600 469.200 256.400 ;
        RECT 468.500 250.400 469.100 255.600 ;
        RECT 471.600 253.600 472.400 254.400 ;
        RECT 471.700 252.400 472.300 253.600 ;
        RECT 473.300 252.400 473.900 257.600 ;
        RECT 478.000 255.600 478.800 256.400 ;
        RECT 476.400 253.600 477.200 254.400 ;
        RECT 470.000 251.600 470.800 252.400 ;
        RECT 471.600 251.600 472.400 252.400 ;
        RECT 473.200 251.600 474.000 252.400 ;
        RECT 474.800 251.600 475.600 252.400 ;
        RECT 470.100 250.400 470.700 251.600 ;
        RECT 474.900 250.400 475.500 251.600 ;
        RECT 468.400 249.600 469.200 250.400 ;
        RECT 470.000 249.600 470.800 250.400 ;
        RECT 474.800 249.600 475.600 250.400 ;
        RECT 466.900 247.700 469.100 248.300 ;
        RECT 455.600 237.600 456.400 238.400 ;
        RECT 458.800 237.600 459.600 238.400 ;
        RECT 465.200 237.600 466.000 238.400 ;
        RECT 455.700 232.400 456.300 237.600 ;
        RECT 460.400 233.600 461.200 234.400 ;
        RECT 466.800 233.600 467.600 234.400 ;
        RECT 455.600 231.600 456.400 232.400 ;
        RECT 457.200 231.600 458.000 232.400 ;
        RECT 463.600 231.600 464.400 232.400 ;
        RECT 465.200 231.600 466.000 232.400 ;
        RECT 465.300 230.400 465.900 231.600 ;
        RECT 452.400 229.600 453.200 230.400 ;
        RECT 454.000 229.600 454.800 230.400 ;
        RECT 455.600 229.600 456.400 230.400 ;
        RECT 458.800 230.300 459.600 230.400 ;
        RECT 458.800 229.700 461.100 230.300 ;
        RECT 458.800 229.600 459.600 229.700 ;
        RECT 450.800 227.600 451.600 228.400 ;
        RECT 452.500 222.400 453.100 229.600 ;
        RECT 452.400 221.600 453.200 222.400 ;
        RECT 449.200 217.600 450.000 218.400 ;
        RECT 436.400 215.600 437.200 216.400 ;
        RECT 438.000 215.600 438.800 216.400 ;
        RECT 441.200 215.600 442.000 216.400 ;
        RECT 444.400 215.600 445.200 216.400 ;
        RECT 446.000 215.600 446.800 216.400 ;
        RECT 447.600 215.600 448.400 216.400 ;
        RECT 434.800 213.600 435.600 214.400 ;
        RECT 436.500 212.400 437.100 215.600 ;
        RECT 434.800 211.600 435.600 212.400 ;
        RECT 436.400 211.600 437.200 212.400 ;
        RECT 441.200 211.600 442.000 212.400 ;
        RECT 442.800 211.600 443.600 212.400 ;
        RECT 433.200 191.600 434.000 192.400 ;
        RECT 434.900 190.400 435.500 211.600 ;
        RECT 436.500 194.400 437.100 211.600 ;
        RECT 441.300 204.400 441.900 211.600 ;
        RECT 441.200 203.600 442.000 204.400 ;
        RECT 436.400 193.600 437.200 194.400 ;
        RECT 436.400 191.600 437.200 192.400 ;
        RECT 436.500 190.400 437.100 191.600 ;
        RECT 441.300 190.400 441.900 203.600 ;
        RECT 442.900 200.400 443.500 211.600 ;
        RECT 446.100 208.400 446.700 215.600 ;
        RECT 447.700 214.400 448.300 215.600 ;
        RECT 455.700 214.400 456.300 229.600 ;
        RECT 460.500 228.400 461.100 229.700 ;
        RECT 465.200 229.600 466.000 230.400 ;
        RECT 458.800 227.600 459.600 228.400 ;
        RECT 460.400 227.600 461.200 228.400 ;
        RECT 457.200 225.600 458.000 226.400 ;
        RECT 447.600 213.600 448.400 214.400 ;
        RECT 452.400 213.600 453.200 214.400 ;
        RECT 454.000 213.600 454.800 214.400 ;
        RECT 455.600 213.600 456.400 214.400 ;
        RECT 452.500 212.400 453.100 213.600 ;
        RECT 449.200 211.600 450.000 212.400 ;
        RECT 452.400 211.600 453.200 212.400 ;
        RECT 449.300 210.400 449.900 211.600 ;
        RECT 447.600 209.600 448.400 210.400 ;
        RECT 449.200 209.600 450.000 210.400 ;
        RECT 444.400 207.600 445.200 208.400 ;
        RECT 446.000 207.600 446.800 208.400 ;
        RECT 442.800 199.600 443.600 200.400 ;
        RECT 447.700 198.400 448.300 209.600 ;
        RECT 449.200 207.600 450.000 208.400 ;
        RECT 447.600 197.600 448.400 198.400 ;
        RECT 446.000 193.600 446.800 194.400 ;
        RECT 434.800 189.600 435.600 190.400 ;
        RECT 436.400 189.600 437.200 190.400 ;
        RECT 441.200 189.600 442.000 190.400 ;
        RECT 433.200 187.600 434.000 188.400 ;
        RECT 433.300 186.400 433.900 187.600 ;
        RECT 431.600 185.600 432.400 186.400 ;
        RECT 433.200 185.600 434.000 186.400 ;
        RECT 431.700 180.400 432.300 185.600 ;
        RECT 434.800 183.600 435.600 184.400 ;
        RECT 439.600 184.300 440.400 184.400 ;
        RECT 438.100 183.700 440.400 184.300 ;
        RECT 431.600 179.600 432.400 180.400 ;
        RECT 428.400 164.200 429.200 177.800 ;
        RECT 430.000 164.200 430.800 177.800 ;
        RECT 431.600 164.200 432.400 177.800 ;
        RECT 433.200 166.200 434.000 177.800 ;
        RECT 434.900 176.400 435.500 183.600 ;
        RECT 434.800 175.600 435.600 176.400 ;
        RECT 433.200 155.600 434.000 156.400 ;
        RECT 420.500 151.700 422.700 152.300 ;
        RECT 406.000 149.600 406.800 150.400 ;
        RECT 407.600 149.600 408.400 150.400 ;
        RECT 410.800 149.600 411.600 150.400 ;
        RECT 412.400 149.600 413.200 150.400 ;
        RECT 412.500 146.400 413.100 149.600 ;
        RECT 412.400 145.600 413.200 146.400 ;
        RECT 404.400 143.600 405.200 144.400 ;
        RECT 402.800 123.600 403.600 124.400 ;
        RECT 404.500 112.400 405.100 143.600 ;
        RECT 414.100 142.300 414.700 151.600 ;
        RECT 418.800 149.600 419.600 150.400 ;
        RECT 420.400 149.600 421.200 150.400 ;
        RECT 418.900 148.400 419.500 149.600 ;
        RECT 418.800 147.600 419.600 148.400 ;
        RECT 415.600 145.600 416.400 146.400 ;
        RECT 415.700 144.400 416.300 145.600 ;
        RECT 420.500 144.400 421.100 149.600 ;
        RECT 415.600 143.600 416.400 144.400 ;
        RECT 417.200 143.600 418.000 144.400 ;
        RECT 420.400 143.600 421.200 144.400 ;
        RECT 414.100 141.700 416.300 142.300 ;
        RECT 406.000 124.200 406.800 137.800 ;
        RECT 407.600 124.200 408.400 137.800 ;
        RECT 409.200 124.200 410.000 137.800 ;
        RECT 410.800 126.200 411.600 137.800 ;
        RECT 412.400 135.600 413.200 136.400 ;
        RECT 412.400 133.600 413.200 134.400 ;
        RECT 407.600 121.600 408.400 122.400 ;
        RECT 404.400 111.600 405.200 112.400 ;
        RECT 407.700 110.400 408.300 121.600 ;
        RECT 412.500 110.400 413.100 133.600 ;
        RECT 414.000 126.200 414.800 137.800 ;
        RECT 415.700 134.400 416.300 141.700 ;
        RECT 415.600 133.600 416.400 134.400 ;
        RECT 417.200 126.200 418.000 137.800 ;
        RECT 418.800 124.200 419.600 137.800 ;
        RECT 420.400 124.200 421.200 137.800 ;
        RECT 422.100 134.400 422.700 151.700 ;
        RECT 423.600 151.600 424.400 152.400 ;
        RECT 425.200 149.600 426.000 150.400 ;
        RECT 426.800 147.600 427.600 148.400 ;
        RECT 426.900 136.400 427.500 147.600 ;
        RECT 426.800 135.600 427.600 136.400 ;
        RECT 422.000 133.600 422.800 134.400 ;
        RECT 425.200 131.600 426.000 132.400 ;
        RECT 425.300 126.400 425.900 131.600 ;
        RECT 425.200 125.600 426.000 126.400 ;
        RECT 420.400 119.600 421.200 120.400 ;
        RECT 431.600 119.600 432.400 120.400 ;
        RECT 415.600 115.600 416.400 116.400 ;
        RECT 414.000 111.600 414.800 112.400 ;
        RECT 407.600 109.600 408.400 110.400 ;
        RECT 412.400 109.600 413.200 110.400 ;
        RECT 415.700 110.300 416.300 115.600 ;
        RECT 420.500 112.400 421.100 119.600 ;
        RECT 417.200 112.300 418.000 112.400 ;
        RECT 417.200 111.700 419.500 112.300 ;
        RECT 417.200 111.600 418.000 111.700 ;
        RECT 418.900 110.400 419.500 111.700 ;
        RECT 420.400 111.600 421.200 112.400 ;
        RECT 431.700 110.400 432.300 119.600 ;
        RECT 433.300 110.400 433.900 155.600 ;
        RECT 434.900 154.300 435.500 175.600 ;
        RECT 436.400 166.200 437.200 177.800 ;
        RECT 438.100 174.400 438.700 183.700 ;
        RECT 439.600 183.600 440.400 183.700 ;
        RECT 446.100 178.400 446.700 193.600 ;
        RECT 447.600 189.600 448.400 190.400 ;
        RECT 447.700 188.400 448.300 189.600 ;
        RECT 447.600 187.600 448.400 188.400 ;
        RECT 447.600 181.600 448.400 182.400 ;
        RECT 438.000 173.600 438.800 174.400 ;
        RECT 439.600 166.200 440.400 177.800 ;
        RECT 441.200 164.200 442.000 177.800 ;
        RECT 442.800 164.200 443.600 177.800 ;
        RECT 446.000 177.600 446.800 178.400 ;
        RECT 447.700 172.400 448.300 181.600 ;
        RECT 452.500 172.400 453.100 211.600 ;
        RECT 454.000 183.600 454.800 184.400 ;
        RECT 454.100 182.400 454.700 183.600 ;
        RECT 454.000 181.600 454.800 182.400 ;
        RECT 457.300 182.300 457.900 225.600 ;
        RECT 458.900 214.400 459.500 227.600 ;
        RECT 468.500 222.300 469.100 247.700 ;
        RECT 478.100 244.400 478.700 255.600 ;
        RECT 478.000 243.600 478.800 244.400 ;
        RECT 476.400 231.600 477.200 232.400 ;
        RECT 478.000 231.600 478.800 232.400 ;
        RECT 478.100 230.400 478.700 231.600 ;
        RECT 479.700 230.400 480.300 267.600 ;
        RECT 481.300 266.400 481.900 303.600 ;
        RECT 487.700 298.400 488.300 343.600 ;
        RECT 497.300 338.300 497.900 349.600 ;
        RECT 495.700 337.700 497.900 338.300 ;
        RECT 494.000 329.600 494.800 330.400 ;
        RECT 490.800 323.600 491.600 324.400 ;
        RECT 490.900 304.400 491.500 323.600 ;
        RECT 495.700 318.400 496.300 337.700 ;
        RECT 497.200 331.600 498.000 332.400 ;
        RECT 497.200 329.600 498.000 330.400 ;
        RECT 495.600 317.600 496.400 318.400 ;
        RECT 495.700 310.400 496.300 317.600 ;
        RECT 495.600 309.600 496.400 310.400 ;
        RECT 497.300 306.400 497.900 329.600 ;
        RECT 498.900 322.400 499.500 349.600 ;
        RECT 502.100 344.400 502.700 373.600 ;
        RECT 505.200 369.600 506.000 370.400 ;
        RECT 503.600 363.600 504.400 364.400 ;
        RECT 503.700 360.400 504.300 363.600 ;
        RECT 503.600 359.600 504.400 360.400 ;
        RECT 505.300 358.400 505.900 369.600 ;
        RECT 506.800 367.600 507.600 368.400 ;
        RECT 508.500 358.400 509.100 373.600 ;
        RECT 521.200 371.600 522.000 372.400 ;
        RECT 510.000 369.600 510.800 370.400 ;
        RECT 513.200 364.300 514.000 364.400 ;
        RECT 513.200 363.700 515.500 364.300 ;
        RECT 522.800 364.200 523.600 377.800 ;
        RECT 524.400 364.200 525.200 377.800 ;
        RECT 526.000 364.200 526.800 377.800 ;
        RECT 527.600 366.200 528.400 377.800 ;
        RECT 529.200 375.600 530.000 376.400 ;
        RECT 529.300 372.400 529.900 375.600 ;
        RECT 529.200 371.600 530.000 372.400 ;
        RECT 530.800 366.200 531.600 377.800 ;
        RECT 532.400 373.600 533.200 374.400 ;
        RECT 532.400 371.600 533.200 372.400 ;
        RECT 513.200 363.600 514.000 363.700 ;
        RECT 505.200 357.600 506.000 358.400 ;
        RECT 508.400 357.600 509.200 358.400 ;
        RECT 508.400 351.600 509.200 352.400 ;
        RECT 503.600 349.600 504.400 350.400 ;
        RECT 502.000 343.600 502.800 344.400 ;
        RECT 503.700 338.400 504.300 349.600 ;
        RECT 508.500 346.400 509.100 351.600 ;
        RECT 513.200 349.600 514.000 350.400 ;
        RECT 511.600 347.600 512.400 348.400 ;
        RECT 506.800 345.600 507.600 346.400 ;
        RECT 508.400 345.600 509.200 346.400 ;
        RECT 506.900 344.400 507.500 345.600 ;
        RECT 506.800 343.600 507.600 344.400 ;
        RECT 503.600 337.600 504.400 338.400 ;
        RECT 506.800 337.600 507.600 338.400 ;
        RECT 506.900 336.400 507.500 337.600 ;
        RECT 503.600 335.600 504.400 336.400 ;
        RECT 506.800 335.600 507.600 336.400 ;
        RECT 503.700 334.400 504.300 335.600 ;
        RECT 503.600 333.600 504.400 334.400 ;
        RECT 508.400 333.600 509.200 334.400 ;
        RECT 502.000 331.600 502.800 332.400 ;
        RECT 502.100 330.400 502.700 331.600 ;
        RECT 502.000 329.600 502.800 330.400 ;
        RECT 503.700 328.400 504.300 333.600 ;
        RECT 510.000 331.600 510.800 332.400 ;
        RECT 503.600 327.600 504.400 328.400 ;
        RECT 506.800 327.600 507.600 328.400 ;
        RECT 505.200 323.600 506.000 324.400 ;
        RECT 498.800 321.600 499.600 322.400 ;
        RECT 498.800 319.600 499.600 320.400 ;
        RECT 498.900 318.400 499.500 319.600 ;
        RECT 498.800 317.600 499.600 318.400 ;
        RECT 503.600 309.600 504.400 310.400 ;
        RECT 503.700 306.400 504.300 309.600 ;
        RECT 494.000 305.600 494.800 306.400 ;
        RECT 497.200 305.600 498.000 306.400 ;
        RECT 503.600 305.600 504.400 306.400 ;
        RECT 490.800 303.600 491.600 304.400 ;
        RECT 487.600 297.600 488.400 298.400 ;
        RECT 494.000 297.600 494.800 298.400 ;
        RECT 486.000 295.600 486.800 296.400 ;
        RECT 492.400 295.600 493.200 296.400 ;
        RECT 486.100 272.400 486.700 295.600 ;
        RECT 492.500 294.400 493.100 295.600 ;
        RECT 489.200 293.600 490.000 294.400 ;
        RECT 492.400 293.600 493.200 294.400 ;
        RECT 494.100 292.400 494.700 297.600 ;
        RECT 490.800 291.600 491.600 292.400 ;
        RECT 494.000 291.600 494.800 292.400 ;
        RECT 495.600 291.600 496.400 292.400 ;
        RECT 489.200 277.600 490.000 278.400 ;
        RECT 486.000 271.600 486.800 272.400 ;
        RECT 482.800 269.600 483.600 270.400 ;
        RECT 481.200 265.600 482.000 266.400 ;
        RECT 481.200 263.600 482.000 264.400 ;
        RECT 473.200 229.600 474.000 230.400 ;
        RECT 478.000 229.600 478.800 230.400 ;
        RECT 479.600 229.600 480.400 230.400 ;
        RECT 473.300 228.400 473.900 229.600 ;
        RECT 470.000 227.600 470.800 228.400 ;
        RECT 473.200 227.600 474.000 228.400 ;
        RECT 470.000 225.600 470.800 226.400 ;
        RECT 474.800 225.600 475.600 226.400 ;
        RECT 470.100 224.400 470.700 225.600 ;
        RECT 474.900 224.400 475.500 225.600 ;
        RECT 470.000 223.600 470.800 224.400 ;
        RECT 473.200 223.600 474.000 224.400 ;
        RECT 474.800 223.600 475.600 224.400 ;
        RECT 468.500 221.700 470.700 222.300 ;
        RECT 458.800 213.600 459.600 214.400 ;
        RECT 462.000 213.600 462.800 214.400 ;
        RECT 460.400 211.600 461.200 212.400 ;
        RECT 463.600 211.600 464.400 212.400 ;
        RECT 465.200 211.600 466.000 212.400 ;
        RECT 460.500 202.400 461.100 211.600 ;
        RECT 468.400 203.600 469.200 204.400 ;
        RECT 460.400 201.600 461.200 202.400 ;
        RECT 465.200 199.600 466.000 200.400 ;
        RECT 465.300 198.400 465.900 199.600 ;
        RECT 468.500 198.400 469.100 203.600 ;
        RECT 470.100 198.400 470.700 221.700 ;
        RECT 473.300 214.400 473.900 223.600 ;
        RECT 473.200 213.600 474.000 214.400 ;
        RECT 478.100 212.400 478.700 229.600 ;
        RECT 479.600 227.600 480.400 228.400 ;
        RECT 479.700 226.400 480.300 227.600 ;
        RECT 479.600 225.600 480.400 226.400 ;
        RECT 481.300 218.400 481.900 263.600 ;
        RECT 482.900 252.400 483.500 269.600 ;
        RECT 490.900 266.400 491.500 291.600 ;
        RECT 497.300 278.400 497.900 305.600 ;
        RECT 505.300 302.400 505.900 323.600 ;
        RECT 506.900 306.400 507.500 327.600 ;
        RECT 511.700 320.400 512.300 347.600 ;
        RECT 514.900 338.400 515.500 363.700 ;
        RECT 522.800 353.600 523.600 354.400 ;
        RECT 516.400 343.600 517.200 344.400 ;
        RECT 516.500 342.400 517.100 343.600 ;
        RECT 516.400 341.600 517.200 342.400 ;
        RECT 514.800 337.600 515.600 338.400 ;
        RECT 514.900 334.400 515.500 337.600 ;
        RECT 516.500 336.400 517.100 341.600 ;
        RECT 522.900 338.400 523.500 353.600 ;
        RECT 526.000 344.200 526.800 357.800 ;
        RECT 527.600 344.200 528.400 357.800 ;
        RECT 529.200 344.200 530.000 357.800 ;
        RECT 530.800 344.200 531.600 355.800 ;
        RECT 532.500 346.400 533.100 371.600 ;
        RECT 534.000 366.200 534.800 377.800 ;
        RECT 535.600 364.200 536.400 377.800 ;
        RECT 537.200 364.200 538.000 377.800 ;
        RECT 548.400 375.600 549.200 376.400 ;
        RECT 542.000 371.600 542.800 372.400 ;
        RECT 532.400 345.600 533.200 346.400 ;
        RECT 524.400 341.600 525.200 342.400 ;
        RECT 522.800 337.600 523.600 338.400 ;
        RECT 524.500 336.400 525.100 341.600 ;
        RECT 516.400 335.600 517.200 336.400 ;
        RECT 521.200 335.600 522.000 336.400 ;
        RECT 524.400 335.600 525.200 336.400 ;
        RECT 514.800 333.600 515.600 334.400 ;
        RECT 516.400 333.600 517.200 334.400 ;
        RECT 516.500 332.400 517.100 333.600 ;
        RECT 514.800 331.600 515.600 332.400 ;
        RECT 516.400 331.600 517.200 332.400 ;
        RECT 518.000 331.600 518.800 332.400 ;
        RECT 521.200 331.600 522.000 332.400 ;
        RECT 524.400 331.600 525.200 332.400 ;
        RECT 530.800 331.600 531.600 332.400 ;
        RECT 513.200 329.600 514.000 330.400 ;
        RECT 513.300 328.400 513.900 329.600 ;
        RECT 513.200 327.600 514.000 328.400 ;
        RECT 511.600 319.600 512.400 320.400 ;
        RECT 514.900 312.400 515.500 331.600 ;
        RECT 514.800 311.600 515.600 312.400 ;
        RECT 510.000 309.600 510.800 310.400 ;
        RECT 511.600 309.600 512.400 310.400 ;
        RECT 508.400 307.600 509.200 308.400 ;
        RECT 511.700 308.300 512.300 309.600 ;
        RECT 510.100 307.700 512.300 308.300 ;
        RECT 506.800 305.600 507.600 306.400 ;
        RECT 506.800 303.600 507.600 304.400 ;
        RECT 505.200 301.600 506.000 302.400 ;
        RECT 500.400 299.600 501.200 300.400 ;
        RECT 500.500 298.400 501.100 299.600 ;
        RECT 500.400 297.600 501.200 298.400 ;
        RECT 502.000 297.600 502.800 298.400 ;
        RECT 498.800 295.600 499.600 296.400 ;
        RECT 498.900 294.400 499.500 295.600 ;
        RECT 502.100 294.400 502.700 297.600 ;
        RECT 503.600 295.600 504.400 296.400 ;
        RECT 503.700 294.400 504.300 295.600 ;
        RECT 498.800 293.600 499.600 294.400 ;
        RECT 502.000 293.600 502.800 294.400 ;
        RECT 503.600 293.600 504.400 294.400 ;
        RECT 506.900 292.400 507.500 303.600 ;
        RECT 510.100 298.400 510.700 307.700 ;
        RECT 513.200 307.600 514.000 308.400 ;
        RECT 511.600 301.600 512.400 302.400 ;
        RECT 510.000 297.600 510.800 298.400 ;
        RECT 511.700 294.400 512.300 301.600 ;
        RECT 513.300 296.400 513.900 307.600 ;
        RECT 516.400 305.600 517.200 306.400 ;
        RECT 514.800 303.600 515.600 304.400 ;
        RECT 513.200 295.600 514.000 296.400 ;
        RECT 511.600 293.600 512.400 294.400 ;
        RECT 498.800 291.600 499.600 292.400 ;
        RECT 506.800 291.600 507.600 292.400 ;
        RECT 508.400 290.300 509.200 290.400 ;
        RECT 506.900 289.700 509.200 290.300 ;
        RECT 506.900 288.400 507.500 289.700 ;
        RECT 508.400 289.600 509.200 289.700 ;
        RECT 506.800 287.600 507.600 288.400 ;
        RECT 497.200 277.600 498.000 278.400 ;
        RECT 497.200 269.600 498.000 270.400 ;
        RECT 490.800 265.600 491.600 266.400 ;
        RECT 490.900 264.400 491.500 265.600 ;
        RECT 490.800 263.600 491.600 264.400 ;
        RECT 495.600 263.600 496.400 264.400 ;
        RECT 498.800 264.200 499.600 277.800 ;
        RECT 500.400 264.200 501.200 277.800 ;
        RECT 502.000 264.200 502.800 277.800 ;
        RECT 503.600 264.200 504.400 275.800 ;
        RECT 505.200 265.600 506.000 266.400 ;
        RECT 505.300 264.400 505.900 265.600 ;
        RECT 505.200 263.600 506.000 264.400 ;
        RECT 506.800 264.200 507.600 275.800 ;
        RECT 508.400 267.600 509.200 268.400 ;
        RECT 510.000 264.200 510.800 275.800 ;
        RECT 511.600 264.200 512.400 277.800 ;
        RECT 513.200 264.200 514.000 277.800 ;
        RECT 514.900 268.400 515.500 303.600 ;
        RECT 516.500 294.400 517.100 305.600 ;
        RECT 518.100 296.400 518.700 331.600 ;
        RECT 521.300 330.400 521.900 331.600 ;
        RECT 519.600 329.600 520.400 330.400 ;
        RECT 521.200 329.600 522.000 330.400 ;
        RECT 519.700 310.400 520.300 329.600 ;
        RECT 519.600 309.600 520.400 310.400 ;
        RECT 521.300 308.400 521.900 329.600 ;
        RECT 524.500 318.400 525.100 331.600 ;
        RECT 524.400 317.600 525.200 318.400 ;
        RECT 530.800 309.600 531.600 310.400 ;
        RECT 521.200 307.600 522.000 308.400 ;
        RECT 526.000 307.600 526.800 308.400 ;
        RECT 529.200 307.600 530.000 308.400 ;
        RECT 532.500 308.300 533.100 345.600 ;
        RECT 534.000 344.200 534.800 355.800 ;
        RECT 535.600 347.600 536.400 348.400 ;
        RECT 535.700 342.300 536.300 347.600 ;
        RECT 537.200 344.200 538.000 355.800 ;
        RECT 538.800 344.200 539.600 357.800 ;
        RECT 540.400 344.200 541.200 357.800 ;
        RECT 542.100 350.400 542.700 371.600 ;
        RECT 546.800 363.600 547.600 364.400 ;
        RECT 542.000 349.600 542.800 350.400 ;
        RECT 534.100 341.700 536.300 342.300 ;
        RECT 534.100 338.400 534.700 341.700 ;
        RECT 534.000 337.600 534.800 338.400 ;
        RECT 537.200 337.600 538.000 338.400 ;
        RECT 535.600 333.600 536.400 334.400 ;
        RECT 534.000 329.600 534.800 330.400 ;
        RECT 534.000 311.600 534.800 312.400 ;
        RECT 535.700 310.300 536.300 333.600 ;
        RECT 537.300 332.400 537.900 337.600 ;
        RECT 543.600 335.600 544.400 336.400 ;
        RECT 537.200 331.600 538.000 332.400 ;
        RECT 537.200 329.600 538.000 330.400 ;
        RECT 540.400 327.600 541.200 328.400 ;
        RECT 540.500 312.400 541.100 327.600 ;
        RECT 537.200 311.600 538.000 312.400 ;
        RECT 540.400 311.600 541.200 312.400 ;
        RECT 537.200 310.300 538.000 310.400 ;
        RECT 535.700 309.700 538.000 310.300 ;
        RECT 537.200 309.600 538.000 309.700 ;
        RECT 530.900 307.700 533.100 308.300 ;
        RECT 526.100 306.400 526.700 307.600 ;
        RECT 524.400 305.600 525.200 306.400 ;
        RECT 526.000 305.600 526.800 306.400 ;
        RECT 524.500 300.400 525.100 305.600 ;
        RECT 524.400 299.600 525.200 300.400 ;
        RECT 518.000 295.600 518.800 296.400 ;
        RECT 516.400 293.600 517.200 294.400 ;
        RECT 514.800 267.600 515.600 268.400 ;
        RECT 482.800 251.600 483.600 252.400 ;
        RECT 482.800 243.600 483.600 244.400 ;
        RECT 487.600 244.200 488.400 257.800 ;
        RECT 489.200 244.200 490.000 257.800 ;
        RECT 490.800 246.200 491.600 257.800 ;
        RECT 492.400 253.600 493.200 254.400 ;
        RECT 494.000 246.200 494.800 257.800 ;
        RECT 495.700 256.400 496.300 263.600 ;
        RECT 495.600 255.600 496.400 256.400 ;
        RECT 482.900 226.300 483.500 243.600 ;
        RECT 487.600 231.600 488.400 232.400 ;
        RECT 489.200 231.600 490.000 232.400 ;
        RECT 484.400 229.600 485.200 230.400 ;
        RECT 484.400 226.300 485.200 226.400 ;
        RECT 482.900 225.700 485.200 226.300 ;
        RECT 484.400 225.600 485.200 225.700 ;
        RECT 481.200 217.600 482.000 218.400 ;
        RECT 471.600 211.600 472.400 212.400 ;
        RECT 474.800 211.600 475.600 212.400 ;
        RECT 476.400 211.600 477.200 212.400 ;
        RECT 478.000 211.600 478.800 212.400 ;
        RECT 474.900 210.400 475.500 211.600 ;
        RECT 474.800 209.600 475.600 210.400 ;
        RECT 465.200 197.600 466.000 198.400 ;
        RECT 468.400 197.600 469.200 198.400 ;
        RECT 470.000 197.600 470.800 198.400 ;
        RECT 458.800 195.600 459.600 196.400 ;
        RECT 458.900 190.400 459.500 195.600 ;
        RECT 460.400 193.600 461.200 194.400 ;
        RECT 463.600 193.600 464.400 194.400 ;
        RECT 460.400 191.600 461.200 192.400 ;
        RECT 462.000 191.600 462.800 192.400 ;
        RECT 458.800 189.600 459.600 190.400 ;
        RECT 458.800 187.600 459.600 188.400 ;
        RECT 455.700 181.700 457.900 182.300 ;
        RECT 455.700 176.400 456.300 181.700 ;
        RECT 460.500 176.400 461.100 191.600 ;
        RECT 462.100 188.400 462.700 191.600 ;
        RECT 462.000 187.600 462.800 188.400 ;
        RECT 463.700 178.400 464.300 193.600 ;
        RECT 465.200 189.600 466.000 190.400 ;
        RECT 466.800 189.600 467.600 190.400 ;
        RECT 466.900 188.400 467.500 189.600 ;
        RECT 474.900 188.400 475.500 209.600 ;
        RECT 466.800 187.600 467.600 188.400 ;
        RECT 474.800 187.600 475.600 188.400 ;
        RECT 474.900 178.400 475.500 187.600 ;
        RECT 476.500 180.400 477.100 211.600 ;
        RECT 478.000 209.600 478.800 210.400 ;
        RECT 478.100 206.400 478.700 209.600 ;
        RECT 489.300 206.400 489.900 231.600 ;
        RECT 495.700 226.400 496.300 255.600 ;
        RECT 497.200 246.200 498.000 257.800 ;
        RECT 498.800 244.200 499.600 257.800 ;
        RECT 500.400 244.200 501.200 257.800 ;
        RECT 502.000 244.200 502.800 257.800 ;
        RECT 511.600 251.600 512.600 252.400 ;
        RECT 516.500 244.400 517.100 293.600 ;
        RECT 519.600 291.600 520.400 292.400 ;
        RECT 522.800 291.600 523.600 292.400 ;
        RECT 519.700 270.400 520.300 291.600 ;
        RECT 524.400 284.200 525.200 297.800 ;
        RECT 526.000 284.200 526.800 297.800 ;
        RECT 527.600 284.200 528.400 297.800 ;
        RECT 529.200 286.200 530.000 297.800 ;
        RECT 530.900 296.400 531.500 307.700 ;
        RECT 535.600 307.600 536.400 308.400 ;
        RECT 537.300 304.400 537.900 309.600 ;
        RECT 534.000 303.600 534.800 304.400 ;
        RECT 537.200 303.600 538.000 304.400 ;
        RECT 543.600 303.600 544.400 304.400 ;
        RECT 530.800 295.600 531.600 296.400 ;
        RECT 530.900 282.400 531.500 295.600 ;
        RECT 532.400 286.200 533.200 297.800 ;
        RECT 534.100 294.400 534.700 303.600 ;
        RECT 534.000 293.600 534.800 294.400 ;
        RECT 535.600 286.200 536.400 297.800 ;
        RECT 537.200 284.200 538.000 297.800 ;
        RECT 538.800 284.200 539.600 297.800 ;
        RECT 527.600 281.600 528.400 282.400 ;
        RECT 530.800 281.600 531.600 282.400 ;
        RECT 519.600 269.600 520.400 270.400 ;
        RECT 524.400 265.600 525.200 266.400 ;
        RECT 526.000 266.200 526.800 271.800 ;
        RECT 527.700 268.400 528.300 281.600 ;
        RECT 530.800 279.600 531.600 280.400 ;
        RECT 527.600 267.600 528.400 268.400 ;
        RECT 527.700 264.400 528.300 267.600 ;
        RECT 522.800 263.600 523.600 264.400 ;
        RECT 527.600 263.600 528.400 264.400 ;
        RECT 529.200 264.200 530.000 275.800 ;
        RECT 530.900 270.200 531.500 279.600 ;
        RECT 530.800 269.400 531.600 270.200 ;
        RECT 535.600 267.600 536.400 268.400 ;
        RECT 516.400 243.600 517.200 244.400 ;
        RECT 505.200 229.600 506.000 230.400 ;
        RECT 497.000 227.600 498.000 228.400 ;
        RECT 495.600 225.600 496.400 226.400 ;
        RECT 490.800 223.600 491.600 224.400 ;
        RECT 490.900 222.400 491.500 223.600 ;
        RECT 490.800 221.600 491.600 222.400 ;
        RECT 495.700 220.300 496.300 225.600 ;
        RECT 505.300 222.300 505.900 229.600 ;
        RECT 506.800 224.200 507.600 237.800 ;
        RECT 508.400 224.200 509.200 237.800 ;
        RECT 510.000 224.200 510.800 237.800 ;
        RECT 511.600 224.200 512.400 235.800 ;
        RECT 513.200 225.600 514.000 226.400 ;
        RECT 505.300 221.700 507.500 222.300 ;
        RECT 495.700 219.700 497.900 220.300 ;
        RECT 478.000 205.600 478.800 206.400 ;
        RECT 489.200 205.600 490.000 206.400 ;
        RECT 481.200 203.600 482.000 204.400 ;
        RECT 490.800 204.200 491.600 217.800 ;
        RECT 492.400 204.200 493.200 217.800 ;
        RECT 494.000 204.200 494.800 217.800 ;
        RECT 495.600 206.200 496.400 217.800 ;
        RECT 497.300 216.400 497.900 219.700 ;
        RECT 497.200 215.600 498.000 216.400 ;
        RECT 497.200 211.600 498.000 212.400 ;
        RECT 481.300 200.400 481.900 203.600 ;
        RECT 481.200 199.600 482.000 200.400 ;
        RECT 478.000 189.600 478.800 190.400 ;
        RECT 478.100 182.400 478.700 189.600 ;
        RECT 479.600 184.200 480.400 197.800 ;
        RECT 481.200 184.200 482.000 197.800 ;
        RECT 482.800 184.200 483.600 197.800 ;
        RECT 489.200 197.600 490.000 198.400 ;
        RECT 484.400 184.200 485.200 195.800 ;
        RECT 486.000 185.600 486.800 186.400 ;
        RECT 486.100 184.400 486.700 185.600 ;
        RECT 486.000 183.600 486.800 184.400 ;
        RECT 487.600 184.200 488.400 195.800 ;
        RECT 489.300 188.400 489.900 197.600 ;
        RECT 489.200 187.600 490.000 188.400 ;
        RECT 490.800 184.200 491.600 195.800 ;
        RECT 492.400 184.200 493.200 197.800 ;
        RECT 494.000 184.200 494.800 197.800 ;
        RECT 497.300 190.400 497.900 211.600 ;
        RECT 498.800 206.200 499.600 217.800 ;
        RECT 500.400 213.600 501.200 214.400 ;
        RECT 500.500 192.400 501.100 213.600 ;
        RECT 502.000 206.200 502.800 217.800 ;
        RECT 503.600 204.200 504.400 217.800 ;
        RECT 505.200 204.200 506.000 217.800 ;
        RECT 506.900 212.400 507.500 221.700 ;
        RECT 508.400 221.600 509.200 222.400 ;
        RECT 506.800 211.600 507.600 212.400 ;
        RECT 508.500 198.400 509.100 221.600 ;
        RECT 513.300 216.400 513.900 225.600 ;
        RECT 514.800 224.200 515.600 235.800 ;
        RECT 516.400 229.600 517.200 230.400 ;
        RECT 516.500 228.400 517.100 229.600 ;
        RECT 516.400 227.600 517.200 228.400 ;
        RECT 518.000 224.200 518.800 235.800 ;
        RECT 519.600 224.200 520.400 237.800 ;
        RECT 521.200 224.200 522.000 237.800 ;
        RECT 522.900 226.400 523.500 263.600 ;
        RECT 527.700 254.400 528.300 263.600 ;
        RECT 527.600 253.600 528.400 254.400 ;
        RECT 532.400 249.600 533.200 250.400 ;
        RECT 530.800 243.600 531.600 244.400 ;
        RECT 530.900 226.400 531.500 243.600 ;
        RECT 532.500 230.300 533.100 249.600 ;
        RECT 534.000 246.200 534.800 257.800 ;
        RECT 535.700 252.400 536.300 267.600 ;
        RECT 538.800 264.200 539.600 275.800 ;
        RECT 543.700 260.300 544.300 303.600 ;
        RECT 543.700 259.700 545.900 260.300 ;
        RECT 535.600 251.600 536.400 252.400 ;
        RECT 542.000 251.800 542.800 252.600 ;
        RECT 537.200 231.600 538.000 232.400 ;
        RECT 532.500 229.700 534.700 230.300 ;
        RECT 534.100 228.400 534.700 229.700 ;
        RECT 537.300 228.400 537.900 231.600 ;
        RECT 542.100 230.400 542.700 251.800 ;
        RECT 543.600 246.200 544.400 257.800 ;
        RECT 543.600 243.600 544.400 244.400 ;
        RECT 542.000 229.600 542.800 230.400 ;
        RECT 534.000 227.600 534.800 228.400 ;
        RECT 537.200 227.600 538.000 228.400 ;
        RECT 537.300 226.400 537.900 227.600 ;
        RECT 522.800 225.600 523.600 226.400 ;
        RECT 530.800 225.600 531.600 226.400 ;
        RECT 537.200 225.600 538.000 226.400 ;
        RECT 542.000 225.600 542.800 226.400 ;
        RECT 532.400 223.600 533.200 224.400 ;
        RECT 537.200 223.600 538.000 224.400 ;
        RECT 532.500 220.400 533.100 223.600 ;
        RECT 532.400 219.600 533.200 220.400 ;
        RECT 514.800 217.600 515.600 218.400 ;
        RECT 513.200 215.600 514.000 216.400 ;
        RECT 514.900 198.400 515.500 217.600 ;
        RECT 518.000 211.600 518.800 212.400 ;
        RECT 518.100 202.400 518.700 211.600 ;
        RECT 522.800 204.200 523.600 217.800 ;
        RECT 524.400 204.200 525.200 217.800 ;
        RECT 526.000 206.200 526.800 217.800 ;
        RECT 527.600 213.600 528.400 214.400 ;
        RECT 529.200 206.200 530.000 217.800 ;
        RECT 530.800 215.600 531.600 216.400 ;
        RECT 518.000 201.600 518.800 202.400 ;
        RECT 522.800 201.600 523.600 202.400 ;
        RECT 508.400 197.600 509.200 198.400 ;
        RECT 514.800 197.600 515.600 198.400 ;
        RECT 500.400 191.600 501.200 192.400 ;
        RECT 516.400 191.600 517.200 192.400 ;
        RECT 519.600 191.600 520.400 192.400 ;
        RECT 497.200 189.600 498.000 190.400 ;
        RECT 505.200 189.600 506.000 190.400 ;
        RECT 508.400 189.600 509.200 190.400 ;
        RECT 511.600 189.600 512.400 190.400 ;
        RECT 513.200 189.600 514.000 190.400 ;
        RECT 505.300 188.400 505.900 189.600 ;
        RECT 498.800 187.600 499.600 188.400 ;
        RECT 503.600 187.600 504.400 188.400 ;
        RECT 505.200 187.600 506.000 188.400 ;
        RECT 478.000 181.600 478.800 182.400 ;
        RECT 487.600 181.600 488.400 182.400 ;
        RECT 476.400 179.600 477.200 180.400 ;
        RECT 487.700 178.400 488.300 181.600 ;
        RECT 463.600 177.600 464.400 178.400 ;
        RECT 474.800 177.600 475.600 178.400 ;
        RECT 487.600 177.600 488.400 178.400 ;
        RECT 455.600 175.600 456.400 176.400 ;
        RECT 460.400 175.600 461.200 176.400 ;
        RECT 468.400 175.600 469.200 176.400 ;
        RECT 470.000 175.600 470.800 176.400 ;
        RECT 486.000 175.600 486.800 176.400 ;
        RECT 460.500 174.400 461.100 175.600 ;
        RECT 460.400 173.600 461.200 174.400 ;
        RECT 463.600 173.600 464.400 174.400 ;
        RECT 447.600 171.600 448.400 172.400 ;
        RECT 452.400 171.600 453.200 172.400 ;
        RECT 455.600 171.600 456.400 172.400 ;
        RECT 452.500 160.400 453.100 171.600 ;
        RECT 454.000 163.600 454.800 164.400 ;
        RECT 452.400 159.600 453.200 160.400 ;
        RECT 434.900 153.700 437.100 154.300 ;
        RECT 434.800 146.200 435.600 151.800 ;
        RECT 436.500 148.400 437.100 153.700 ;
        RECT 436.400 147.600 437.200 148.400 ;
        RECT 438.000 144.200 438.800 155.800 ;
        RECT 446.000 151.600 446.800 152.400 ;
        RECT 444.400 149.600 445.200 150.400 ;
        RECT 442.800 139.600 443.600 140.400 ;
        RECT 441.200 137.600 442.000 138.400 ;
        RECT 436.400 135.600 437.200 136.400 ;
        RECT 434.800 131.600 435.600 132.400 ;
        RECT 414.100 109.700 416.300 110.300 ;
        RECT 406.000 107.600 406.800 108.400 ;
        RECT 412.400 107.600 413.200 108.400 ;
        RECT 404.400 105.600 405.200 106.400 ;
        RECT 402.800 103.600 403.600 104.400 ;
        RECT 407.600 103.600 408.400 104.400 ;
        RECT 402.900 94.400 403.500 103.600 ;
        RECT 407.700 94.400 408.300 103.600 ;
        RECT 412.500 100.300 413.100 107.600 ;
        RECT 410.900 99.700 413.100 100.300 ;
        RECT 409.200 97.600 410.000 98.400 ;
        RECT 410.900 96.400 411.500 99.700 ;
        RECT 410.800 95.600 411.600 96.400 ;
        RECT 399.600 93.700 401.900 94.300 ;
        RECT 399.600 93.600 400.400 93.700 ;
        RECT 402.800 93.600 403.600 94.400 ;
        RECT 404.400 93.600 405.200 94.400 ;
        RECT 407.600 93.600 408.400 94.400 ;
        RECT 396.500 90.400 397.100 93.600 ;
        RECT 396.400 89.600 397.200 90.400 ;
        RECT 402.800 89.600 403.600 90.400 ;
        RECT 404.400 89.600 405.200 90.400 ;
        RECT 407.600 89.600 408.400 90.400 ;
        RECT 402.900 86.400 403.500 89.600 ;
        RECT 402.800 85.600 403.600 86.400 ;
        RECT 396.400 83.600 397.200 84.400 ;
        RECT 401.200 83.600 402.000 84.400 ;
        RECT 396.500 72.400 397.100 83.600 ;
        RECT 391.600 71.600 392.400 72.400 ;
        RECT 394.800 71.600 395.600 72.400 ;
        RECT 396.400 71.600 397.200 72.400 ;
        RECT 401.300 70.400 401.900 83.600 ;
        RECT 380.400 69.600 381.200 70.400 ;
        RECT 385.200 69.600 386.000 70.400 ;
        RECT 388.400 69.600 389.200 70.400 ;
        RECT 401.200 69.600 402.000 70.400 ;
        RECT 380.500 68.400 381.100 69.600 ;
        RECT 372.400 67.600 373.200 68.400 ;
        RECT 378.800 67.600 379.600 68.400 ;
        RECT 380.400 67.600 381.200 68.400 ;
        RECT 386.800 67.600 387.600 68.400 ;
        RECT 393.200 67.600 394.000 68.400 ;
        RECT 399.600 67.600 400.400 68.400 ;
        RECT 404.500 66.400 405.100 89.600 ;
        RECT 410.900 78.400 411.500 95.600 ;
        RECT 412.400 91.600 413.200 92.400 ;
        RECT 412.500 90.400 413.100 91.600 ;
        RECT 412.400 89.600 413.200 90.400 ;
        RECT 410.800 77.600 411.600 78.400 ;
        RECT 394.800 65.600 395.600 66.400 ;
        RECT 398.000 65.600 398.800 66.400 ;
        RECT 404.400 65.600 405.200 66.400 ;
        RECT 406.000 65.600 406.800 66.400 ;
        RECT 394.900 64.400 395.500 65.600 ;
        RECT 380.400 63.600 381.200 64.400 ;
        RECT 391.600 63.600 392.400 64.400 ;
        RECT 394.800 63.600 395.600 64.400 ;
        RECT 380.500 62.400 381.100 63.600 ;
        RECT 377.200 61.600 378.000 62.400 ;
        RECT 380.400 61.600 381.200 62.400 ;
        RECT 372.400 55.600 373.200 56.400 ;
        RECT 372.500 54.400 373.100 55.600 ;
        RECT 372.400 53.600 373.200 54.400 ;
        RECT 377.300 52.400 377.900 61.600 ;
        RECT 391.700 60.400 392.300 63.600 ;
        RECT 391.600 59.600 392.400 60.400 ;
        RECT 343.600 51.600 344.400 52.400 ;
        RECT 354.800 51.600 355.600 52.400 ;
        RECT 358.000 51.600 358.800 52.400 ;
        RECT 359.600 51.600 360.400 52.400 ;
        RECT 364.400 51.600 365.200 52.400 ;
        RECT 369.200 51.600 370.000 52.400 ;
        RECT 377.200 51.600 378.000 52.400 ;
        RECT 324.200 29.600 325.200 30.400 ;
        RECT 334.000 24.200 334.800 37.800 ;
        RECT 335.600 24.200 336.400 37.800 ;
        RECT 337.200 24.200 338.000 37.800 ;
        RECT 338.800 24.200 339.600 35.800 ;
        RECT 340.400 25.600 341.200 26.400 ;
        RECT 335.600 21.600 336.400 22.400 ;
        RECT 335.700 18.400 336.300 21.600 ;
        RECT 340.500 20.400 341.100 25.600 ;
        RECT 342.000 24.200 342.800 35.800 ;
        RECT 343.700 30.400 344.300 51.600 ;
        RECT 369.300 50.400 369.900 51.600 ;
        RECT 369.200 49.600 370.000 50.400 ;
        RECT 343.600 29.600 344.400 30.400 ;
        RECT 343.600 27.600 344.400 28.400 ;
        RECT 343.700 22.400 344.300 27.600 ;
        RECT 345.200 24.200 346.000 35.800 ;
        RECT 346.800 24.200 347.600 37.800 ;
        RECT 348.400 24.200 349.200 37.800 ;
        RECT 377.300 30.400 377.900 51.600 ;
        RECT 382.000 44.200 382.800 57.800 ;
        RECT 383.600 44.200 384.400 57.800 ;
        RECT 385.200 46.200 386.000 57.800 ;
        RECT 386.800 53.600 387.600 54.400 ;
        RECT 388.400 46.200 389.200 57.800 ;
        RECT 390.000 55.600 390.800 56.400 ;
        RECT 390.100 44.300 390.700 55.600 ;
        RECT 391.600 46.200 392.400 57.800 ;
        RECT 388.500 43.700 390.700 44.300 ;
        RECT 393.200 44.200 394.000 57.800 ;
        RECT 394.800 44.200 395.600 57.800 ;
        RECT 396.400 44.200 397.200 57.800 ;
        RECT 377.200 29.600 378.000 30.400 ;
        RECT 359.600 23.600 360.400 24.400 ;
        RECT 343.600 21.600 344.400 22.400 ;
        RECT 359.700 20.400 360.300 23.600 ;
        RECT 377.300 22.400 377.900 29.600 ;
        RECT 380.400 24.200 381.200 37.800 ;
        RECT 382.000 24.200 382.800 37.800 ;
        RECT 383.600 24.200 384.400 35.800 ;
        RECT 385.200 27.600 386.000 28.400 ;
        RECT 386.800 24.200 387.600 35.800 ;
        RECT 388.500 26.400 389.100 43.700 ;
        RECT 388.400 25.600 389.200 26.400 ;
        RECT 367.600 21.600 368.400 22.400 ;
        RECT 377.200 21.600 378.000 22.400 ;
        RECT 340.400 19.600 341.200 20.400 ;
        RECT 354.800 19.600 355.600 20.400 ;
        RECT 359.600 19.600 360.400 20.400 ;
        RECT 335.600 17.600 336.400 18.400 ;
        RECT 324.400 13.600 325.200 14.400 ;
        RECT 330.800 13.600 331.600 14.400 ;
        RECT 329.200 11.600 330.000 12.400 ;
        RECT 332.400 11.600 333.200 12.400 ;
        RECT 332.500 10.400 333.100 11.600 ;
        RECT 321.200 9.600 322.000 10.400 ;
        RECT 332.400 9.600 333.200 10.400 ;
        RECT 338.800 9.600 339.600 10.400 ;
        RECT 348.400 4.200 349.200 17.800 ;
        RECT 350.000 4.200 350.800 17.800 ;
        RECT 351.600 4.200 352.400 17.800 ;
        RECT 353.200 6.200 354.000 17.800 ;
        RECT 354.900 16.400 355.500 19.600 ;
        RECT 354.800 15.600 355.600 16.400 ;
        RECT 356.400 6.200 357.200 17.800 ;
        RECT 358.000 13.600 358.800 14.400 ;
        RECT 358.100 12.400 358.700 13.600 ;
        RECT 358.000 11.600 358.800 12.400 ;
        RECT 359.600 6.200 360.400 17.800 ;
        RECT 361.200 4.200 362.000 17.800 ;
        RECT 362.800 4.200 363.600 17.800 ;
        RECT 367.700 12.400 368.300 21.600 ;
        RECT 386.800 20.300 387.600 20.400 ;
        RECT 388.500 20.300 389.100 25.600 ;
        RECT 390.000 24.200 390.800 35.800 ;
        RECT 391.600 24.200 392.400 37.800 ;
        RECT 393.200 24.200 394.000 37.800 ;
        RECT 394.800 24.200 395.600 37.800 ;
        RECT 396.400 29.600 397.200 30.400 ;
        RECT 390.000 21.600 390.800 22.400 ;
        RECT 386.800 19.700 389.100 20.300 ;
        RECT 386.800 19.600 387.600 19.700 ;
        RECT 367.600 11.600 368.400 12.400 ;
        RECT 382.000 6.200 382.800 17.800 ;
        RECT 386.900 16.400 387.500 19.600 ;
        RECT 386.800 15.600 387.600 16.400 ;
        RECT 386.900 14.400 387.500 15.600 ;
        RECT 386.800 13.600 387.600 14.400 ;
        RECT 390.100 12.600 390.700 21.600 ;
        RECT 390.000 11.800 390.800 12.600 ;
        RECT 390.100 11.700 390.700 11.800 ;
        RECT 391.600 6.200 392.400 17.800 ;
        RECT 394.800 10.200 395.600 15.800 ;
        RECT 396.500 12.400 397.100 29.600 ;
        RECT 398.100 22.400 398.700 65.600 ;
        RECT 402.800 63.600 403.600 64.400 ;
        RECT 404.400 63.600 405.200 64.400 ;
        RECT 402.900 28.400 403.500 63.600 ;
        RECT 404.500 38.400 405.100 63.600 ;
        RECT 406.100 58.400 406.700 65.600 ;
        RECT 406.000 57.600 406.800 58.400 ;
        RECT 409.200 53.600 410.000 54.400 ;
        RECT 410.800 53.600 411.600 54.400 ;
        RECT 404.400 37.600 405.200 38.400 ;
        RECT 407.600 33.600 408.400 34.400 ;
        RECT 402.800 27.600 403.600 28.400 ;
        RECT 407.700 26.400 408.300 33.600 ;
        RECT 407.600 25.600 408.400 26.400 ;
        RECT 398.000 21.600 398.800 22.400 ;
        RECT 396.400 11.600 397.200 12.400 ;
        RECT 399.600 11.600 400.400 12.400 ;
        RECT 404.400 4.200 405.200 17.800 ;
        RECT 406.000 4.200 406.800 17.800 ;
        RECT 407.600 6.200 408.400 17.800 ;
        RECT 409.300 14.400 409.900 53.600 ;
        RECT 410.900 52.400 411.500 53.600 ;
        RECT 412.500 52.400 413.100 89.600 ;
        RECT 410.800 51.600 411.600 52.400 ;
        RECT 412.400 51.600 413.200 52.400 ;
        RECT 414.100 38.400 414.700 109.700 ;
        RECT 417.200 109.600 418.000 110.400 ;
        RECT 418.800 109.600 419.600 110.400 ;
        RECT 431.600 109.600 432.400 110.400 ;
        RECT 433.200 109.600 434.000 110.400 ;
        RECT 418.800 108.300 419.600 108.400 ;
        RECT 417.300 107.700 419.600 108.300 ;
        RECT 417.300 98.400 417.900 107.700 ;
        RECT 418.800 107.600 419.600 107.700 ;
        RECT 423.600 107.600 424.400 108.400 ;
        RECT 431.600 107.600 432.400 108.400 ;
        RECT 433.200 107.600 434.000 108.400 ;
        RECT 423.700 106.400 424.300 107.600 ;
        RECT 423.600 105.600 424.400 106.400 ;
        RECT 431.700 104.400 432.300 107.600 ;
        RECT 433.300 106.400 433.900 107.600 ;
        RECT 433.200 105.600 434.000 106.400 ;
        RECT 422.000 103.600 422.800 104.400 ;
        RECT 431.600 103.600 432.400 104.400 ;
        RECT 422.100 102.400 422.700 103.600 ;
        RECT 422.000 101.600 422.800 102.400 ;
        RECT 431.700 98.400 432.300 103.600 ;
        RECT 415.600 97.600 416.400 98.400 ;
        RECT 417.200 97.600 418.000 98.400 ;
        RECT 431.600 97.600 432.400 98.400 ;
        RECT 415.700 96.400 416.300 97.600 ;
        RECT 415.600 95.600 416.400 96.400 ;
        RECT 430.000 95.600 430.800 96.400 ;
        RECT 433.200 96.300 434.000 96.400 ;
        RECT 434.900 96.300 435.500 131.600 ;
        RECT 436.500 130.400 437.100 135.600 ;
        RECT 441.300 132.400 441.900 137.600 ;
        RECT 442.900 134.400 443.500 139.600 ;
        RECT 442.800 133.600 443.600 134.400 ;
        RECT 439.600 132.300 440.400 132.400 ;
        RECT 438.100 131.700 440.400 132.300 ;
        RECT 436.400 129.600 437.200 130.400 ;
        RECT 438.100 110.400 438.700 131.700 ;
        RECT 439.600 131.600 440.400 131.700 ;
        RECT 441.200 131.600 442.000 132.400 ;
        RECT 444.500 118.400 445.100 149.600 ;
        RECT 446.100 136.400 446.700 151.600 ;
        RECT 447.600 144.200 448.400 155.800 ;
        RECT 452.500 150.400 453.100 159.600 ;
        RECT 454.100 152.400 454.700 163.600 ;
        RECT 455.700 154.400 456.300 171.600 ;
        RECT 462.000 159.600 462.800 160.400 ;
        RECT 462.100 158.400 462.700 159.600 ;
        RECT 463.700 158.400 464.300 173.600 ;
        RECT 468.500 168.400 469.100 175.600 ;
        RECT 470.100 172.400 470.700 175.600 ;
        RECT 470.000 171.600 470.800 172.400 ;
        RECT 484.400 171.600 485.200 172.400 ;
        RECT 484.500 168.400 485.100 171.600 ;
        RECT 486.100 168.400 486.700 175.600 ;
        RECT 498.900 174.400 499.500 187.600 ;
        RECT 500.400 185.600 501.200 186.400 ;
        RECT 498.800 173.600 499.600 174.400 ;
        RECT 468.400 167.600 469.200 168.400 ;
        RECT 474.800 167.600 475.600 168.400 ;
        RECT 479.600 167.600 480.400 168.400 ;
        RECT 484.400 167.600 485.200 168.400 ;
        RECT 486.000 167.600 486.800 168.400 ;
        RECT 489.200 167.600 490.000 168.400 ;
        RECT 494.000 167.600 494.800 168.400 ;
        RECT 468.500 166.400 469.100 167.600 ;
        RECT 474.900 166.400 475.500 167.600 ;
        RECT 466.800 165.600 467.600 166.400 ;
        RECT 468.400 165.600 469.200 166.400 ;
        RECT 474.800 165.600 475.600 166.400 ;
        RECT 462.000 157.600 462.800 158.400 ;
        RECT 463.600 157.600 464.400 158.400 ;
        RECT 458.800 155.600 459.600 156.400 ;
        RECT 455.600 153.600 456.400 154.400 ;
        RECT 457.200 153.600 458.000 154.400 ;
        RECT 454.000 151.600 454.800 152.400 ;
        RECT 457.300 150.400 457.900 153.600 ;
        RECT 452.400 149.600 453.200 150.400 ;
        RECT 455.600 149.600 456.400 150.400 ;
        RECT 457.200 149.600 458.000 150.400 ;
        RECT 452.400 147.600 453.200 148.400 ;
        RECT 454.000 145.600 454.800 146.400 ;
        RECT 450.800 143.600 451.600 144.400 ;
        RECT 450.900 138.400 451.500 143.600 ;
        RECT 454.000 141.600 454.800 142.400 ;
        RECT 450.800 137.600 451.600 138.400 ;
        RECT 446.000 135.600 446.800 136.400 ;
        RECT 454.100 134.400 454.700 141.600 ;
        RECT 454.000 133.600 454.800 134.400 ;
        RECT 455.700 132.400 456.300 149.600 ;
        RECT 458.900 132.400 459.500 155.600 ;
        RECT 463.600 153.600 464.400 154.400 ;
        RECT 479.700 152.400 480.300 167.600 ;
        RECT 497.200 165.600 498.000 166.400 ;
        RECT 487.600 163.600 488.400 164.400 ;
        RECT 495.600 163.600 496.400 164.400 ;
        RECT 481.200 157.600 482.000 158.400 ;
        RECT 471.600 151.600 472.400 152.400 ;
        RECT 479.600 151.600 480.400 152.400 ;
        RECT 471.700 150.400 472.300 151.600 ;
        RECT 481.300 150.400 481.900 157.600 ;
        RECT 487.700 156.400 488.300 163.600 ;
        RECT 495.700 160.400 496.300 163.600 ;
        RECT 495.600 159.600 496.400 160.400 ;
        RECT 487.600 155.600 488.400 156.400 ;
        RECT 487.700 154.400 488.300 155.600 ;
        RECT 487.600 153.600 488.400 154.400 ;
        RECT 494.000 153.600 494.800 154.400 ;
        RECT 494.100 150.400 494.700 153.600 ;
        RECT 471.600 149.600 472.400 150.400 ;
        RECT 481.200 149.600 482.000 150.400 ;
        RECT 486.000 149.600 486.800 150.400 ;
        RECT 487.600 149.600 488.400 150.400 ;
        RECT 494.000 149.600 494.800 150.400 ;
        RECT 495.700 150.300 496.300 159.600 ;
        RECT 497.300 158.400 497.900 165.600 ;
        RECT 497.200 157.600 498.000 158.400 ;
        RECT 498.800 153.600 499.600 154.400 ;
        RECT 497.200 150.300 498.000 150.400 ;
        RECT 495.700 149.700 498.000 150.300 ;
        RECT 486.100 146.400 486.700 149.600 ;
        RECT 492.400 147.600 493.200 148.400 ;
        RECT 486.000 145.600 486.800 146.400 ;
        RECT 489.200 145.600 490.000 146.400 ;
        RECT 490.800 145.600 491.600 146.400 ;
        RECT 470.000 143.600 470.800 144.400 ;
        RECT 482.800 143.600 483.600 144.400 ;
        RECT 463.600 141.600 464.400 142.400 ;
        RECT 463.700 136.400 464.300 141.600 ;
        RECT 463.600 135.600 464.400 136.400 ;
        RECT 470.100 134.400 470.700 143.600 ;
        RECT 482.900 142.400 483.500 143.600 ;
        RECT 478.000 141.600 478.800 142.400 ;
        RECT 482.800 141.600 483.600 142.400 ;
        RECT 470.000 133.600 470.800 134.400 ;
        RECT 449.200 131.600 450.000 132.400 ;
        RECT 455.600 131.600 456.400 132.400 ;
        RECT 458.800 131.600 459.600 132.400 ;
        RECT 470.000 131.600 470.800 132.400 ;
        RECT 449.300 130.400 449.900 131.600 ;
        RECT 447.600 129.600 448.400 130.400 ;
        RECT 449.200 129.600 450.000 130.400 ;
        RECT 447.700 128.400 448.300 129.600 ;
        RECT 470.100 128.400 470.700 131.600 ;
        RECT 447.600 127.600 448.400 128.400 ;
        RECT 454.000 127.600 454.800 128.400 ;
        RECT 470.000 127.600 470.800 128.400 ;
        RECT 454.100 126.400 454.700 127.600 ;
        RECT 454.000 125.600 454.800 126.400 ;
        RECT 442.800 117.600 443.600 118.400 ;
        RECT 444.400 117.600 445.200 118.400 ;
        RECT 442.900 114.400 443.500 117.600 ;
        RECT 442.800 113.600 443.600 114.400 ;
        RECT 439.600 111.600 440.400 112.400 ;
        RECT 452.400 111.600 453.200 112.400 ;
        RECT 438.000 109.600 438.800 110.400 ;
        RECT 441.200 109.600 442.000 110.400 ;
        RECT 446.000 109.600 446.800 110.400 ;
        RECT 447.600 109.600 448.400 110.400 ;
        RECT 438.000 107.600 438.800 108.400 ;
        RECT 438.100 96.400 438.700 107.600 ;
        RECT 441.300 102.400 441.900 109.600 ;
        RECT 446.100 104.400 446.700 109.600 ;
        RECT 447.700 108.400 448.300 109.600 ;
        RECT 447.600 107.600 448.400 108.400 ;
        RECT 449.200 107.600 450.000 108.400 ;
        RECT 446.000 103.600 446.800 104.400 ;
        RECT 441.200 101.600 442.000 102.400 ;
        RECT 446.000 99.600 446.800 100.400 ;
        RECT 433.200 95.700 435.500 96.300 ;
        RECT 433.200 95.600 434.000 95.700 ;
        RECT 438.000 95.600 438.800 96.400 ;
        RECT 415.700 92.400 416.300 95.600 ;
        RECT 415.600 91.600 416.400 92.400 ;
        RECT 430.100 86.400 430.700 95.600 ;
        RECT 446.100 94.400 446.700 99.600 ;
        RECT 452.500 96.400 453.100 111.600 ;
        RECT 454.100 98.400 454.700 125.600 ;
        RECT 457.200 123.600 458.000 124.400 ;
        RECT 462.000 123.600 462.800 124.400 ;
        RECT 473.200 124.200 474.000 137.800 ;
        RECT 474.800 124.200 475.600 137.800 ;
        RECT 476.400 126.200 477.200 137.800 ;
        RECT 478.100 134.400 478.700 141.600 ;
        RECT 489.200 139.600 490.000 140.400 ;
        RECT 478.000 133.600 478.800 134.400 ;
        RECT 479.600 126.200 480.400 137.800 ;
        RECT 481.200 135.600 482.000 136.400 ;
        RECT 481.200 129.600 482.000 130.400 ;
        RECT 455.600 119.600 456.400 120.400 ;
        RECT 455.700 110.400 456.300 119.600 ;
        RECT 457.300 110.400 457.900 123.600 ;
        RECT 460.400 113.600 461.200 114.400 ;
        RECT 455.600 109.600 456.400 110.400 ;
        RECT 457.200 109.600 458.000 110.400 ;
        RECT 458.800 109.600 459.600 110.400 ;
        RECT 458.900 108.400 459.500 109.600 ;
        RECT 455.600 107.600 456.400 108.400 ;
        RECT 457.200 107.600 458.000 108.400 ;
        RECT 458.800 107.600 459.600 108.400 ;
        RECT 454.000 97.600 454.800 98.400 ;
        RECT 455.600 97.600 456.400 98.400 ;
        RECT 452.400 95.600 453.200 96.400 ;
        RECT 436.400 93.600 437.200 94.400 ;
        RECT 438.000 93.600 438.800 94.400 ;
        RECT 441.200 93.600 442.000 94.400 ;
        RECT 446.000 93.600 446.800 94.400 ;
        RECT 436.500 86.400 437.100 93.600 ;
        RECT 438.100 92.400 438.700 93.600 ;
        RECT 441.300 92.400 441.900 93.600 ;
        RECT 455.700 92.400 456.300 97.600 ;
        RECT 438.000 91.600 438.800 92.400 ;
        RECT 441.200 91.600 442.000 92.400 ;
        RECT 455.600 91.600 456.400 92.400 ;
        RECT 439.600 89.600 440.400 90.400 ;
        RECT 449.200 89.600 450.000 90.400 ;
        RECT 455.600 89.600 456.400 90.400 ;
        RECT 439.700 88.400 440.300 89.600 ;
        RECT 439.600 87.600 440.400 88.400 ;
        RECT 441.200 87.600 442.000 88.400 ;
        RECT 417.200 85.600 418.000 86.400 ;
        RECT 430.000 85.600 430.800 86.400 ;
        RECT 436.400 85.600 437.200 86.400 ;
        RECT 417.300 78.400 417.900 85.600 ;
        RECT 441.300 84.400 441.900 87.600 ;
        RECT 442.800 85.600 443.600 86.400 ;
        RECT 418.800 83.600 419.600 84.400 ;
        RECT 433.200 83.600 434.000 84.400 ;
        RECT 441.200 83.600 442.000 84.400 ;
        RECT 436.400 81.600 437.200 82.400 ;
        RECT 417.200 77.600 418.000 78.400 ;
        RECT 425.200 71.600 426.000 72.400 ;
        RECT 418.800 55.600 419.600 56.400 ;
        RECT 420.400 55.600 421.200 56.400 ;
        RECT 418.900 52.400 419.500 55.600 ;
        RECT 425.300 54.400 425.900 71.600 ;
        RECT 426.800 64.200 427.600 77.800 ;
        RECT 428.400 64.200 429.200 77.800 ;
        RECT 430.000 64.200 430.800 77.800 ;
        RECT 431.600 64.200 432.400 75.800 ;
        RECT 433.200 65.600 434.000 66.400 ;
        RECT 425.200 53.600 426.000 54.400 ;
        RECT 430.000 53.600 430.800 54.400 ;
        RECT 425.300 52.400 425.900 53.600 ;
        RECT 415.600 51.600 416.400 52.400 ;
        RECT 417.200 51.600 418.000 52.400 ;
        RECT 418.800 51.600 419.600 52.400 ;
        RECT 425.200 51.600 426.000 52.400 ;
        RECT 415.700 48.400 416.300 51.600 ;
        RECT 415.600 47.600 416.400 48.400 ;
        RECT 418.800 47.600 419.600 48.400 ;
        RECT 430.000 47.600 430.800 48.400 ;
        RECT 414.000 37.600 414.800 38.400 ;
        RECT 420.400 29.600 421.200 30.400 ;
        RECT 409.200 13.600 410.000 14.400 ;
        RECT 410.800 6.200 411.600 17.800 ;
        RECT 412.400 15.600 413.200 16.400 ;
        RECT 414.000 6.200 414.800 17.800 ;
        RECT 415.600 4.200 416.400 17.800 ;
        RECT 417.200 4.200 418.000 17.800 ;
        RECT 418.800 4.200 419.600 17.800 ;
        RECT 420.500 12.400 421.100 29.600 ;
        RECT 425.200 24.200 426.000 37.800 ;
        RECT 426.800 24.200 427.600 37.800 ;
        RECT 428.400 24.200 429.200 35.800 ;
        RECT 430.100 28.400 430.700 47.600 ;
        RECT 430.000 27.600 430.800 28.400 ;
        RECT 431.600 24.200 432.400 35.800 ;
        RECT 433.300 26.400 433.900 65.600 ;
        RECT 434.800 64.200 435.600 75.800 ;
        RECT 436.500 68.400 437.100 81.600 ;
        RECT 436.400 67.600 437.200 68.400 ;
        RECT 438.000 64.200 438.800 75.800 ;
        RECT 439.600 64.200 440.400 77.800 ;
        RECT 441.200 64.200 442.000 77.800 ;
        RECT 442.900 58.400 443.500 85.600 ;
        RECT 444.400 83.600 445.200 84.400 ;
        RECT 447.600 83.600 448.400 84.400 ;
        RECT 454.000 83.600 454.800 84.400 ;
        RECT 447.700 74.400 448.300 83.600 ;
        RECT 447.600 73.600 448.400 74.400 ;
        RECT 450.800 73.600 451.600 74.400 ;
        RECT 450.900 72.400 451.500 73.600 ;
        RECT 450.800 71.600 451.600 72.400 ;
        RECT 454.100 70.400 454.700 83.600 ;
        RECT 455.700 70.400 456.300 89.600 ;
        RECT 457.300 78.400 457.900 107.600 ;
        RECT 458.800 97.600 459.600 98.400 ;
        RECT 458.900 94.400 459.500 97.600 ;
        RECT 458.800 93.600 459.600 94.400 ;
        RECT 460.500 92.300 461.100 113.600 ;
        RECT 462.100 112.400 462.700 123.600 ;
        RECT 481.300 118.400 481.900 129.600 ;
        RECT 482.800 126.200 483.600 137.800 ;
        RECT 484.400 124.200 485.200 137.800 ;
        RECT 486.000 124.200 486.800 137.800 ;
        RECT 487.600 124.200 488.400 137.800 ;
        RECT 481.200 117.600 482.000 118.400 ;
        RECT 484.400 113.600 485.200 114.400 ;
        RECT 487.600 113.600 488.400 114.400 ;
        RECT 462.000 111.600 462.800 112.400 ;
        RECT 471.600 111.600 472.400 112.400 ;
        RECT 473.200 111.600 474.000 112.400 ;
        RECT 462.000 109.600 462.800 110.400 ;
        RECT 463.600 109.600 464.400 110.400 ;
        RECT 466.800 109.600 467.600 110.400 ;
        RECT 471.600 109.600 472.400 110.400 ;
        RECT 462.100 106.300 462.700 109.600 ;
        RECT 471.700 106.400 472.300 109.600 ;
        RECT 473.300 108.400 473.900 111.600 ;
        RECT 484.500 110.400 485.100 113.600 ;
        RECT 476.400 109.600 477.200 110.400 ;
        RECT 479.600 109.600 480.400 110.400 ;
        RECT 482.800 109.600 483.600 110.400 ;
        RECT 484.400 109.600 485.200 110.400 ;
        RECT 486.000 109.600 486.800 110.400 ;
        RECT 473.200 107.600 474.000 108.400 ;
        RECT 478.000 107.600 478.800 108.400 ;
        RECT 463.600 106.300 464.400 106.400 ;
        RECT 462.100 105.700 464.400 106.300 ;
        RECT 463.600 105.600 464.400 105.700 ;
        RECT 471.600 105.600 472.400 106.400 ;
        RECT 465.200 103.600 466.000 104.400 ;
        RECT 470.000 103.600 470.800 104.400 ;
        RECT 465.300 96.400 465.900 103.600 ;
        RECT 468.400 101.600 469.200 102.400 ;
        RECT 468.500 98.400 469.100 101.600 ;
        RECT 468.400 97.600 469.200 98.400 ;
        RECT 465.200 95.600 466.000 96.400 ;
        RECT 468.400 95.600 469.200 96.400 ;
        RECT 465.200 93.600 466.000 94.400 ;
        RECT 466.800 93.600 467.600 94.400 ;
        RECT 465.300 92.400 465.900 93.600 ;
        RECT 462.000 92.300 462.800 92.400 ;
        RECT 460.500 91.700 462.800 92.300 ;
        RECT 462.000 91.600 462.800 91.700 ;
        RECT 463.600 91.600 464.400 92.400 ;
        RECT 465.200 91.600 466.000 92.400 ;
        RECT 460.400 83.600 461.200 84.400 ;
        RECT 457.200 77.600 458.000 78.400 ;
        RECT 460.500 70.400 461.100 83.600 ;
        RECT 446.000 69.600 446.800 70.400 ;
        RECT 454.000 69.600 454.800 70.400 ;
        RECT 455.600 69.600 456.400 70.400 ;
        RECT 460.400 69.600 461.200 70.400 ;
        RECT 449.200 65.600 450.000 66.400 ;
        RECT 447.600 63.600 448.400 64.400 ;
        RECT 442.800 57.600 443.600 58.400 ;
        RECT 438.000 54.300 438.800 54.400 ;
        RECT 434.900 53.700 438.800 54.300 ;
        RECT 434.900 52.400 435.500 53.700 ;
        RECT 438.000 53.600 438.800 53.700 ;
        RECT 434.800 51.600 435.600 52.400 ;
        RECT 436.400 51.600 437.200 52.400 ;
        RECT 442.800 51.600 443.600 52.400 ;
        RECT 436.500 50.400 437.100 51.600 ;
        RECT 436.400 49.600 437.200 50.400 ;
        RECT 433.200 25.600 434.000 26.400 ;
        RECT 428.400 21.600 429.200 22.400 ;
        RECT 428.500 18.400 429.100 21.600 ;
        RECT 428.400 17.600 429.200 18.400 ;
        RECT 433.300 16.400 433.900 25.600 ;
        RECT 434.800 24.200 435.600 35.800 ;
        RECT 436.400 24.200 437.200 37.800 ;
        RECT 438.000 24.200 438.800 37.800 ;
        RECT 439.600 24.200 440.400 37.800 ;
        RECT 433.200 15.600 434.000 16.400 ;
        RECT 420.400 11.600 421.200 12.400 ;
        RECT 438.000 10.200 438.800 15.800 ;
        RECT 441.200 6.200 442.000 17.800 ;
        RECT 442.900 12.600 443.500 51.600 ;
        RECT 447.700 48.400 448.300 63.600 ;
        RECT 449.300 52.400 449.900 65.600 ;
        RECT 450.800 63.600 451.600 64.400 ;
        RECT 454.100 62.400 454.700 69.600 ;
        RECT 455.700 64.400 456.300 69.600 ;
        RECT 465.300 68.400 465.900 91.600 ;
        RECT 466.900 78.400 467.500 93.600 ;
        RECT 466.800 77.600 467.600 78.400 ;
        RECT 466.800 72.300 467.600 72.400 ;
        RECT 468.500 72.300 469.100 95.600 ;
        RECT 470.100 72.400 470.700 103.600 ;
        RECT 471.700 94.400 472.300 105.600 ;
        RECT 478.100 98.400 478.700 107.600 ;
        RECT 474.800 97.600 475.600 98.400 ;
        RECT 478.000 97.600 478.800 98.400 ;
        RECT 479.700 94.400 480.300 109.600 ;
        RECT 486.100 108.400 486.700 109.600 ;
        RECT 481.200 107.600 482.000 108.400 ;
        RECT 482.800 107.600 483.600 108.400 ;
        RECT 486.000 107.600 486.800 108.400 ;
        RECT 481.300 106.400 481.900 107.600 ;
        RECT 481.200 105.600 482.000 106.400 ;
        RECT 482.900 98.400 483.500 107.600 ;
        RECT 482.800 97.600 483.600 98.400 ;
        RECT 471.600 93.600 472.400 94.400 ;
        RECT 479.600 93.600 480.400 94.400 ;
        RECT 479.700 92.400 480.300 93.600 ;
        RECT 487.700 92.400 488.300 113.600 ;
        RECT 489.300 106.400 489.900 139.600 ;
        RECT 490.900 110.400 491.500 145.600 ;
        RECT 492.500 116.400 493.100 147.600 ;
        RECT 492.400 115.600 493.200 116.400 ;
        RECT 495.700 112.400 496.300 149.700 ;
        RECT 497.200 149.600 498.000 149.700 ;
        RECT 498.900 148.400 499.500 153.600 ;
        RECT 500.500 152.300 501.100 185.600 ;
        RECT 502.000 175.600 502.800 176.400 ;
        RECT 502.000 173.600 502.800 174.400 ;
        RECT 503.700 166.400 504.300 187.600 ;
        RECT 508.500 182.400 509.100 189.600 ;
        RECT 510.000 187.600 510.800 188.400 ;
        RECT 508.400 181.600 509.200 182.400 ;
        RECT 505.200 173.600 506.000 174.400 ;
        RECT 506.800 173.600 507.600 174.400 ;
        RECT 508.400 173.600 509.200 174.400 ;
        RECT 506.900 172.400 507.500 173.600 ;
        RECT 505.200 171.600 506.000 172.400 ;
        RECT 506.800 171.600 507.600 172.400 ;
        RECT 503.600 165.600 504.400 166.400 ;
        RECT 502.000 163.600 502.800 164.400 ;
        RECT 500.500 151.700 502.700 152.300 ;
        RECT 502.100 150.400 502.700 151.700 ;
        RECT 500.400 149.600 501.200 150.400 ;
        RECT 502.000 149.600 502.800 150.400 ;
        RECT 498.800 147.600 499.600 148.400 ;
        RECT 497.200 145.600 498.000 146.400 ;
        RECT 497.300 138.400 497.900 145.600 ;
        RECT 497.200 137.600 498.000 138.400 ;
        RECT 500.500 132.400 501.100 149.600 ;
        RECT 503.600 143.600 504.400 144.400 ;
        RECT 503.700 142.400 504.300 143.600 ;
        RECT 503.600 141.600 504.400 142.400 ;
        RECT 500.400 131.600 501.200 132.400 ;
        RECT 502.000 131.600 502.800 132.400 ;
        RECT 497.200 129.600 498.000 130.400 ;
        RECT 497.300 112.400 497.900 129.600 ;
        RECT 500.500 114.400 501.100 131.600 ;
        RECT 500.400 113.600 501.200 114.400 ;
        RECT 495.600 111.600 496.400 112.400 ;
        RECT 497.200 111.600 498.000 112.400 ;
        RECT 490.800 109.600 491.600 110.400 ;
        RECT 500.400 109.600 501.200 110.400 ;
        RECT 490.800 107.600 491.600 108.400 ;
        RECT 492.400 107.600 493.200 108.400 ;
        RECT 498.800 107.600 499.600 108.400 ;
        RECT 490.900 106.400 491.500 107.600 ;
        RECT 500.500 106.400 501.100 109.600 ;
        RECT 489.200 105.600 490.000 106.400 ;
        RECT 490.800 105.600 491.600 106.400 ;
        RECT 500.400 105.600 501.200 106.400 ;
        RECT 497.200 103.600 498.000 104.400 ;
        RECT 497.300 100.400 497.900 103.600 ;
        RECT 497.200 99.600 498.000 100.400 ;
        RECT 502.100 98.400 502.700 131.600 ;
        RECT 505.300 126.400 505.900 171.600 ;
        RECT 508.500 164.400 509.100 173.600 ;
        RECT 510.100 172.400 510.700 187.600 ;
        RECT 511.600 181.600 512.400 182.400 ;
        RECT 511.700 178.400 512.300 181.600 ;
        RECT 511.600 177.600 512.400 178.400 ;
        RECT 513.300 174.400 513.900 189.600 ;
        RECT 514.800 187.600 515.600 188.400 ;
        RECT 514.900 178.400 515.500 187.600 ;
        RECT 514.800 177.600 515.600 178.400 ;
        RECT 513.200 173.600 514.000 174.400 ;
        RECT 510.000 171.600 510.800 172.400 ;
        RECT 511.600 169.600 512.400 170.400 ;
        RECT 510.000 165.600 510.800 166.400 ;
        RECT 508.400 163.600 509.200 164.400 ;
        RECT 510.100 158.400 510.700 165.600 ;
        RECT 511.700 162.400 512.300 169.600 ;
        RECT 511.600 161.600 512.400 162.400 ;
        RECT 510.000 157.600 510.800 158.400 ;
        RECT 516.500 154.400 517.100 191.600 ;
        RECT 518.000 189.600 518.800 190.400 ;
        RECT 518.100 188.400 518.700 189.600 ;
        RECT 518.000 187.600 518.800 188.400 ;
        RECT 506.800 153.600 507.600 154.400 ;
        RECT 511.600 153.600 512.400 154.400 ;
        RECT 516.400 153.600 517.200 154.400 ;
        RECT 506.900 150.400 507.500 153.600 ;
        RECT 508.400 151.600 509.200 152.400 ;
        RECT 510.000 151.600 510.800 152.400 ;
        RECT 508.500 150.400 509.100 151.600 ;
        RECT 506.800 149.600 507.600 150.400 ;
        RECT 508.400 149.600 509.200 150.400 ;
        RECT 510.100 148.400 510.700 151.600 ;
        RECT 516.400 149.600 517.200 150.400 ;
        RECT 518.000 149.600 518.800 150.400 ;
        RECT 518.100 148.400 518.700 149.600 ;
        RECT 510.000 147.600 510.800 148.400 ;
        RECT 511.600 147.600 512.400 148.400 ;
        RECT 518.000 147.600 518.800 148.400 ;
        RECT 511.700 146.400 512.300 147.600 ;
        RECT 511.600 146.300 512.400 146.400 ;
        RECT 510.100 145.700 512.400 146.300 ;
        RECT 510.100 134.400 510.700 145.700 ;
        RECT 511.600 145.600 512.400 145.700 ;
        RECT 514.800 145.600 515.600 146.400 ;
        RECT 514.900 136.400 515.500 145.600 ;
        RECT 514.800 135.600 515.600 136.400 ;
        RECT 510.000 133.600 510.800 134.400 ;
        RECT 506.800 131.600 507.600 132.400 ;
        RECT 513.200 129.600 514.000 130.400 ;
        RECT 510.000 127.600 510.800 128.400 ;
        RECT 505.200 125.600 506.000 126.400 ;
        RECT 505.200 123.600 506.000 124.400 ;
        RECT 505.300 114.400 505.900 123.600 ;
        RECT 505.200 113.600 506.000 114.400 ;
        RECT 510.100 112.400 510.700 127.600 ;
        RECT 514.800 119.600 515.600 120.400 ;
        RECT 513.200 113.600 514.000 114.400 ;
        RECT 505.200 111.600 506.000 112.400 ;
        RECT 510.000 111.600 510.800 112.400 ;
        RECT 513.300 110.400 513.900 113.600 ;
        RECT 513.200 109.600 514.000 110.400 ;
        RECT 514.900 108.400 515.500 119.600 ;
        RECT 518.100 118.400 518.700 147.600 ;
        RECT 519.700 130.400 520.300 191.600 ;
        RECT 521.200 186.200 522.000 191.800 ;
        RECT 521.200 183.600 522.000 184.400 ;
        RECT 521.300 158.400 521.900 183.600 ;
        RECT 522.900 174.400 523.500 201.600 ;
        RECT 524.400 184.200 525.200 195.800 ;
        RECT 530.900 190.400 531.500 215.600 ;
        RECT 532.400 206.200 533.200 217.800 ;
        RECT 534.000 204.200 534.800 217.800 ;
        RECT 535.600 204.200 536.400 217.800 ;
        RECT 537.200 204.200 538.000 217.800 ;
        RECT 542.000 213.600 542.800 214.400 ;
        RECT 540.400 211.600 541.200 212.400 ;
        RECT 527.600 189.600 528.400 190.400 ;
        RECT 530.800 189.600 531.600 190.400 ;
        RECT 527.700 182.400 528.300 189.600 ;
        RECT 527.600 181.600 528.400 182.400 ;
        RECT 522.800 173.600 523.600 174.400 ;
        RECT 522.800 171.600 523.600 172.400 ;
        RECT 521.200 157.600 522.000 158.400 ;
        RECT 519.600 129.600 520.400 130.400 ;
        RECT 518.000 117.600 518.800 118.400 ;
        RECT 508.400 107.600 509.200 108.400 ;
        RECT 511.600 107.600 512.400 108.400 ;
        RECT 514.800 107.600 515.600 108.400 ;
        RECT 503.600 103.600 504.400 104.400 ;
        RECT 503.700 100.400 504.300 103.600 ;
        RECT 503.600 99.600 504.400 100.400 ;
        RECT 508.500 98.400 509.100 107.600 ;
        RECT 511.700 106.400 512.300 107.600 ;
        RECT 511.600 105.600 512.400 106.400 ;
        RECT 471.600 91.600 472.400 92.400 ;
        RECT 473.200 91.600 474.000 92.400 ;
        RECT 479.600 91.600 480.400 92.400 ;
        RECT 487.600 91.600 488.400 92.400 ;
        RECT 471.700 74.400 472.300 91.600 ;
        RECT 473.300 90.400 473.900 91.600 ;
        RECT 473.200 89.600 474.000 90.400 ;
        RECT 478.000 89.600 478.800 90.400 ;
        RECT 471.600 73.600 472.400 74.400 ;
        RECT 466.800 71.700 469.100 72.300 ;
        RECT 466.800 71.600 467.600 71.700 ;
        RECT 470.000 71.600 470.800 72.400 ;
        RECT 478.100 70.400 478.700 89.600 ;
        RECT 484.400 77.600 485.200 78.400 ;
        RECT 484.500 74.400 485.100 77.600 ;
        RECT 484.400 73.600 485.200 74.400 ;
        RECT 484.500 70.400 485.100 73.600 ;
        RECT 487.700 70.400 488.300 91.600 ;
        RECT 492.400 84.200 493.200 97.800 ;
        RECT 494.000 84.200 494.800 97.800 ;
        RECT 495.600 84.200 496.400 97.800 ;
        RECT 497.200 86.200 498.000 97.800 ;
        RECT 498.800 95.600 499.600 96.400 ;
        RECT 500.400 86.200 501.200 97.800 ;
        RECT 502.000 97.600 502.800 98.400 ;
        RECT 502.000 93.600 502.800 94.400 ;
        RECT 502.100 78.400 502.700 93.600 ;
        RECT 503.600 86.200 504.400 97.800 ;
        RECT 505.200 84.200 506.000 97.800 ;
        RECT 506.800 84.200 507.600 97.800 ;
        RECT 508.400 97.600 509.200 98.400 ;
        RECT 511.600 91.600 512.400 92.400 ;
        RECT 502.000 77.600 502.800 78.400 ;
        RECT 514.900 76.400 515.500 107.600 ;
        RECT 518.000 97.600 518.800 98.400 ;
        RECT 498.800 75.600 499.600 76.400 ;
        RECT 503.600 75.600 504.400 76.400 ;
        RECT 506.800 75.600 507.600 76.400 ;
        RECT 514.800 75.600 515.600 76.400 ;
        RECT 498.900 72.400 499.500 75.600 ;
        RECT 490.800 71.600 491.600 72.400 ;
        RECT 497.200 71.600 498.000 72.400 ;
        RECT 498.800 71.600 499.600 72.400 ;
        RECT 497.300 70.400 497.900 71.600 ;
        RECT 466.800 69.600 467.600 70.400 ;
        RECT 476.400 69.600 477.200 70.400 ;
        RECT 478.000 69.600 478.800 70.400 ;
        RECT 484.400 69.600 485.200 70.400 ;
        RECT 487.600 70.300 488.400 70.400 ;
        RECT 487.600 69.700 489.900 70.300 ;
        RECT 487.600 69.600 488.400 69.700 ;
        RECT 458.800 67.600 459.600 68.400 ;
        RECT 465.200 67.600 466.000 68.400 ;
        RECT 458.800 65.600 459.600 66.400 ;
        RECT 460.400 65.600 461.200 66.400 ;
        RECT 455.600 63.600 456.400 64.400 ;
        RECT 450.800 61.600 451.600 62.400 ;
        RECT 454.000 61.600 454.800 62.400 ;
        RECT 450.900 52.400 451.500 61.600 ;
        RECT 460.500 60.400 461.100 65.600 ;
        RECT 466.900 60.400 467.500 69.600 ;
        RECT 474.800 67.600 475.600 68.400 ;
        RECT 468.400 65.600 469.200 66.400 ;
        RECT 471.600 65.600 472.400 66.400 ;
        RECT 468.500 62.400 469.100 65.600 ;
        RECT 468.400 61.600 469.200 62.400 ;
        RECT 460.400 59.600 461.200 60.400 ;
        RECT 466.800 59.600 467.600 60.400 ;
        RECT 471.700 58.400 472.300 65.600 ;
        RECT 449.200 51.600 450.000 52.400 ;
        RECT 450.800 51.600 451.600 52.400 ;
        RECT 447.600 47.600 448.400 48.400 ;
        RECT 449.300 38.400 449.900 51.600 ;
        RECT 452.400 44.200 453.200 57.800 ;
        RECT 454.000 44.200 454.800 57.800 ;
        RECT 455.600 44.200 456.400 57.800 ;
        RECT 457.200 46.200 458.000 57.800 ;
        RECT 458.800 55.600 459.600 56.400 ;
        RECT 449.200 37.600 450.000 38.400 ;
        RECT 449.200 25.600 450.000 26.400 ;
        RECT 442.800 11.800 443.600 12.600 ;
        RECT 449.300 12.400 449.900 25.600 ;
        RECT 457.200 24.200 458.000 35.800 ;
        RECT 458.900 30.400 459.500 55.600 ;
        RECT 460.400 46.200 461.200 57.800 ;
        RECT 462.000 55.600 462.800 56.400 ;
        RECT 462.100 54.400 462.700 55.600 ;
        RECT 462.000 53.600 462.800 54.400 ;
        RECT 463.600 46.200 464.400 57.800 ;
        RECT 465.200 44.200 466.000 57.800 ;
        RECT 466.800 44.200 467.600 57.800 ;
        RECT 471.600 57.600 472.400 58.400 ;
        RECT 476.500 56.400 477.100 69.600 ;
        RECT 476.400 55.600 477.200 56.400 ;
        RECT 476.400 53.600 477.200 54.400 ;
        RECT 473.200 51.600 474.000 52.400 ;
        RECT 465.200 41.600 466.000 42.400 ;
        RECT 458.800 29.600 459.600 30.400 ;
        RECT 465.300 30.200 465.900 41.600 ;
        RECT 465.200 29.400 466.000 30.200 ;
        RECT 458.800 25.600 459.600 26.400 ;
        RECT 442.900 11.700 443.500 11.800 ;
        RECT 449.200 11.600 450.000 12.400 ;
        RECT 450.800 6.200 451.600 17.800 ;
        RECT 458.900 12.400 459.500 25.600 ;
        RECT 466.800 24.200 467.600 35.800 ;
        RECT 468.400 27.600 469.200 28.400 ;
        RECT 468.500 26.400 469.100 27.600 ;
        RECT 468.400 25.600 469.200 26.400 ;
        RECT 470.000 26.200 470.800 31.800 ;
        RECT 471.600 25.600 472.400 26.400 ;
        RECT 471.700 24.400 472.300 25.600 ;
        RECT 471.600 23.600 472.400 24.400 ;
        RECT 473.300 12.400 473.900 51.600 ;
        RECT 478.100 46.400 478.700 69.600 ;
        RECT 482.800 67.600 483.600 68.400 ;
        RECT 487.600 67.600 488.400 68.400 ;
        RECT 482.900 66.400 483.500 67.600 ;
        RECT 482.800 65.600 483.600 66.400 ;
        RECT 479.600 63.600 480.400 64.400 ;
        RECT 479.700 50.400 480.300 63.600 ;
        RECT 487.700 60.400 488.300 67.600 ;
        RECT 487.600 59.600 488.400 60.400 ;
        RECT 487.700 52.400 488.300 59.600 ;
        RECT 489.300 52.400 489.900 69.700 ;
        RECT 490.800 69.600 491.600 70.400 ;
        RECT 492.400 69.600 493.200 70.400 ;
        RECT 494.000 69.600 494.800 70.400 ;
        RECT 497.200 69.600 498.000 70.400 ;
        RECT 502.000 69.600 502.800 70.400 ;
        RECT 490.900 68.400 491.500 69.600 ;
        RECT 490.800 67.600 491.600 68.400 ;
        RECT 494.100 58.400 494.700 69.600 ;
        RECT 502.100 68.400 502.700 69.600 ;
        RECT 503.700 68.400 504.300 75.600 ;
        RECT 505.200 71.600 506.000 72.400 ;
        RECT 502.000 67.600 502.800 68.400 ;
        RECT 503.600 67.600 504.400 68.400 ;
        RECT 503.600 65.600 504.400 66.400 ;
        RECT 497.200 63.600 498.000 64.400 ;
        RECT 494.000 57.600 494.800 58.400 ;
        RECT 492.400 55.600 493.200 56.400 ;
        RECT 492.500 52.400 493.100 55.600 ;
        RECT 497.300 54.400 497.900 63.600 ;
        RECT 500.400 57.600 501.200 58.400 ;
        RECT 500.500 54.400 501.100 57.600 ;
        RECT 503.700 54.400 504.300 65.600 ;
        RECT 505.200 63.600 506.000 64.400 ;
        RECT 497.200 53.600 498.000 54.400 ;
        RECT 500.400 53.600 501.200 54.400 ;
        RECT 502.000 53.600 502.800 54.400 ;
        RECT 503.600 53.600 504.400 54.400 ;
        RECT 482.800 51.600 483.600 52.400 ;
        RECT 484.400 51.600 485.200 52.400 ;
        RECT 487.600 51.600 488.400 52.400 ;
        RECT 489.200 51.600 490.000 52.400 ;
        RECT 492.400 51.600 493.200 52.400 ;
        RECT 497.200 51.600 498.000 52.400 ;
        RECT 479.600 49.600 480.400 50.400 ;
        RECT 478.000 45.600 478.800 46.400 ;
        RECT 478.000 43.600 478.800 44.400 ;
        RECT 476.400 33.600 477.200 34.400 ;
        RECT 476.500 30.400 477.100 33.600 ;
        RECT 478.100 32.300 478.700 43.600 ;
        RECT 479.700 34.400 480.300 49.600 ;
        RECT 487.700 38.400 488.300 51.600 ;
        RECT 497.300 44.400 497.900 51.600 ;
        RECT 497.200 43.600 498.000 44.400 ;
        RECT 482.800 37.600 483.600 38.400 ;
        RECT 487.600 37.600 488.400 38.400 ;
        RECT 479.600 33.600 480.400 34.400 ;
        RECT 479.600 32.300 480.400 32.400 ;
        RECT 478.100 31.700 480.400 32.300 ;
        RECT 479.600 31.600 480.400 31.700 ;
        RECT 476.400 29.600 477.200 30.400 ;
        RECT 490.800 29.600 491.600 30.400 ;
        RECT 482.800 25.600 483.600 26.400 ;
        RECT 479.600 23.600 480.400 24.400 ;
        RECT 458.800 11.600 459.600 12.400 ;
        RECT 462.000 11.600 462.800 12.400 ;
        RECT 473.200 11.600 474.000 12.400 ;
        RECT 474.800 4.200 475.600 17.800 ;
        RECT 476.400 4.200 477.200 17.800 ;
        RECT 478.000 6.200 478.800 17.800 ;
        RECT 479.700 14.400 480.300 23.600 ;
        RECT 479.600 13.600 480.400 14.400 ;
        RECT 481.200 6.200 482.000 17.800 ;
        RECT 482.900 16.400 483.500 25.600 ;
        RECT 482.800 15.600 483.600 16.400 ;
        RECT 484.400 6.200 485.200 17.800 ;
        RECT 486.000 4.200 486.800 17.800 ;
        RECT 487.600 4.200 488.400 17.800 ;
        RECT 489.200 4.200 490.000 17.800 ;
        RECT 490.900 12.400 491.500 29.600 ;
        RECT 492.400 24.200 493.200 37.800 ;
        RECT 494.000 24.200 494.800 37.800 ;
        RECT 495.600 24.200 496.400 37.800 ;
        RECT 497.200 24.200 498.000 35.800 ;
        RECT 498.800 25.600 499.600 26.400 ;
        RECT 498.800 23.600 499.600 24.400 ;
        RECT 500.400 24.200 501.200 35.800 ;
        RECT 502.100 28.400 502.700 53.600 ;
        RECT 505.300 50.400 505.900 63.600 ;
        RECT 506.900 58.400 507.500 75.600 ;
        RECT 510.000 73.600 510.800 74.400 ;
        RECT 508.400 71.600 509.200 72.400 ;
        RECT 510.100 68.400 510.700 73.600 ;
        RECT 510.000 67.600 510.800 68.400 ;
        RECT 514.800 67.600 515.600 68.400 ;
        RECT 516.200 67.600 517.200 68.400 ;
        RECT 511.600 63.600 512.400 64.400 ;
        RECT 506.800 57.600 507.600 58.400 ;
        RECT 506.900 54.400 507.500 57.600 ;
        RECT 511.700 56.300 512.300 63.600 ;
        RECT 514.900 58.400 515.500 67.600 ;
        RECT 514.800 57.600 515.600 58.400 ;
        RECT 514.900 56.400 515.500 57.600 ;
        RECT 511.700 55.700 513.900 56.300 ;
        RECT 506.800 53.600 507.600 54.400 ;
        RECT 511.600 53.600 512.400 54.400 ;
        RECT 508.400 51.600 509.200 52.400 ;
        RECT 510.000 51.600 510.800 52.400 ;
        RECT 505.200 49.600 506.000 50.400 ;
        RECT 502.000 27.600 502.800 28.400 ;
        RECT 502.000 23.600 502.800 24.400 ;
        RECT 503.600 24.200 504.400 35.800 ;
        RECT 505.200 24.200 506.000 37.800 ;
        RECT 506.800 24.200 507.600 37.800 ;
        RECT 510.100 30.400 510.700 51.600 ;
        RECT 513.300 50.400 513.900 55.700 ;
        RECT 514.800 55.600 515.600 56.400 ;
        RECT 513.200 49.600 514.000 50.400 ;
        RECT 521.200 49.600 522.000 50.400 ;
        RECT 519.600 37.600 520.400 38.400 ;
        RECT 518.000 31.600 518.800 32.400 ;
        RECT 518.100 30.400 518.700 31.600 ;
        RECT 510.000 29.600 510.800 30.400 ;
        RECT 518.000 29.600 518.800 30.400 ;
        RECT 498.900 18.400 499.500 23.600 ;
        RECT 498.800 17.600 499.600 18.400 ;
        RECT 502.100 16.400 502.700 23.600 ;
        RECT 503.600 21.600 504.400 22.400 ;
        RECT 503.700 18.400 504.300 21.600 ;
        RECT 503.600 17.600 504.400 18.400 ;
        RECT 502.000 15.600 502.800 16.400 ;
        RECT 510.100 12.400 510.700 29.600 ;
        RECT 518.000 27.600 518.800 28.400 ;
        RECT 490.800 11.600 491.600 12.400 ;
        RECT 510.000 11.600 510.800 12.400 ;
        RECT 513.200 4.200 514.000 17.800 ;
        RECT 514.800 4.200 515.600 17.800 ;
        RECT 516.400 6.200 517.200 17.800 ;
        RECT 518.100 14.400 518.700 27.600 ;
        RECT 521.300 26.400 521.900 49.600 ;
        RECT 522.900 30.400 523.500 171.600 ;
        RECT 524.400 164.200 525.200 177.800 ;
        RECT 526.000 164.200 526.800 177.800 ;
        RECT 527.600 164.200 528.400 177.800 ;
        RECT 529.200 166.200 530.000 177.800 ;
        RECT 530.900 176.400 531.500 189.600 ;
        RECT 534.000 184.200 534.800 195.800 ;
        RECT 540.500 188.400 541.100 211.600 ;
        RECT 542.100 198.400 542.700 213.600 ;
        RECT 542.000 197.600 542.800 198.400 ;
        RECT 542.000 189.600 542.800 190.400 ;
        RECT 540.400 187.600 541.200 188.400 ;
        RECT 538.800 183.600 539.600 184.400 ;
        RECT 538.900 180.400 539.500 183.600 ;
        RECT 538.800 179.600 539.600 180.400 ;
        RECT 530.800 175.600 531.600 176.400 ;
        RECT 532.400 166.200 533.200 177.800 ;
        RECT 534.000 173.600 534.800 174.400 ;
        RECT 524.400 149.600 525.200 150.400 ;
        RECT 524.500 146.400 525.100 149.600 ;
        RECT 524.400 145.600 525.200 146.400 ;
        RECT 526.000 146.200 526.800 151.800 ;
        RECT 529.200 144.200 530.000 155.800 ;
        RECT 530.900 150.200 531.500 150.300 ;
        RECT 530.800 149.400 531.600 150.200 ;
        RECT 530.900 144.400 531.500 149.400 ;
        RECT 532.400 147.600 533.200 148.400 ;
        RECT 530.800 143.600 531.600 144.400 ;
        RECT 526.000 124.200 526.800 137.800 ;
        RECT 527.600 124.200 528.400 137.800 ;
        RECT 529.200 124.200 530.000 137.800 ;
        RECT 530.800 126.200 531.600 137.800 ;
        RECT 532.500 136.400 533.100 147.600 ;
        RECT 534.100 140.400 534.700 173.600 ;
        RECT 535.600 166.200 536.400 177.800 ;
        RECT 537.200 164.200 538.000 177.800 ;
        RECT 538.800 164.200 539.600 177.800 ;
        RECT 540.500 174.300 541.100 187.600 ;
        RECT 542.100 184.400 542.700 189.600 ;
        RECT 542.000 183.600 542.800 184.400 ;
        RECT 540.500 173.700 542.700 174.300 ;
        RECT 538.800 144.200 539.600 155.800 ;
        RECT 535.600 141.600 536.400 142.400 ;
        RECT 534.000 139.600 534.800 140.400 ;
        RECT 532.400 135.600 533.200 136.400 ;
        RECT 532.500 124.300 533.100 135.600 ;
        RECT 534.000 126.200 534.800 137.800 ;
        RECT 535.700 134.400 536.300 141.600 ;
        RECT 535.600 133.600 536.400 134.400 ;
        RECT 537.200 126.200 538.000 137.800 ;
        RECT 532.500 123.700 534.700 124.300 ;
        RECT 538.800 124.200 539.600 137.800 ;
        RECT 540.400 124.200 541.200 137.800 ;
        RECT 527.600 104.200 528.400 117.800 ;
        RECT 529.200 104.200 530.000 117.800 ;
        RECT 530.800 104.200 531.600 117.800 ;
        RECT 532.400 104.200 533.200 115.800 ;
        RECT 534.100 106.400 534.700 123.700 ;
        RECT 542.100 120.400 542.700 173.700 ;
        RECT 543.700 158.400 544.300 243.600 ;
        RECT 545.300 230.400 545.900 259.700 ;
        RECT 546.900 258.400 547.500 363.600 ;
        RECT 548.500 344.400 549.100 375.600 ;
        RECT 548.400 343.600 549.200 344.400 ;
        RECT 548.400 331.600 549.200 332.400 ;
        RECT 546.800 257.600 547.600 258.400 ;
        RECT 546.800 250.200 547.600 255.800 ;
        RECT 548.500 244.400 549.100 331.600 ;
        RECT 548.400 243.600 549.200 244.400 ;
        RECT 545.200 229.600 546.000 230.400 ;
        RECT 546.800 229.600 547.600 230.400 ;
        RECT 546.900 226.400 547.500 229.600 ;
        RECT 546.800 225.600 547.600 226.400 ;
        RECT 550.000 207.600 550.800 208.400 ;
        RECT 546.800 191.600 547.600 192.400 ;
        RECT 550.100 190.400 550.700 207.600 ;
        RECT 550.000 189.600 550.800 190.400 ;
        RECT 550.100 188.400 550.700 189.600 ;
        RECT 550.000 187.600 550.800 188.400 ;
        RECT 543.600 157.600 544.400 158.400 ;
        RECT 545.200 151.600 546.000 152.400 ;
        RECT 545.300 150.400 545.900 151.600 ;
        RECT 545.200 149.600 546.000 150.400 ;
        RECT 543.600 131.600 544.400 132.400 ;
        RECT 542.000 119.600 542.800 120.400 ;
        RECT 534.000 105.600 534.800 106.400 ;
        RECT 526.000 91.600 526.800 92.400 ;
        RECT 527.600 84.200 528.400 97.800 ;
        RECT 529.200 84.200 530.000 97.800 ;
        RECT 530.800 84.200 531.600 97.800 ;
        RECT 532.400 86.200 533.200 97.800 ;
        RECT 534.100 96.400 534.700 105.600 ;
        RECT 535.600 104.200 536.400 115.800 ;
        RECT 537.200 107.600 538.000 108.400 ;
        RECT 537.300 106.400 537.900 107.600 ;
        RECT 537.200 105.600 538.000 106.400 ;
        RECT 538.800 104.200 539.600 115.800 ;
        RECT 540.400 104.200 541.200 117.800 ;
        RECT 542.000 104.200 542.800 117.800 ;
        RECT 543.700 110.400 544.300 131.600 ;
        RECT 543.600 109.600 544.400 110.400 ;
        RECT 545.200 109.600 546.000 110.400 ;
        RECT 537.200 99.600 538.000 100.400 ;
        RECT 534.000 95.600 534.800 96.400 ;
        RECT 534.100 84.300 534.700 95.600 ;
        RECT 535.600 86.200 536.400 97.800 ;
        RECT 537.300 94.400 537.900 99.600 ;
        RECT 537.200 93.600 538.000 94.400 ;
        RECT 538.800 86.200 539.600 97.800 ;
        RECT 532.500 83.700 534.700 84.300 ;
        RECT 540.400 84.200 541.200 97.800 ;
        RECT 542.000 84.200 542.800 97.800 ;
        RECT 545.300 92.400 545.900 109.600 ;
        RECT 545.200 91.600 546.000 92.400 ;
        RECT 526.000 64.200 526.800 77.800 ;
        RECT 527.600 64.200 528.400 77.800 ;
        RECT 529.200 64.200 530.000 77.800 ;
        RECT 530.800 64.200 531.600 75.800 ;
        RECT 532.500 66.400 533.100 83.700 ;
        RECT 545.300 82.400 545.900 91.600 ;
        RECT 542.000 81.600 542.800 82.400 ;
        RECT 545.200 81.600 546.000 82.400 ;
        RECT 532.400 65.600 533.200 66.400 ;
        RECT 532.500 62.300 533.100 65.600 ;
        RECT 534.000 64.200 534.800 75.800 ;
        RECT 535.600 67.600 536.400 68.400 ;
        RECT 535.700 66.400 536.300 67.600 ;
        RECT 535.600 65.600 536.400 66.400 ;
        RECT 537.200 64.200 538.000 75.800 ;
        RECT 538.800 64.200 539.600 77.800 ;
        RECT 540.400 64.200 541.200 77.800 ;
        RECT 542.100 70.400 542.700 81.600 ;
        RECT 542.000 69.600 542.800 70.400 ;
        RECT 530.900 61.700 533.100 62.300 ;
        RECT 524.400 44.200 525.200 57.800 ;
        RECT 526.000 44.200 526.800 57.800 ;
        RECT 527.600 44.200 528.400 57.800 ;
        RECT 529.200 46.200 530.000 57.800 ;
        RECT 530.900 56.400 531.500 61.700 ;
        RECT 530.800 55.600 531.600 56.400 ;
        RECT 530.900 50.400 531.500 55.600 ;
        RECT 530.800 49.600 531.600 50.400 ;
        RECT 532.400 46.200 533.200 57.800 ;
        RECT 534.000 53.600 534.800 54.400 ;
        RECT 534.000 51.600 534.800 52.400 ;
        RECT 535.600 46.200 536.400 57.800 ;
        RECT 537.200 44.200 538.000 57.800 ;
        RECT 538.800 44.200 539.600 57.800 ;
        RECT 542.100 52.400 542.700 69.600 ;
        RECT 542.000 51.600 542.800 52.400 ;
        RECT 546.800 49.600 547.600 50.400 ;
        RECT 546.900 38.400 547.500 49.600 ;
        RECT 530.800 37.600 531.600 38.400 ;
        RECT 546.800 37.600 547.600 38.400 ;
        RECT 527.600 33.600 528.400 34.400 ;
        RECT 527.700 30.400 528.300 33.600 ;
        RECT 532.400 31.600 533.200 32.400 ;
        RECT 532.500 30.400 533.100 31.600 ;
        RECT 522.800 29.600 523.600 30.400 ;
        RECT 524.400 29.600 525.200 30.400 ;
        RECT 527.600 29.600 528.400 30.400 ;
        RECT 532.400 29.600 533.200 30.400 ;
        RECT 521.200 25.600 522.000 26.400 ;
        RECT 518.000 13.600 518.800 14.400 ;
        RECT 519.600 6.200 520.400 17.800 ;
        RECT 521.300 16.400 521.900 25.600 ;
        RECT 521.200 15.600 522.000 16.400 ;
        RECT 522.800 6.200 523.600 17.800 ;
        RECT 524.400 4.200 525.200 17.800 ;
        RECT 526.000 4.200 526.800 17.800 ;
        RECT 527.600 4.200 528.400 17.800 ;
        RECT 545.200 11.600 546.000 12.400 ;
      LAYER via2 ;
        RECT 105.200 229.600 106.000 230.400 ;
        RECT 129.200 191.600 130.000 192.400 ;
        RECT 297.200 349.600 298.000 350.400 ;
        RECT 68.400 11.600 69.200 12.400 ;
        RECT 183.600 131.600 184.400 132.400 ;
        RECT 122.800 51.600 123.600 52.400 ;
        RECT 116.400 11.600 117.200 12.400 ;
        RECT 270.000 267.600 270.800 268.400 ;
        RECT 268.400 189.600 269.200 190.400 ;
        RECT 311.600 231.600 312.400 232.400 ;
        RECT 426.800 373.600 427.600 374.400 ;
        RECT 438.000 371.600 438.800 372.400 ;
        RECT 295.600 149.600 296.400 150.400 ;
        RECT 274.800 109.600 275.600 110.400 ;
        RECT 236.400 51.600 237.200 52.400 ;
        RECT 434.800 253.600 435.600 254.400 ;
        RECT 378.800 189.600 379.600 190.400 ;
        RECT 290.800 11.600 291.600 12.400 ;
        RECT 511.600 251.600 512.400 252.400 ;
        RECT 497.200 227.600 498.000 228.400 ;
        RECT 324.400 29.600 325.200 30.400 ;
        RECT 516.400 67.600 517.200 68.400 ;
      LAYER metal3 ;
        RECT 196.400 378.300 197.200 378.400 ;
        RECT 218.800 378.300 219.600 378.400 ;
        RECT 196.400 377.700 219.600 378.300 ;
        RECT 196.400 377.600 197.200 377.700 ;
        RECT 218.800 377.600 219.600 377.700 ;
        RECT 327.600 378.300 328.400 378.400 ;
        RECT 388.400 378.300 389.200 378.400 ;
        RECT 327.600 377.700 389.200 378.300 ;
        RECT 327.600 377.600 328.400 377.700 ;
        RECT 388.400 377.600 389.200 377.700 ;
        RECT 18.800 376.300 19.600 376.400 ;
        RECT 52.400 376.300 53.200 376.400 ;
        RECT 89.200 376.300 90.000 376.400 ;
        RECT 18.800 375.700 90.000 376.300 ;
        RECT 18.800 375.600 19.600 375.700 ;
        RECT 52.400 375.600 53.200 375.700 ;
        RECT 89.200 375.600 90.000 375.700 ;
        RECT 134.000 376.300 134.800 376.400 ;
        RECT 249.200 376.300 250.000 376.400 ;
        RECT 134.000 375.700 250.000 376.300 ;
        RECT 134.000 375.600 134.800 375.700 ;
        RECT 249.200 375.600 250.000 375.700 ;
        RECT 273.200 376.300 274.000 376.400 ;
        RECT 302.000 376.300 302.800 376.400 ;
        RECT 273.200 375.700 302.800 376.300 ;
        RECT 273.200 375.600 274.000 375.700 ;
        RECT 302.000 375.600 302.800 375.700 ;
        RECT 314.800 376.300 315.600 376.400 ;
        RECT 330.800 376.300 331.600 376.400 ;
        RECT 314.800 375.700 331.600 376.300 ;
        RECT 314.800 375.600 315.600 375.700 ;
        RECT 330.800 375.600 331.600 375.700 ;
        RECT 335.600 376.300 336.400 376.400 ;
        RECT 342.000 376.300 342.800 376.400 ;
        RECT 335.600 375.700 342.800 376.300 ;
        RECT 335.600 375.600 336.400 375.700 ;
        RECT 342.000 375.600 342.800 375.700 ;
        RECT 410.800 376.300 411.600 376.400 ;
        RECT 454.000 376.300 454.800 376.400 ;
        RECT 410.800 375.700 454.800 376.300 ;
        RECT 410.800 375.600 411.600 375.700 ;
        RECT 454.000 375.600 454.800 375.700 ;
        RECT 487.600 376.300 488.400 376.400 ;
        RECT 529.200 376.300 530.000 376.400 ;
        RECT 487.600 375.700 530.000 376.300 ;
        RECT 487.600 375.600 488.400 375.700 ;
        RECT 529.200 375.600 530.000 375.700 ;
        RECT 22.000 374.300 22.800 374.400 ;
        RECT 26.800 374.300 27.600 374.400 ;
        RECT 22.000 373.700 27.600 374.300 ;
        RECT 22.000 373.600 22.800 373.700 ;
        RECT 26.800 373.600 27.600 373.700 ;
        RECT 92.400 374.300 93.200 374.400 ;
        RECT 236.400 374.300 237.200 374.400 ;
        RECT 92.400 373.700 237.200 374.300 ;
        RECT 92.400 373.600 93.200 373.700 ;
        RECT 236.400 373.600 237.200 373.700 ;
        RECT 242.800 374.300 243.600 374.400 ;
        RECT 247.600 374.300 248.400 374.400 ;
        RECT 242.800 373.700 248.400 374.300 ;
        RECT 242.800 373.600 243.600 373.700 ;
        RECT 247.600 373.600 248.400 373.700 ;
        RECT 295.600 374.300 296.400 374.400 ;
        RECT 300.400 374.300 301.200 374.400 ;
        RECT 295.600 373.700 301.200 374.300 ;
        RECT 295.600 373.600 296.400 373.700 ;
        RECT 300.400 373.600 301.200 373.700 ;
        RECT 319.600 374.300 320.400 374.400 ;
        RECT 337.200 374.300 338.000 374.400 ;
        RECT 319.600 373.700 338.000 374.300 ;
        RECT 319.600 373.600 320.400 373.700 ;
        RECT 337.200 373.600 338.000 373.700 ;
        RECT 340.400 374.300 341.200 374.400 ;
        RECT 346.800 374.300 347.600 374.400 ;
        RECT 340.400 373.700 347.600 374.300 ;
        RECT 340.400 373.600 341.200 373.700 ;
        RECT 346.800 373.600 347.600 373.700 ;
        RECT 359.600 374.300 360.400 374.400 ;
        RECT 361.200 374.300 362.000 374.400 ;
        RECT 359.600 373.700 362.000 374.300 ;
        RECT 359.600 373.600 360.400 373.700 ;
        RECT 361.200 373.600 362.000 373.700 ;
        RECT 386.800 374.300 387.600 374.400 ;
        RECT 393.200 374.300 394.000 374.400 ;
        RECT 426.800 374.300 427.600 374.400 ;
        RECT 386.800 373.700 427.600 374.300 ;
        RECT 386.800 373.600 387.600 373.700 ;
        RECT 393.200 373.600 394.000 373.700 ;
        RECT 426.800 373.600 427.600 373.700 ;
        RECT 446.000 374.300 446.800 374.400 ;
        RECT 484.400 374.300 485.200 374.400 ;
        RECT 446.000 373.700 485.200 374.300 ;
        RECT 446.000 373.600 446.800 373.700 ;
        RECT 484.400 373.600 485.200 373.700 ;
        RECT 502.000 374.300 502.800 374.400 ;
        RECT 506.800 374.300 507.600 374.400 ;
        RECT 502.000 373.700 507.600 374.300 ;
        RECT 502.000 373.600 502.800 373.700 ;
        RECT 506.800 373.600 507.600 373.700 ;
        RECT 508.400 374.300 509.200 374.400 ;
        RECT 532.400 374.300 533.200 374.400 ;
        RECT 508.400 373.700 533.200 374.300 ;
        RECT 508.400 373.600 509.200 373.700 ;
        RECT 532.400 373.600 533.200 373.700 ;
        RECT 31.600 372.300 32.400 372.400 ;
        RECT 38.000 372.300 38.800 372.400 ;
        RECT 31.600 371.700 38.800 372.300 ;
        RECT 31.600 371.600 32.400 371.700 ;
        RECT 38.000 371.600 38.800 371.700 ;
        RECT 161.200 372.300 162.000 372.400 ;
        RECT 175.600 372.300 176.400 372.400 ;
        RECT 161.200 371.700 176.400 372.300 ;
        RECT 161.200 371.600 162.000 371.700 ;
        RECT 175.600 371.600 176.400 371.700 ;
        RECT 228.400 372.300 229.200 372.400 ;
        RECT 234.800 372.300 235.600 372.400 ;
        RECT 246.000 372.300 246.800 372.400 ;
        RECT 298.800 372.300 299.600 372.400 ;
        RECT 228.400 371.700 299.600 372.300 ;
        RECT 228.400 371.600 229.200 371.700 ;
        RECT 234.800 371.600 235.600 371.700 ;
        RECT 246.000 371.600 246.800 371.700 ;
        RECT 298.800 371.600 299.600 371.700 ;
        RECT 310.000 372.300 310.800 372.400 ;
        RECT 314.800 372.300 315.600 372.400 ;
        RECT 310.000 371.700 315.600 372.300 ;
        RECT 310.000 371.600 310.800 371.700 ;
        RECT 314.800 371.600 315.600 371.700 ;
        RECT 318.000 372.300 318.800 372.400 ;
        RECT 322.800 372.300 323.600 372.400 ;
        RECT 318.000 371.700 323.600 372.300 ;
        RECT 318.000 371.600 318.800 371.700 ;
        RECT 322.800 371.600 323.600 371.700 ;
        RECT 337.200 372.300 338.000 372.400 ;
        RECT 345.200 372.300 346.000 372.400 ;
        RECT 382.000 372.300 382.800 372.400 ;
        RECT 337.200 371.700 382.800 372.300 ;
        RECT 337.200 371.600 338.000 371.700 ;
        RECT 345.200 371.600 346.000 371.700 ;
        RECT 382.000 371.600 382.800 371.700 ;
        RECT 391.600 372.300 392.400 372.400 ;
        RECT 438.000 372.300 438.800 372.400 ;
        RECT 391.600 371.700 438.800 372.300 ;
        RECT 391.600 371.600 392.400 371.700 ;
        RECT 438.000 371.600 438.800 371.700 ;
        RECT 463.600 372.300 464.400 372.400 ;
        RECT 474.800 372.300 475.600 372.400 ;
        RECT 463.600 371.700 475.600 372.300 ;
        RECT 463.600 371.600 464.400 371.700 ;
        RECT 474.800 371.600 475.600 371.700 ;
        RECT 495.600 372.300 496.400 372.400 ;
        RECT 521.200 372.300 522.000 372.400 ;
        RECT 495.600 371.700 522.000 372.300 ;
        RECT 495.600 371.600 496.400 371.700 ;
        RECT 521.200 371.600 522.000 371.700 ;
        RECT 529.200 372.300 530.000 372.400 ;
        RECT 532.400 372.300 533.200 372.400 ;
        RECT 529.200 371.700 533.200 372.300 ;
        RECT 529.200 371.600 530.000 371.700 ;
        RECT 532.400 371.600 533.200 371.700 ;
        RECT 172.400 370.300 173.200 370.400 ;
        RECT 186.800 370.300 187.600 370.400 ;
        RECT 172.400 369.700 187.600 370.300 ;
        RECT 172.400 369.600 173.200 369.700 ;
        RECT 186.800 369.600 187.600 369.700 ;
        RECT 215.600 370.300 216.400 370.400 ;
        RECT 222.000 370.300 222.800 370.400 ;
        RECT 215.600 369.700 222.800 370.300 ;
        RECT 215.600 369.600 216.400 369.700 ;
        RECT 222.000 369.600 222.800 369.700 ;
        RECT 226.800 370.300 227.600 370.400 ;
        RECT 233.200 370.300 234.000 370.400 ;
        RECT 244.400 370.300 245.200 370.400 ;
        RECT 297.200 370.300 298.000 370.400 ;
        RECT 327.600 370.300 328.400 370.400 ;
        RECT 226.800 369.700 328.400 370.300 ;
        RECT 226.800 369.600 227.600 369.700 ;
        RECT 233.200 369.600 234.000 369.700 ;
        RECT 244.400 369.600 245.200 369.700 ;
        RECT 297.200 369.600 298.000 369.700 ;
        RECT 327.600 369.600 328.400 369.700 ;
        RECT 329.200 370.300 330.000 370.400 ;
        RECT 334.000 370.300 334.800 370.400 ;
        RECT 329.200 369.700 334.800 370.300 ;
        RECT 329.200 369.600 330.000 369.700 ;
        RECT 334.000 369.600 334.800 369.700 ;
        RECT 505.200 370.300 506.000 370.400 ;
        RECT 510.000 370.300 510.800 370.400 ;
        RECT 505.200 369.700 510.800 370.300 ;
        RECT 505.200 369.600 506.000 369.700 ;
        RECT 510.000 369.600 510.800 369.700 ;
        RECT 73.200 368.300 74.000 368.400 ;
        RECT 230.000 368.300 230.800 368.400 ;
        RECT 73.200 367.700 230.800 368.300 ;
        RECT 73.200 367.600 74.000 367.700 ;
        RECT 230.000 367.600 230.800 367.700 ;
        RECT 233.200 368.300 234.000 368.400 ;
        RECT 236.400 368.300 237.200 368.400 ;
        RECT 233.200 367.700 237.200 368.300 ;
        RECT 233.200 367.600 234.000 367.700 ;
        RECT 236.400 367.600 237.200 367.700 ;
        RECT 250.800 368.300 251.600 368.400 ;
        RECT 313.200 368.300 314.000 368.400 ;
        RECT 332.400 368.300 333.200 368.400 ;
        RECT 250.800 367.700 314.000 368.300 ;
        RECT 250.800 367.600 251.600 367.700 ;
        RECT 313.200 367.600 314.000 367.700 ;
        RECT 319.700 367.700 333.200 368.300 ;
        RECT 92.400 366.300 93.200 366.400 ;
        RECT 114.800 366.300 115.600 366.400 ;
        RECT 239.600 366.300 240.400 366.400 ;
        RECT 92.400 365.700 240.400 366.300 ;
        RECT 92.400 365.600 93.200 365.700 ;
        RECT 114.800 365.600 115.600 365.700 ;
        RECT 239.600 365.600 240.400 365.700 ;
        RECT 241.200 366.300 242.000 366.400 ;
        RECT 252.400 366.300 253.200 366.400 ;
        RECT 241.200 365.700 253.200 366.300 ;
        RECT 241.200 365.600 242.000 365.700 ;
        RECT 252.400 365.600 253.200 365.700 ;
        RECT 255.600 366.300 256.400 366.400 ;
        RECT 305.200 366.300 306.000 366.400 ;
        RECT 308.400 366.300 309.200 366.400 ;
        RECT 255.600 365.700 309.200 366.300 ;
        RECT 255.600 365.600 256.400 365.700 ;
        RECT 305.200 365.600 306.000 365.700 ;
        RECT 308.400 365.600 309.200 365.700 ;
        RECT 311.600 366.300 312.400 366.400 ;
        RECT 319.700 366.300 320.300 367.700 ;
        RECT 332.400 367.600 333.200 367.700 ;
        RECT 366.000 368.300 366.800 368.400 ;
        RECT 388.400 368.300 389.200 368.400 ;
        RECT 366.000 367.700 389.200 368.300 ;
        RECT 366.000 367.600 366.800 367.700 ;
        RECT 388.400 367.600 389.200 367.700 ;
        RECT 390.000 368.300 390.800 368.400 ;
        RECT 407.600 368.300 408.400 368.400 ;
        RECT 390.000 367.700 408.400 368.300 ;
        RECT 390.000 367.600 390.800 367.700 ;
        RECT 407.600 367.600 408.400 367.700 ;
        RECT 506.800 368.300 507.600 368.400 ;
        RECT 526.000 368.300 526.800 368.400 ;
        RECT 506.800 367.700 526.800 368.300 ;
        RECT 506.800 367.600 507.600 367.700 ;
        RECT 526.000 367.600 526.800 367.700 ;
        RECT 311.600 365.700 320.300 366.300 ;
        RECT 321.200 366.300 322.000 366.400 ;
        RECT 351.600 366.300 352.400 366.400 ;
        RECT 399.600 366.300 400.400 366.400 ;
        RECT 321.200 365.700 400.400 366.300 ;
        RECT 311.600 365.600 312.400 365.700 ;
        RECT 321.200 365.600 322.000 365.700 ;
        RECT 351.600 365.600 352.400 365.700 ;
        RECT 399.600 365.600 400.400 365.700 ;
        RECT 68.400 364.300 69.200 364.400 ;
        RECT 71.600 364.300 72.400 364.400 ;
        RECT 68.400 363.700 72.400 364.300 ;
        RECT 68.400 363.600 69.200 363.700 ;
        RECT 71.600 363.600 72.400 363.700 ;
        RECT 218.800 364.300 219.600 364.400 ;
        RECT 246.000 364.300 246.800 364.400 ;
        RECT 218.800 363.700 246.800 364.300 ;
        RECT 218.800 363.600 219.600 363.700 ;
        RECT 246.000 363.600 246.800 363.700 ;
        RECT 254.000 364.300 254.800 364.400 ;
        RECT 292.400 364.300 293.200 364.400 ;
        RECT 254.000 363.700 293.200 364.300 ;
        RECT 254.000 363.600 254.800 363.700 ;
        RECT 292.400 363.600 293.200 363.700 ;
        RECT 324.400 364.300 325.200 364.400 ;
        RECT 364.400 364.300 365.200 364.400 ;
        RECT 410.800 364.300 411.600 364.400 ;
        RECT 324.400 363.700 411.600 364.300 ;
        RECT 324.400 363.600 325.200 363.700 ;
        RECT 364.400 363.600 365.200 363.700 ;
        RECT 410.800 363.600 411.600 363.700 ;
        RECT 193.200 362.300 194.000 362.400 ;
        RECT 199.600 362.300 200.400 362.400 ;
        RECT 193.200 361.700 200.400 362.300 ;
        RECT 193.200 361.600 194.000 361.700 ;
        RECT 199.600 361.600 200.400 361.700 ;
        RECT 298.800 362.300 299.600 362.400 ;
        RECT 306.800 362.300 307.600 362.400 ;
        RECT 361.200 362.300 362.000 362.400 ;
        RECT 298.800 361.700 362.000 362.300 ;
        RECT 298.800 361.600 299.600 361.700 ;
        RECT 306.800 361.600 307.600 361.700 ;
        RECT 361.200 361.600 362.000 361.700 ;
        RECT 369.200 362.300 370.000 362.400 ;
        RECT 390.000 362.300 390.800 362.400 ;
        RECT 369.200 361.700 390.800 362.300 ;
        RECT 369.200 361.600 370.000 361.700 ;
        RECT 390.000 361.600 390.800 361.700 ;
        RECT 391.600 362.300 392.400 362.400 ;
        RECT 394.800 362.300 395.600 362.400 ;
        RECT 412.400 362.300 413.200 362.400 ;
        RECT 391.600 361.700 395.600 362.300 ;
        RECT 391.600 361.600 392.400 361.700 ;
        RECT 394.800 361.600 395.600 361.700 ;
        RECT 396.500 361.700 413.200 362.300 ;
        RECT 302.000 360.300 302.800 360.400 ;
        RECT 388.400 360.300 389.200 360.400 ;
        RECT 302.000 359.700 389.200 360.300 ;
        RECT 302.000 359.600 302.800 359.700 ;
        RECT 388.400 359.600 389.200 359.700 ;
        RECT 393.200 360.300 394.000 360.400 ;
        RECT 396.500 360.300 397.100 361.700 ;
        RECT 412.400 361.600 413.200 361.700 ;
        RECT 393.200 359.700 397.100 360.300 ;
        RECT 398.000 360.300 398.800 360.400 ;
        RECT 406.000 360.300 406.800 360.400 ;
        RECT 398.000 359.700 406.800 360.300 ;
        RECT 393.200 359.600 394.000 359.700 ;
        RECT 398.000 359.600 398.800 359.700 ;
        RECT 406.000 359.600 406.800 359.700 ;
        RECT 487.600 360.300 488.400 360.400 ;
        RECT 503.600 360.300 504.400 360.400 ;
        RECT 487.600 359.700 504.400 360.300 ;
        RECT 487.600 359.600 488.400 359.700 ;
        RECT 503.600 359.600 504.400 359.700 ;
        RECT 38.000 358.300 38.800 358.400 ;
        RECT 44.400 358.300 45.200 358.400 ;
        RECT 49.200 358.300 50.000 358.400 ;
        RECT 73.200 358.300 74.000 358.400 ;
        RECT 38.000 357.700 74.000 358.300 ;
        RECT 38.000 357.600 38.800 357.700 ;
        RECT 44.400 357.600 45.200 357.700 ;
        RECT 49.200 357.600 50.000 357.700 ;
        RECT 73.200 357.600 74.000 357.700 ;
        RECT 97.200 358.300 98.000 358.400 ;
        RECT 254.000 358.300 254.800 358.400 ;
        RECT 97.200 357.700 254.800 358.300 ;
        RECT 97.200 357.600 98.000 357.700 ;
        RECT 254.000 357.600 254.800 357.700 ;
        RECT 324.400 358.300 325.200 358.400 ;
        RECT 346.800 358.300 347.600 358.400 ;
        RECT 372.400 358.300 373.200 358.400 ;
        RECT 324.400 357.700 373.200 358.300 ;
        RECT 324.400 357.600 325.200 357.700 ;
        RECT 346.800 357.600 347.600 357.700 ;
        RECT 372.400 357.600 373.200 357.700 ;
        RECT 382.000 358.300 382.800 358.400 ;
        RECT 396.400 358.300 397.200 358.400 ;
        RECT 382.000 357.700 397.200 358.300 ;
        RECT 382.000 357.600 382.800 357.700 ;
        RECT 396.400 357.600 397.200 357.700 ;
        RECT 398.000 358.300 398.800 358.400 ;
        RECT 441.200 358.300 442.000 358.400 ;
        RECT 398.000 357.700 442.000 358.300 ;
        RECT 398.000 357.600 398.800 357.700 ;
        RECT 441.200 357.600 442.000 357.700 ;
        RECT 442.800 358.300 443.600 358.400 ;
        RECT 479.600 358.300 480.400 358.400 ;
        RECT 442.800 357.700 480.400 358.300 ;
        RECT 442.800 357.600 443.600 357.700 ;
        RECT 479.600 357.600 480.400 357.700 ;
        RECT 249.200 356.300 250.000 356.400 ;
        RECT 254.000 356.300 254.800 356.400 ;
        RECT 303.600 356.300 304.400 356.400 ;
        RECT 249.200 355.700 304.400 356.300 ;
        RECT 249.200 355.600 250.000 355.700 ;
        RECT 254.000 355.600 254.800 355.700 ;
        RECT 303.600 355.600 304.400 355.700 ;
        RECT 310.000 356.300 310.800 356.400 ;
        RECT 378.800 356.300 379.600 356.400 ;
        RECT 310.000 355.700 379.600 356.300 ;
        RECT 310.000 355.600 310.800 355.700 ;
        RECT 378.800 355.600 379.600 355.700 ;
        RECT 386.800 356.300 387.600 356.400 ;
        RECT 409.200 356.300 410.000 356.400 ;
        RECT 473.200 356.300 474.000 356.400 ;
        RECT 386.800 355.700 410.000 356.300 ;
        RECT 386.800 355.600 387.600 355.700 ;
        RECT 409.200 355.600 410.000 355.700 ;
        RECT 410.900 355.700 474.000 356.300 ;
        RECT 281.200 354.300 282.000 354.400 ;
        RECT 311.600 354.300 312.400 354.400 ;
        RECT 321.200 354.300 322.000 354.400 ;
        RECT 281.200 353.700 322.000 354.300 ;
        RECT 281.200 353.600 282.000 353.700 ;
        RECT 311.600 353.600 312.400 353.700 ;
        RECT 321.200 353.600 322.000 353.700 ;
        RECT 322.800 354.300 323.600 354.400 ;
        RECT 338.800 354.300 339.600 354.400 ;
        RECT 322.800 353.700 339.600 354.300 ;
        RECT 322.800 353.600 323.600 353.700 ;
        RECT 338.800 353.600 339.600 353.700 ;
        RECT 375.600 354.300 376.400 354.400 ;
        RECT 378.800 354.300 379.600 354.400 ;
        RECT 375.600 353.700 379.600 354.300 ;
        RECT 375.600 353.600 376.400 353.700 ;
        RECT 378.800 353.600 379.600 353.700 ;
        RECT 383.600 354.300 384.400 354.400 ;
        RECT 399.600 354.300 400.400 354.400 ;
        RECT 383.600 353.700 400.400 354.300 ;
        RECT 383.600 353.600 384.400 353.700 ;
        RECT 399.600 353.600 400.400 353.700 ;
        RECT 401.200 354.300 402.000 354.400 ;
        RECT 406.000 354.300 406.800 354.400 ;
        RECT 401.200 353.700 406.800 354.300 ;
        RECT 401.200 353.600 402.000 353.700 ;
        RECT 406.000 353.600 406.800 353.700 ;
        RECT 407.600 354.300 408.400 354.400 ;
        RECT 410.900 354.300 411.500 355.700 ;
        RECT 473.200 355.600 474.000 355.700 ;
        RECT 476.400 356.300 477.200 356.400 ;
        RECT 498.800 356.300 499.600 356.400 ;
        RECT 476.400 355.700 499.600 356.300 ;
        RECT 476.400 355.600 477.200 355.700 ;
        RECT 498.800 355.600 499.600 355.700 ;
        RECT 407.600 353.700 411.500 354.300 ;
        RECT 412.400 354.300 413.200 354.400 ;
        RECT 442.800 354.300 443.600 354.400 ;
        RECT 412.400 353.700 443.600 354.300 ;
        RECT 407.600 353.600 408.400 353.700 ;
        RECT 412.400 353.600 413.200 353.700 ;
        RECT 442.800 353.600 443.600 353.700 ;
        RECT 444.400 354.300 445.200 354.400 ;
        RECT 449.200 354.300 450.000 354.400 ;
        RECT 444.400 353.700 450.000 354.300 ;
        RECT 444.400 353.600 445.200 353.700 ;
        RECT 449.200 353.600 450.000 353.700 ;
        RECT 454.000 354.300 454.800 354.400 ;
        RECT 474.800 354.300 475.600 354.400 ;
        RECT 454.000 353.700 475.600 354.300 ;
        RECT 454.000 353.600 454.800 353.700 ;
        RECT 474.800 353.600 475.600 353.700 ;
        RECT 482.800 354.300 483.600 354.400 ;
        RECT 492.400 354.300 493.200 354.400 ;
        RECT 482.800 353.700 493.200 354.300 ;
        RECT 482.800 353.600 483.600 353.700 ;
        RECT 492.400 353.600 493.200 353.700 ;
        RECT 494.000 354.300 494.800 354.400 ;
        RECT 500.400 354.300 501.200 354.400 ;
        RECT 522.800 354.300 523.600 354.400 ;
        RECT 494.000 353.700 523.600 354.300 ;
        RECT 494.000 353.600 494.800 353.700 ;
        RECT 500.400 353.600 501.200 353.700 ;
        RECT 522.800 353.600 523.600 353.700 ;
        RECT 42.800 352.300 43.600 352.400 ;
        RECT 47.600 352.300 48.400 352.400 ;
        RECT 54.000 352.300 54.800 352.400 ;
        RECT 215.600 352.300 216.400 352.400 ;
        RECT 42.800 351.700 216.400 352.300 ;
        RECT 42.800 351.600 43.600 351.700 ;
        RECT 47.600 351.600 48.400 351.700 ;
        RECT 54.000 351.600 54.800 351.700 ;
        RECT 215.600 351.600 216.400 351.700 ;
        RECT 250.800 352.300 251.600 352.400 ;
        RECT 255.600 352.300 256.400 352.400 ;
        RECT 250.800 351.700 256.400 352.300 ;
        RECT 250.800 351.600 251.600 351.700 ;
        RECT 255.600 351.600 256.400 351.700 ;
        RECT 266.800 352.300 267.600 352.400 ;
        RECT 270.000 352.300 270.800 352.400 ;
        RECT 266.800 351.700 270.800 352.300 ;
        RECT 266.800 351.600 267.600 351.700 ;
        RECT 270.000 351.600 270.800 351.700 ;
        RECT 303.600 352.300 304.400 352.400 ;
        RECT 314.800 352.300 315.600 352.400 ;
        RECT 303.600 351.700 315.600 352.300 ;
        RECT 303.600 351.600 304.400 351.700 ;
        RECT 314.800 351.600 315.600 351.700 ;
        RECT 321.200 352.300 322.000 352.400 ;
        RECT 337.200 352.300 338.000 352.400 ;
        RECT 396.400 352.300 397.200 352.400 ;
        RECT 402.800 352.300 403.600 352.400 ;
        RECT 321.200 351.700 403.600 352.300 ;
        RECT 321.200 351.600 322.000 351.700 ;
        RECT 337.200 351.600 338.000 351.700 ;
        RECT 396.400 351.600 397.200 351.700 ;
        RECT 402.800 351.600 403.600 351.700 ;
        RECT 407.600 352.300 408.400 352.400 ;
        RECT 420.400 352.300 421.200 352.400 ;
        RECT 407.600 351.700 421.200 352.300 ;
        RECT 407.600 351.600 408.400 351.700 ;
        RECT 420.400 351.600 421.200 351.700 ;
        RECT 434.800 352.300 435.600 352.400 ;
        RECT 439.600 352.300 440.400 352.400 ;
        RECT 450.800 352.300 451.600 352.400 ;
        RECT 462.000 352.300 462.800 352.400 ;
        RECT 434.800 351.700 462.800 352.300 ;
        RECT 434.800 351.600 435.600 351.700 ;
        RECT 439.600 351.600 440.400 351.700 ;
        RECT 450.800 351.600 451.600 351.700 ;
        RECT 462.000 351.600 462.800 351.700 ;
        RECT 465.200 352.300 466.000 352.400 ;
        RECT 508.400 352.300 509.200 352.400 ;
        RECT 465.200 351.700 509.200 352.300 ;
        RECT 465.200 351.600 466.000 351.700 ;
        RECT 508.400 351.600 509.200 351.700 ;
        RECT 82.800 350.300 83.600 350.400 ;
        RECT 100.400 350.300 101.200 350.400 ;
        RECT 82.800 349.700 101.200 350.300 ;
        RECT 82.800 349.600 83.600 349.700 ;
        RECT 100.400 349.600 101.200 349.700 ;
        RECT 122.800 350.300 123.600 350.400 ;
        RECT 140.400 350.300 141.200 350.400 ;
        RECT 143.600 350.300 144.400 350.400 ;
        RECT 122.800 349.700 144.400 350.300 ;
        RECT 122.800 349.600 123.600 349.700 ;
        RECT 140.400 349.600 141.200 349.700 ;
        RECT 143.600 349.600 144.400 349.700 ;
        RECT 206.000 350.300 206.800 350.400 ;
        RECT 209.200 350.300 210.000 350.400 ;
        RECT 220.400 350.300 221.200 350.400 ;
        RECT 206.000 349.700 221.200 350.300 ;
        RECT 206.000 349.600 206.800 349.700 ;
        RECT 209.200 349.600 210.000 349.700 ;
        RECT 220.400 349.600 221.200 349.700 ;
        RECT 242.800 350.300 243.600 350.400 ;
        RECT 268.400 350.300 269.200 350.400 ;
        RECT 242.800 349.700 269.200 350.300 ;
        RECT 242.800 349.600 243.600 349.700 ;
        RECT 268.400 349.600 269.200 349.700 ;
        RECT 297.200 350.300 298.000 350.400 ;
        RECT 306.800 350.300 307.600 350.400 ;
        RECT 297.200 349.700 307.600 350.300 ;
        RECT 297.200 349.600 298.000 349.700 ;
        RECT 306.800 349.600 307.600 349.700 ;
        RECT 310.000 350.300 310.800 350.400 ;
        RECT 314.800 350.300 315.600 350.400 ;
        RECT 321.200 350.300 322.000 350.400 ;
        RECT 310.000 349.700 322.000 350.300 ;
        RECT 310.000 349.600 310.800 349.700 ;
        RECT 314.800 349.600 315.600 349.700 ;
        RECT 321.200 349.600 322.000 349.700 ;
        RECT 337.200 350.300 338.000 350.400 ;
        RECT 342.000 350.300 342.800 350.400 ;
        RECT 337.200 349.700 342.800 350.300 ;
        RECT 337.200 349.600 338.000 349.700 ;
        RECT 342.000 349.600 342.800 349.700 ;
        RECT 346.800 350.300 347.600 350.400 ;
        RECT 353.200 350.300 354.000 350.400 ;
        RECT 346.800 349.700 354.000 350.300 ;
        RECT 346.800 349.600 347.600 349.700 ;
        RECT 353.200 349.600 354.000 349.700 ;
        RECT 372.400 349.600 373.200 350.400 ;
        RECT 374.000 350.300 374.800 350.400 ;
        RECT 404.400 350.300 405.200 350.400 ;
        RECT 374.000 349.700 405.200 350.300 ;
        RECT 374.000 349.600 374.800 349.700 ;
        RECT 404.400 349.600 405.200 349.700 ;
        RECT 406.000 350.300 406.800 350.400 ;
        RECT 410.800 350.300 411.600 350.400 ;
        RECT 406.000 349.700 411.600 350.300 ;
        RECT 406.000 349.600 406.800 349.700 ;
        RECT 410.800 349.600 411.600 349.700 ;
        RECT 412.400 350.300 413.200 350.400 ;
        RECT 422.000 350.300 422.800 350.400 ;
        RECT 412.400 349.700 422.800 350.300 ;
        RECT 412.400 349.600 413.200 349.700 ;
        RECT 422.000 349.600 422.800 349.700 ;
        RECT 436.400 350.300 437.200 350.400 ;
        RECT 442.800 350.300 443.600 350.400 ;
        RECT 436.400 349.700 443.600 350.300 ;
        RECT 436.400 349.600 437.200 349.700 ;
        RECT 442.800 349.600 443.600 349.700 ;
        RECT 449.200 349.600 450.000 350.400 ;
        RECT 458.800 350.300 459.600 350.400 ;
        RECT 462.000 350.300 462.800 350.400 ;
        RECT 458.800 349.700 462.800 350.300 ;
        RECT 458.800 349.600 459.600 349.700 ;
        RECT 462.000 349.600 462.800 349.700 ;
        RECT 465.200 350.300 466.000 350.400 ;
        RECT 478.000 350.300 478.800 350.400 ;
        RECT 465.200 349.700 478.800 350.300 ;
        RECT 465.200 349.600 466.000 349.700 ;
        RECT 478.000 349.600 478.800 349.700 ;
        RECT 479.600 350.300 480.400 350.400 ;
        RECT 484.400 350.300 485.200 350.400 ;
        RECT 479.600 349.700 485.200 350.300 ;
        RECT 479.600 349.600 480.400 349.700 ;
        RECT 484.400 349.600 485.200 349.700 ;
        RECT 492.400 350.300 493.200 350.400 ;
        RECT 497.200 350.300 498.000 350.400 ;
        RECT 492.400 349.700 498.000 350.300 ;
        RECT 492.400 349.600 493.200 349.700 ;
        RECT 497.200 349.600 498.000 349.700 ;
        RECT 498.800 350.300 499.600 350.400 ;
        RECT 513.200 350.300 514.000 350.400 ;
        RECT 498.800 349.700 514.000 350.300 ;
        RECT 498.800 349.600 499.600 349.700 ;
        RECT 513.200 349.600 514.000 349.700 ;
        RECT 22.000 348.300 22.800 348.400 ;
        RECT 44.400 348.300 45.200 348.400 ;
        RECT 22.000 347.700 45.200 348.300 ;
        RECT 22.000 347.600 22.800 347.700 ;
        RECT 44.400 347.600 45.200 347.700 ;
        RECT 111.600 348.300 112.400 348.400 ;
        RECT 170.800 348.300 171.600 348.400 ;
        RECT 111.600 347.700 171.600 348.300 ;
        RECT 111.600 347.600 112.400 347.700 ;
        RECT 170.800 347.600 171.600 347.700 ;
        RECT 257.200 348.300 258.000 348.400 ;
        RECT 322.800 348.300 323.600 348.400 ;
        RECT 338.800 348.300 339.600 348.400 ;
        RECT 345.200 348.300 346.000 348.400 ;
        RECT 257.200 347.700 323.600 348.300 ;
        RECT 257.200 347.600 258.000 347.700 ;
        RECT 322.800 347.600 323.600 347.700 ;
        RECT 324.500 347.700 346.000 348.300 ;
        RECT 193.200 346.300 194.000 346.400 ;
        RECT 228.400 346.300 229.200 346.400 ;
        RECT 193.200 345.700 229.200 346.300 ;
        RECT 193.200 345.600 194.000 345.700 ;
        RECT 228.400 345.600 229.200 345.700 ;
        RECT 278.000 346.300 278.800 346.400 ;
        RECT 286.000 346.300 286.800 346.400 ;
        RECT 278.000 345.700 286.800 346.300 ;
        RECT 278.000 345.600 278.800 345.700 ;
        RECT 286.000 345.600 286.800 345.700 ;
        RECT 318.000 346.300 318.800 346.400 ;
        RECT 324.500 346.300 325.100 347.700 ;
        RECT 338.800 347.600 339.600 347.700 ;
        RECT 345.200 347.600 346.000 347.700 ;
        RECT 351.600 348.300 352.400 348.400 ;
        RECT 410.800 348.300 411.600 348.400 ;
        RECT 452.400 348.300 453.200 348.400 ;
        RECT 466.800 348.300 467.600 348.400 ;
        RECT 471.600 348.300 472.400 348.400 ;
        RECT 487.600 348.300 488.400 348.400 ;
        RECT 351.600 347.700 488.400 348.300 ;
        RECT 351.600 347.600 352.400 347.700 ;
        RECT 410.800 347.600 411.600 347.700 ;
        RECT 452.400 347.600 453.200 347.700 ;
        RECT 466.800 347.600 467.600 347.700 ;
        RECT 471.600 347.600 472.400 347.700 ;
        RECT 487.600 347.600 488.400 347.700 ;
        RECT 318.000 345.700 325.100 346.300 ;
        RECT 334.000 346.300 334.800 346.400 ;
        RECT 340.400 346.300 341.200 346.400 ;
        RECT 364.400 346.300 365.200 346.400 ;
        RECT 385.200 346.300 386.000 346.400 ;
        RECT 420.400 346.300 421.200 346.400 ;
        RECT 334.000 345.700 421.200 346.300 ;
        RECT 318.000 345.600 318.800 345.700 ;
        RECT 334.000 345.600 334.800 345.700 ;
        RECT 340.400 345.600 341.200 345.700 ;
        RECT 364.400 345.600 365.200 345.700 ;
        RECT 385.200 345.600 386.000 345.700 ;
        RECT 409.300 344.400 409.900 345.700 ;
        RECT 420.400 345.600 421.200 345.700 ;
        RECT 442.800 346.300 443.600 346.400 ;
        RECT 454.000 346.300 454.800 346.400 ;
        RECT 442.800 345.700 454.800 346.300 ;
        RECT 442.800 345.600 443.600 345.700 ;
        RECT 454.000 345.600 454.800 345.700 ;
        RECT 465.200 346.300 466.000 346.400 ;
        RECT 468.400 346.300 469.200 346.400 ;
        RECT 465.200 345.700 469.200 346.300 ;
        RECT 465.200 345.600 466.000 345.700 ;
        RECT 468.400 345.600 469.200 345.700 ;
        RECT 473.200 346.300 474.000 346.400 ;
        RECT 479.600 346.300 480.400 346.400 ;
        RECT 473.200 345.700 480.400 346.300 ;
        RECT 473.200 345.600 474.000 345.700 ;
        RECT 479.600 345.600 480.400 345.700 ;
        RECT 2.800 344.300 3.600 344.400 ;
        RECT 39.600 344.300 40.400 344.400 ;
        RECT 2.800 343.700 40.400 344.300 ;
        RECT 2.800 343.600 3.600 343.700 ;
        RECT 39.600 343.600 40.400 343.700 ;
        RECT 74.800 344.300 75.600 344.400 ;
        RECT 89.200 344.300 90.000 344.400 ;
        RECT 74.800 343.700 90.000 344.300 ;
        RECT 74.800 343.600 75.600 343.700 ;
        RECT 89.200 343.600 90.000 343.700 ;
        RECT 231.600 344.300 232.400 344.400 ;
        RECT 238.000 344.300 238.800 344.400 ;
        RECT 231.600 343.700 238.800 344.300 ;
        RECT 231.600 343.600 232.400 343.700 ;
        RECT 238.000 343.600 238.800 343.700 ;
        RECT 265.200 344.300 266.000 344.400 ;
        RECT 281.200 344.300 282.000 344.400 ;
        RECT 290.800 344.300 291.600 344.400 ;
        RECT 265.200 343.700 291.600 344.300 ;
        RECT 265.200 343.600 266.000 343.700 ;
        RECT 281.200 343.600 282.000 343.700 ;
        RECT 290.800 343.600 291.600 343.700 ;
        RECT 306.800 344.300 307.600 344.400 ;
        RECT 326.000 344.300 326.800 344.400 ;
        RECT 306.800 343.700 326.800 344.300 ;
        RECT 306.800 343.600 307.600 343.700 ;
        RECT 326.000 343.600 326.800 343.700 ;
        RECT 329.200 344.300 330.000 344.400 ;
        RECT 351.600 344.300 352.400 344.400 ;
        RECT 366.000 344.300 366.800 344.400 ;
        RECT 329.200 343.700 366.800 344.300 ;
        RECT 329.200 343.600 330.000 343.700 ;
        RECT 351.600 343.600 352.400 343.700 ;
        RECT 366.000 343.600 366.800 343.700 ;
        RECT 367.600 344.300 368.400 344.400 ;
        RECT 370.800 344.300 371.600 344.400 ;
        RECT 394.800 344.300 395.600 344.400 ;
        RECT 367.600 343.700 395.600 344.300 ;
        RECT 367.600 343.600 368.400 343.700 ;
        RECT 370.800 343.600 371.600 343.700 ;
        RECT 394.800 343.600 395.600 343.700 ;
        RECT 396.400 344.300 397.200 344.400 ;
        RECT 401.200 344.300 402.000 344.400 ;
        RECT 396.400 343.700 402.000 344.300 ;
        RECT 396.400 343.600 397.200 343.700 ;
        RECT 401.200 343.600 402.000 343.700 ;
        RECT 409.200 343.600 410.000 344.400 ;
        RECT 410.800 343.600 411.600 344.400 ;
        RECT 460.400 344.300 461.200 344.400 ;
        RECT 486.000 344.300 486.800 344.400 ;
        RECT 460.400 343.700 486.800 344.300 ;
        RECT 460.400 343.600 461.200 343.700 ;
        RECT 486.000 343.600 486.800 343.700 ;
        RECT 487.600 344.300 488.400 344.400 ;
        RECT 502.000 344.300 502.800 344.400 ;
        RECT 487.600 343.700 502.800 344.300 ;
        RECT 487.600 343.600 488.400 343.700 ;
        RECT 502.000 343.600 502.800 343.700 ;
        RECT 506.800 344.300 507.600 344.400 ;
        RECT 522.800 344.300 523.600 344.400 ;
        RECT 506.800 343.700 523.600 344.300 ;
        RECT 506.800 343.600 507.600 343.700 ;
        RECT 522.800 343.600 523.600 343.700 ;
        RECT 538.800 344.300 539.600 344.400 ;
        RECT 548.400 344.300 549.200 344.400 ;
        RECT 538.800 343.700 549.200 344.300 ;
        RECT 538.800 343.600 539.600 343.700 ;
        RECT 548.400 343.600 549.200 343.700 ;
        RECT 50.800 342.300 51.600 342.400 ;
        RECT 68.400 342.300 69.200 342.400 ;
        RECT 50.800 341.700 69.200 342.300 ;
        RECT 50.800 341.600 51.600 341.700 ;
        RECT 68.400 341.600 69.200 341.700 ;
        RECT 111.600 342.300 112.400 342.400 ;
        RECT 114.800 342.300 115.600 342.400 ;
        RECT 129.200 342.300 130.000 342.400 ;
        RECT 151.600 342.300 152.400 342.400 ;
        RECT 156.400 342.300 157.200 342.400 ;
        RECT 164.400 342.300 165.200 342.400 ;
        RECT 193.200 342.300 194.000 342.400 ;
        RECT 111.600 341.700 194.000 342.300 ;
        RECT 111.600 341.600 112.400 341.700 ;
        RECT 114.800 341.600 115.600 341.700 ;
        RECT 129.200 341.600 130.000 341.700 ;
        RECT 151.600 341.600 152.400 341.700 ;
        RECT 156.400 341.600 157.200 341.700 ;
        RECT 164.400 341.600 165.200 341.700 ;
        RECT 193.200 341.600 194.000 341.700 ;
        RECT 196.400 342.300 197.200 342.400 ;
        RECT 199.600 342.300 200.400 342.400 ;
        RECT 196.400 341.700 200.400 342.300 ;
        RECT 196.400 341.600 197.200 341.700 ;
        RECT 199.600 341.600 200.400 341.700 ;
        RECT 345.200 342.300 346.000 342.400 ;
        RECT 364.400 342.300 365.200 342.400 ;
        RECT 345.200 341.700 365.200 342.300 ;
        RECT 366.100 342.300 366.700 343.600 ;
        RECT 455.600 342.300 456.400 342.400 ;
        RECT 366.100 341.700 456.400 342.300 ;
        RECT 345.200 341.600 346.000 341.700 ;
        RECT 364.400 341.600 365.200 341.700 ;
        RECT 455.600 341.600 456.400 341.700 ;
        RECT 457.200 342.300 458.000 342.400 ;
        RECT 473.200 342.300 474.000 342.400 ;
        RECT 457.200 341.700 474.000 342.300 ;
        RECT 457.200 341.600 458.000 341.700 ;
        RECT 473.200 341.600 474.000 341.700 ;
        RECT 516.400 342.300 517.200 342.400 ;
        RECT 524.400 342.300 525.200 342.400 ;
        RECT 516.400 341.700 525.200 342.300 ;
        RECT 516.400 341.600 517.200 341.700 ;
        RECT 524.400 341.600 525.200 341.700 ;
        RECT 18.800 340.300 19.600 340.400 ;
        RECT 22.000 340.300 22.800 340.400 ;
        RECT 18.800 339.700 22.800 340.300 ;
        RECT 18.800 339.600 19.600 339.700 ;
        RECT 22.000 339.600 22.800 339.700 ;
        RECT 52.400 340.300 53.200 340.400 ;
        RECT 81.200 340.300 82.000 340.400 ;
        RECT 52.400 339.700 82.000 340.300 ;
        RECT 52.400 339.600 53.200 339.700 ;
        RECT 81.200 339.600 82.000 339.700 ;
        RECT 153.200 339.600 154.000 340.400 ;
        RECT 177.200 340.300 178.000 340.400 ;
        RECT 191.600 340.300 192.400 340.400 ;
        RECT 177.200 339.700 192.400 340.300 ;
        RECT 177.200 339.600 178.000 339.700 ;
        RECT 191.600 339.600 192.400 339.700 ;
        RECT 327.600 340.300 328.400 340.400 ;
        RECT 337.200 340.300 338.000 340.400 ;
        RECT 327.600 339.700 338.000 340.300 ;
        RECT 327.600 339.600 328.400 339.700 ;
        RECT 337.200 339.600 338.000 339.700 ;
        RECT 342.000 340.300 342.800 340.400 ;
        RECT 354.800 340.300 355.600 340.400 ;
        RECT 342.000 339.700 355.600 340.300 ;
        RECT 342.000 339.600 342.800 339.700 ;
        RECT 354.800 339.600 355.600 339.700 ;
        RECT 356.400 340.300 357.200 340.400 ;
        RECT 366.000 340.300 366.800 340.400 ;
        RECT 447.600 340.300 448.400 340.400 ;
        RECT 356.400 339.700 448.400 340.300 ;
        RECT 356.400 339.600 357.200 339.700 ;
        RECT 366.000 339.600 366.800 339.700 ;
        RECT 447.600 339.600 448.400 339.700 ;
        RECT 468.400 340.300 469.200 340.400 ;
        RECT 470.000 340.300 470.800 340.400 ;
        RECT 468.400 339.700 470.800 340.300 ;
        RECT 468.400 339.600 469.200 339.700 ;
        RECT 470.000 339.600 470.800 339.700 ;
        RECT 57.200 338.300 58.000 338.400 ;
        RECT 73.200 338.300 74.000 338.400 ;
        RECT 95.600 338.300 96.400 338.400 ;
        RECT 57.200 337.700 96.400 338.300 ;
        RECT 153.300 338.300 153.900 339.600 ;
        RECT 194.800 338.300 195.600 338.400 ;
        RECT 153.300 337.700 195.600 338.300 ;
        RECT 57.200 337.600 58.000 337.700 ;
        RECT 73.200 337.600 74.000 337.700 ;
        RECT 95.600 337.600 96.400 337.700 ;
        RECT 194.800 337.600 195.600 337.700 ;
        RECT 290.800 338.300 291.600 338.400 ;
        RECT 308.400 338.300 309.200 338.400 ;
        RECT 324.400 338.300 325.200 338.400 ;
        RECT 326.000 338.300 326.800 338.400 ;
        RECT 290.800 337.700 326.800 338.300 ;
        RECT 290.800 337.600 291.600 337.700 ;
        RECT 308.400 337.600 309.200 337.700 ;
        RECT 324.400 337.600 325.200 337.700 ;
        RECT 326.000 337.600 326.800 337.700 ;
        RECT 362.800 338.300 363.600 338.400 ;
        RECT 382.000 338.300 382.800 338.400 ;
        RECT 362.800 337.700 382.800 338.300 ;
        RECT 362.800 337.600 363.600 337.700 ;
        RECT 382.000 337.600 382.800 337.700 ;
        RECT 399.600 338.300 400.400 338.400 ;
        RECT 412.400 338.300 413.200 338.400 ;
        RECT 436.400 338.300 437.200 338.400 ;
        RECT 399.600 337.700 437.200 338.300 ;
        RECT 399.600 337.600 400.400 337.700 ;
        RECT 412.400 337.600 413.200 337.700 ;
        RECT 436.400 337.600 437.200 337.700 ;
        RECT 458.800 338.300 459.600 338.400 ;
        RECT 503.600 338.300 504.400 338.400 ;
        RECT 458.800 337.700 504.400 338.300 ;
        RECT 458.800 337.600 459.600 337.700 ;
        RECT 503.600 337.600 504.400 337.700 ;
        RECT 506.800 338.300 507.600 338.400 ;
        RECT 514.800 338.300 515.600 338.400 ;
        RECT 506.800 337.700 515.600 338.300 ;
        RECT 506.800 337.600 507.600 337.700 ;
        RECT 514.800 337.600 515.600 337.700 ;
        RECT 522.800 338.300 523.600 338.400 ;
        RECT 537.200 338.300 538.000 338.400 ;
        RECT 522.800 337.700 538.000 338.300 ;
        RECT 522.800 337.600 523.600 337.700 ;
        RECT 537.200 337.600 538.000 337.700 ;
        RECT 49.200 336.300 50.000 336.400 ;
        RECT 74.800 336.300 75.600 336.400 ;
        RECT 49.200 335.700 75.600 336.300 ;
        RECT 49.200 335.600 50.000 335.700 ;
        RECT 74.800 335.600 75.600 335.700 ;
        RECT 228.400 336.300 229.200 336.400 ;
        RECT 236.400 336.300 237.200 336.400 ;
        RECT 228.400 335.700 237.200 336.300 ;
        RECT 228.400 335.600 229.200 335.700 ;
        RECT 236.400 335.600 237.200 335.700 ;
        RECT 247.600 336.300 248.400 336.400 ;
        RECT 356.400 336.300 357.200 336.400 ;
        RECT 247.600 335.700 357.200 336.300 ;
        RECT 247.600 335.600 248.400 335.700 ;
        RECT 356.400 335.600 357.200 335.700 ;
        RECT 364.400 336.300 365.200 336.400 ;
        RECT 374.000 336.300 374.800 336.400 ;
        RECT 364.400 335.700 374.800 336.300 ;
        RECT 364.400 335.600 365.200 335.700 ;
        RECT 374.000 335.600 374.800 335.700 ;
        RECT 375.600 336.300 376.400 336.400 ;
        RECT 391.600 336.300 392.400 336.400 ;
        RECT 375.600 335.700 392.400 336.300 ;
        RECT 375.600 335.600 376.400 335.700 ;
        RECT 391.600 335.600 392.400 335.700 ;
        RECT 398.000 336.300 398.800 336.400 ;
        RECT 417.200 336.300 418.000 336.400 ;
        RECT 398.000 335.700 418.000 336.300 ;
        RECT 398.000 335.600 398.800 335.700 ;
        RECT 417.200 335.600 418.000 335.700 ;
        RECT 422.000 336.300 422.800 336.400 ;
        RECT 444.400 336.300 445.200 336.400 ;
        RECT 465.200 336.300 466.000 336.400 ;
        RECT 474.800 336.300 475.600 336.400 ;
        RECT 422.000 335.700 475.600 336.300 ;
        RECT 422.000 335.600 422.800 335.700 ;
        RECT 444.400 335.600 445.200 335.700 ;
        RECT 465.200 335.600 466.000 335.700 ;
        RECT 474.800 335.600 475.600 335.700 ;
        RECT 503.600 336.300 504.400 336.400 ;
        RECT 516.400 336.300 517.200 336.400 ;
        RECT 503.600 335.700 517.200 336.300 ;
        RECT 503.600 335.600 504.400 335.700 ;
        RECT 516.400 335.600 517.200 335.700 ;
        RECT 521.200 336.300 522.000 336.400 ;
        RECT 543.600 336.300 544.400 336.400 ;
        RECT 521.200 335.700 544.400 336.300 ;
        RECT 521.200 335.600 522.000 335.700 ;
        RECT 543.600 335.600 544.400 335.700 ;
        RECT 46.000 334.300 46.800 334.400 ;
        RECT 52.400 334.300 53.200 334.400 ;
        RECT 46.000 333.700 53.200 334.300 ;
        RECT 46.000 333.600 46.800 333.700 ;
        RECT 52.400 333.600 53.200 333.700 ;
        RECT 79.600 334.300 80.400 334.400 ;
        RECT 89.200 334.300 90.000 334.400 ;
        RECT 97.200 334.300 98.000 334.400 ;
        RECT 79.600 333.700 98.000 334.300 ;
        RECT 79.600 333.600 80.400 333.700 ;
        RECT 89.200 333.600 90.000 333.700 ;
        RECT 97.200 333.600 98.000 333.700 ;
        RECT 159.600 334.300 160.400 334.400 ;
        RECT 169.200 334.300 170.000 334.400 ;
        RECT 159.600 333.700 170.000 334.300 ;
        RECT 159.600 333.600 160.400 333.700 ;
        RECT 169.200 333.600 170.000 333.700 ;
        RECT 186.800 334.300 187.600 334.400 ;
        RECT 193.200 334.300 194.000 334.400 ;
        RECT 201.200 334.300 202.000 334.400 ;
        RECT 186.800 333.700 202.000 334.300 ;
        RECT 186.800 333.600 187.600 333.700 ;
        RECT 193.200 333.600 194.000 333.700 ;
        RECT 201.200 333.600 202.000 333.700 ;
        RECT 239.600 334.300 240.400 334.400 ;
        RECT 255.600 334.300 256.400 334.400 ;
        RECT 239.600 333.700 256.400 334.300 ;
        RECT 239.600 333.600 240.400 333.700 ;
        RECT 255.600 333.600 256.400 333.700 ;
        RECT 353.200 334.300 354.000 334.400 ;
        RECT 401.200 334.300 402.000 334.400 ;
        RECT 422.100 334.300 422.700 335.600 ;
        RECT 353.200 333.700 422.700 334.300 ;
        RECT 436.400 334.300 437.200 334.400 ;
        RECT 471.600 334.300 472.400 334.400 ;
        RECT 436.400 333.700 472.400 334.300 ;
        RECT 353.200 333.600 354.000 333.700 ;
        RECT 401.200 333.600 402.000 333.700 ;
        RECT 436.400 333.600 437.200 333.700 ;
        RECT 471.600 333.600 472.400 333.700 ;
        RECT 508.400 334.300 509.200 334.400 ;
        RECT 516.400 334.300 517.200 334.400 ;
        RECT 535.600 334.300 536.400 334.400 ;
        RECT 508.400 333.700 536.400 334.300 ;
        RECT 508.400 333.600 509.200 333.700 ;
        RECT 516.400 333.600 517.200 333.700 ;
        RECT 535.600 333.600 536.400 333.700 ;
        RECT 41.200 332.300 42.000 332.400 ;
        RECT 57.200 332.300 58.000 332.400 ;
        RECT 41.200 331.700 58.000 332.300 ;
        RECT 41.200 331.600 42.000 331.700 ;
        RECT 57.200 331.600 58.000 331.700 ;
        RECT 63.600 332.300 64.400 332.400 ;
        RECT 66.800 332.300 67.600 332.400 ;
        RECT 63.600 331.700 67.600 332.300 ;
        RECT 63.600 331.600 64.400 331.700 ;
        RECT 66.800 331.600 67.600 331.700 ;
        RECT 82.800 332.300 83.600 332.400 ;
        RECT 87.600 332.300 88.400 332.400 ;
        RECT 90.800 332.300 91.600 332.400 ;
        RECT 82.800 331.700 91.600 332.300 ;
        RECT 82.800 331.600 83.600 331.700 ;
        RECT 87.600 331.600 88.400 331.700 ;
        RECT 90.800 331.600 91.600 331.700 ;
        RECT 220.400 332.300 221.200 332.400 ;
        RECT 228.400 332.300 229.200 332.400 ;
        RECT 220.400 331.700 229.200 332.300 ;
        RECT 220.400 331.600 221.200 331.700 ;
        RECT 228.400 331.600 229.200 331.700 ;
        RECT 310.000 332.300 310.800 332.400 ;
        RECT 337.200 332.300 338.000 332.400 ;
        RECT 343.600 332.300 344.400 332.400 ;
        RECT 310.000 331.700 344.400 332.300 ;
        RECT 310.000 331.600 310.800 331.700 ;
        RECT 337.200 331.600 338.000 331.700 ;
        RECT 343.600 331.600 344.400 331.700 ;
        RECT 354.800 332.300 355.600 332.400 ;
        RECT 362.800 332.300 363.600 332.400 ;
        RECT 375.600 332.300 376.400 332.400 ;
        RECT 354.800 331.700 376.400 332.300 ;
        RECT 354.800 331.600 355.600 331.700 ;
        RECT 362.800 331.600 363.600 331.700 ;
        RECT 375.600 331.600 376.400 331.700 ;
        RECT 382.000 332.300 382.800 332.400 ;
        RECT 434.800 332.300 435.600 332.400 ;
        RECT 382.000 331.700 435.600 332.300 ;
        RECT 382.000 331.600 382.800 331.700 ;
        RECT 434.800 331.600 435.600 331.700 ;
        RECT 447.600 332.300 448.400 332.400 ;
        RECT 449.200 332.300 450.000 332.400 ;
        RECT 455.600 332.300 456.400 332.400 ;
        RECT 447.600 331.700 456.400 332.300 ;
        RECT 447.600 331.600 448.400 331.700 ;
        RECT 449.200 331.600 450.000 331.700 ;
        RECT 455.600 331.600 456.400 331.700 ;
        RECT 497.200 332.300 498.000 332.400 ;
        RECT 510.000 332.300 510.800 332.400 ;
        RECT 497.200 331.700 510.800 332.300 ;
        RECT 497.200 331.600 498.000 331.700 ;
        RECT 510.000 331.600 510.800 331.700 ;
        RECT 524.400 332.300 525.200 332.400 ;
        RECT 530.800 332.300 531.600 332.400 ;
        RECT 524.400 331.700 531.600 332.300 ;
        RECT 524.400 331.600 525.200 331.700 ;
        RECT 530.800 331.600 531.600 331.700 ;
        RECT 25.200 330.300 26.000 330.400 ;
        RECT 44.400 330.300 45.200 330.400 ;
        RECT 25.200 329.700 45.200 330.300 ;
        RECT 25.200 329.600 26.000 329.700 ;
        RECT 44.400 329.600 45.200 329.700 ;
        RECT 50.800 330.300 51.600 330.400 ;
        RECT 58.800 330.300 59.600 330.400 ;
        RECT 50.800 329.700 59.600 330.300 ;
        RECT 50.800 329.600 51.600 329.700 ;
        RECT 58.800 329.600 59.600 329.700 ;
        RECT 70.000 330.300 70.800 330.400 ;
        RECT 74.800 330.300 75.600 330.400 ;
        RECT 86.000 330.300 86.800 330.400 ;
        RECT 103.600 330.300 104.400 330.400 ;
        RECT 70.000 329.700 104.400 330.300 ;
        RECT 70.000 329.600 70.800 329.700 ;
        RECT 74.800 329.600 75.600 329.700 ;
        RECT 86.000 329.600 86.800 329.700 ;
        RECT 103.600 329.600 104.400 329.700 ;
        RECT 114.800 330.300 115.600 330.400 ;
        RECT 140.400 330.300 141.200 330.400 ;
        RECT 114.800 329.700 141.200 330.300 ;
        RECT 114.800 329.600 115.600 329.700 ;
        RECT 140.400 329.600 141.200 329.700 ;
        RECT 175.600 330.300 176.400 330.400 ;
        RECT 180.400 330.300 181.200 330.400 ;
        RECT 175.600 329.700 181.200 330.300 ;
        RECT 175.600 329.600 176.400 329.700 ;
        RECT 180.400 329.600 181.200 329.700 ;
        RECT 188.400 330.300 189.200 330.400 ;
        RECT 204.400 330.300 205.200 330.400 ;
        RECT 212.400 330.300 213.200 330.400 ;
        RECT 188.400 329.700 213.200 330.300 ;
        RECT 188.400 329.600 189.200 329.700 ;
        RECT 204.400 329.600 205.200 329.700 ;
        RECT 212.400 329.600 213.200 329.700 ;
        RECT 351.600 330.300 352.400 330.400 ;
        RECT 358.000 330.300 358.800 330.400 ;
        RECT 359.600 330.300 360.400 330.400 ;
        RECT 372.400 330.300 373.200 330.400 ;
        RECT 383.600 330.300 384.400 330.400 ;
        RECT 388.400 330.300 389.200 330.400 ;
        RECT 394.800 330.300 395.600 330.400 ;
        RECT 407.600 330.300 408.400 330.400 ;
        RECT 351.600 329.700 408.400 330.300 ;
        RECT 351.600 329.600 352.400 329.700 ;
        RECT 358.000 329.600 358.800 329.700 ;
        RECT 359.600 329.600 360.400 329.700 ;
        RECT 372.400 329.600 373.200 329.700 ;
        RECT 383.600 329.600 384.400 329.700 ;
        RECT 388.400 329.600 389.200 329.700 ;
        RECT 394.800 329.600 395.600 329.700 ;
        RECT 407.600 329.600 408.400 329.700 ;
        RECT 409.200 330.300 410.000 330.400 ;
        RECT 436.400 330.300 437.200 330.400 ;
        RECT 409.200 329.700 437.200 330.300 ;
        RECT 409.200 329.600 410.000 329.700 ;
        RECT 436.400 329.600 437.200 329.700 ;
        RECT 441.200 330.300 442.000 330.400 ;
        RECT 446.000 330.300 446.800 330.400 ;
        RECT 441.200 329.700 446.800 330.300 ;
        RECT 441.200 329.600 442.000 329.700 ;
        RECT 446.000 329.600 446.800 329.700 ;
        RECT 486.000 330.300 486.800 330.400 ;
        RECT 494.000 330.300 494.800 330.400 ;
        RECT 486.000 329.700 494.800 330.300 ;
        RECT 486.000 329.600 486.800 329.700 ;
        RECT 494.000 329.600 494.800 329.700 ;
        RECT 502.000 330.300 502.800 330.400 ;
        RECT 521.200 330.300 522.000 330.400 ;
        RECT 502.000 329.700 522.000 330.300 ;
        RECT 502.000 329.600 502.800 329.700 ;
        RECT 521.200 329.600 522.000 329.700 ;
        RECT 534.000 330.300 534.800 330.400 ;
        RECT 537.200 330.300 538.000 330.400 ;
        RECT 534.000 329.700 538.000 330.300 ;
        RECT 534.000 329.600 534.800 329.700 ;
        RECT 537.200 329.600 538.000 329.700 ;
        RECT 42.800 328.300 43.600 328.400 ;
        RECT 65.200 328.300 66.000 328.400 ;
        RECT 42.800 327.700 66.000 328.300 ;
        RECT 42.800 327.600 43.600 327.700 ;
        RECT 65.200 327.600 66.000 327.700 ;
        RECT 94.000 328.300 94.800 328.400 ;
        RECT 111.600 328.300 112.400 328.400 ;
        RECT 94.000 327.700 112.400 328.300 ;
        RECT 94.000 327.600 94.800 327.700 ;
        RECT 111.600 327.600 112.400 327.700 ;
        RECT 359.600 327.600 360.400 328.400 ;
        RECT 361.200 328.300 362.000 328.400 ;
        RECT 375.600 328.300 376.400 328.400 ;
        RECT 361.200 327.700 376.400 328.300 ;
        RECT 361.200 327.600 362.000 327.700 ;
        RECT 375.600 327.600 376.400 327.700 ;
        RECT 398.000 328.300 398.800 328.400 ;
        RECT 399.600 328.300 400.400 328.400 ;
        RECT 398.000 327.700 400.400 328.300 ;
        RECT 398.000 327.600 398.800 327.700 ;
        RECT 399.600 327.600 400.400 327.700 ;
        RECT 404.400 328.300 405.200 328.400 ;
        RECT 407.600 328.300 408.400 328.400 ;
        RECT 452.400 328.300 453.200 328.400 ;
        RECT 404.400 327.700 453.200 328.300 ;
        RECT 404.400 327.600 405.200 327.700 ;
        RECT 407.600 327.600 408.400 327.700 ;
        RECT 452.400 327.600 453.200 327.700 ;
        RECT 503.600 328.300 504.400 328.400 ;
        RECT 506.800 328.300 507.600 328.400 ;
        RECT 503.600 327.700 507.600 328.300 ;
        RECT 503.600 327.600 504.400 327.700 ;
        RECT 506.800 327.600 507.600 327.700 ;
        RECT 513.200 328.300 514.000 328.400 ;
        RECT 540.400 328.300 541.200 328.400 ;
        RECT 513.200 327.700 541.200 328.300 ;
        RECT 513.200 327.600 514.000 327.700 ;
        RECT 540.400 327.600 541.200 327.700 ;
        RECT 47.600 326.300 48.400 326.400 ;
        RECT 52.400 326.300 53.200 326.400 ;
        RECT 92.400 326.300 93.200 326.400 ;
        RECT 47.600 325.700 93.200 326.300 ;
        RECT 47.600 325.600 48.400 325.700 ;
        RECT 52.400 325.600 53.200 325.700 ;
        RECT 92.400 325.600 93.200 325.700 ;
        RECT 306.800 326.300 307.600 326.400 ;
        RECT 356.400 326.300 357.200 326.400 ;
        RECT 378.800 326.300 379.600 326.400 ;
        RECT 401.200 326.300 402.000 326.400 ;
        RECT 306.800 325.700 379.600 326.300 ;
        RECT 306.800 325.600 307.600 325.700 ;
        RECT 356.400 325.600 357.200 325.700 ;
        RECT 378.800 325.600 379.600 325.700 ;
        RECT 380.500 325.700 402.000 326.300 ;
        RECT 286.000 324.300 286.800 324.400 ;
        RECT 369.200 324.300 370.000 324.400 ;
        RECT 286.000 323.700 370.000 324.300 ;
        RECT 286.000 323.600 286.800 323.700 ;
        RECT 369.200 323.600 370.000 323.700 ;
        RECT 370.800 324.300 371.600 324.400 ;
        RECT 380.500 324.300 381.100 325.700 ;
        RECT 401.200 325.600 402.000 325.700 ;
        RECT 404.400 326.300 405.200 326.400 ;
        RECT 428.400 326.300 429.200 326.400 ;
        RECT 404.400 325.700 429.200 326.300 ;
        RECT 404.400 325.600 405.200 325.700 ;
        RECT 428.400 325.600 429.200 325.700 ;
        RECT 370.800 323.700 381.100 324.300 ;
        RECT 393.200 324.300 394.000 324.400 ;
        RECT 412.400 324.300 413.200 324.400 ;
        RECT 438.000 324.300 438.800 324.400 ;
        RECT 393.200 323.700 413.200 324.300 ;
        RECT 370.800 323.600 371.600 323.700 ;
        RECT 393.200 323.600 394.000 323.700 ;
        RECT 412.400 323.600 413.200 323.700 ;
        RECT 420.500 323.700 438.800 324.300 ;
        RECT 26.800 322.300 27.600 322.400 ;
        RECT 30.000 322.300 30.800 322.400 ;
        RECT 26.800 321.700 30.800 322.300 ;
        RECT 26.800 321.600 27.600 321.700 ;
        RECT 30.000 321.600 30.800 321.700 ;
        RECT 71.600 322.300 72.400 322.400 ;
        RECT 106.800 322.300 107.600 322.400 ;
        RECT 71.600 321.700 107.600 322.300 ;
        RECT 71.600 321.600 72.400 321.700 ;
        RECT 106.800 321.600 107.600 321.700 ;
        RECT 151.600 322.300 152.400 322.400 ;
        RECT 156.400 322.300 157.200 322.400 ;
        RECT 151.600 321.700 157.200 322.300 ;
        RECT 151.600 321.600 152.400 321.700 ;
        RECT 156.400 321.600 157.200 321.700 ;
        RECT 182.000 322.300 182.800 322.400 ;
        RECT 206.000 322.300 206.800 322.400 ;
        RECT 212.400 322.300 213.200 322.400 ;
        RECT 182.000 321.700 213.200 322.300 ;
        RECT 182.000 321.600 182.800 321.700 ;
        RECT 206.000 321.600 206.800 321.700 ;
        RECT 212.400 321.600 213.200 321.700 ;
        RECT 238.000 322.300 238.800 322.400 ;
        RECT 244.400 322.300 245.200 322.400 ;
        RECT 238.000 321.700 245.200 322.300 ;
        RECT 238.000 321.600 238.800 321.700 ;
        RECT 244.400 321.600 245.200 321.700 ;
        RECT 314.800 322.300 315.600 322.400 ;
        RECT 318.000 322.300 318.800 322.400 ;
        RECT 314.800 321.700 318.800 322.300 ;
        RECT 314.800 321.600 315.600 321.700 ;
        RECT 318.000 321.600 318.800 321.700 ;
        RECT 353.200 322.300 354.000 322.400 ;
        RECT 364.400 322.300 365.200 322.400 ;
        RECT 353.200 321.700 365.200 322.300 ;
        RECT 353.200 321.600 354.000 321.700 ;
        RECT 364.400 321.600 365.200 321.700 ;
        RECT 366.000 322.300 366.800 322.400 ;
        RECT 369.200 322.300 370.000 322.400 ;
        RECT 366.000 321.700 370.000 322.300 ;
        RECT 366.000 321.600 366.800 321.700 ;
        RECT 369.200 321.600 370.000 321.700 ;
        RECT 375.600 322.300 376.400 322.400 ;
        RECT 391.600 322.300 392.400 322.400 ;
        RECT 375.600 321.700 392.400 322.300 ;
        RECT 375.600 321.600 376.400 321.700 ;
        RECT 391.600 321.600 392.400 321.700 ;
        RECT 407.600 322.300 408.400 322.400 ;
        RECT 420.500 322.300 421.100 323.700 ;
        RECT 438.000 323.600 438.800 323.700 ;
        RECT 407.600 321.700 421.100 322.300 ;
        RECT 441.200 322.300 442.000 322.400 ;
        RECT 478.000 322.300 478.800 322.400 ;
        RECT 498.800 322.300 499.600 322.400 ;
        RECT 441.200 321.700 499.600 322.300 ;
        RECT 407.600 321.600 408.400 321.700 ;
        RECT 441.200 321.600 442.000 321.700 ;
        RECT 478.000 321.600 478.800 321.700 ;
        RECT 498.800 321.600 499.600 321.700 ;
        RECT 159.600 320.300 160.400 320.400 ;
        RECT 167.600 320.300 168.400 320.400 ;
        RECT 233.200 320.300 234.000 320.400 ;
        RECT 159.600 319.700 168.400 320.300 ;
        RECT 159.600 319.600 160.400 319.700 ;
        RECT 167.600 319.600 168.400 319.700 ;
        RECT 210.900 319.700 234.000 320.300 ;
        RECT 210.900 318.400 211.500 319.700 ;
        RECT 233.200 319.600 234.000 319.700 ;
        RECT 306.800 320.300 307.600 320.400 ;
        RECT 332.400 320.300 333.200 320.400 ;
        RECT 306.800 319.700 333.200 320.300 ;
        RECT 306.800 319.600 307.600 319.700 ;
        RECT 332.400 319.600 333.200 319.700 ;
        RECT 375.600 320.300 376.400 320.400 ;
        RECT 402.800 320.300 403.600 320.400 ;
        RECT 409.200 320.300 410.000 320.400 ;
        RECT 375.600 319.700 410.000 320.300 ;
        RECT 375.600 319.600 376.400 319.700 ;
        RECT 402.800 319.600 403.600 319.700 ;
        RECT 409.200 319.600 410.000 319.700 ;
        RECT 484.400 320.300 485.200 320.400 ;
        RECT 498.800 320.300 499.600 320.400 ;
        RECT 511.600 320.300 512.400 320.400 ;
        RECT 484.400 319.700 512.400 320.300 ;
        RECT 484.400 319.600 485.200 319.700 ;
        RECT 498.800 319.600 499.600 319.700 ;
        RECT 511.600 319.600 512.400 319.700 ;
        RECT 2.800 318.300 3.600 318.400 ;
        RECT 17.200 318.300 18.000 318.400 ;
        RECT 25.200 318.300 26.000 318.400 ;
        RECT 31.600 318.300 32.400 318.400 ;
        RECT 2.800 317.700 32.400 318.300 ;
        RECT 2.800 317.600 3.600 317.700 ;
        RECT 17.200 317.600 18.000 317.700 ;
        RECT 25.200 317.600 26.000 317.700 ;
        RECT 31.600 317.600 32.400 317.700 ;
        RECT 148.400 318.300 149.200 318.400 ;
        RECT 167.600 318.300 168.400 318.400 ;
        RECT 148.400 317.700 168.400 318.300 ;
        RECT 148.400 317.600 149.200 317.700 ;
        RECT 167.600 317.600 168.400 317.700 ;
        RECT 172.400 318.300 173.200 318.400 ;
        RECT 182.000 318.300 182.800 318.400 ;
        RECT 172.400 317.700 182.800 318.300 ;
        RECT 172.400 317.600 173.200 317.700 ;
        RECT 182.000 317.600 182.800 317.700 ;
        RECT 191.600 318.300 192.400 318.400 ;
        RECT 210.800 318.300 211.600 318.400 ;
        RECT 191.600 317.700 211.600 318.300 ;
        RECT 191.600 317.600 192.400 317.700 ;
        RECT 210.800 317.600 211.600 317.700 ;
        RECT 214.000 318.300 214.800 318.400 ;
        RECT 226.800 318.300 227.600 318.400 ;
        RECT 238.000 318.300 238.800 318.400 ;
        RECT 214.000 317.700 238.800 318.300 ;
        RECT 214.000 317.600 214.800 317.700 ;
        RECT 226.800 317.600 227.600 317.700 ;
        RECT 238.000 317.600 238.800 317.700 ;
        RECT 287.600 318.300 288.400 318.400 ;
        RECT 330.800 318.300 331.600 318.400 ;
        RECT 287.600 317.700 331.600 318.300 ;
        RECT 287.600 317.600 288.400 317.700 ;
        RECT 330.800 317.600 331.600 317.700 ;
        RECT 346.800 318.300 347.600 318.400 ;
        RECT 442.800 318.300 443.600 318.400 ;
        RECT 346.800 317.700 443.600 318.300 ;
        RECT 346.800 317.600 347.600 317.700 ;
        RECT 442.800 317.600 443.600 317.700 ;
        RECT 473.200 318.300 474.000 318.400 ;
        RECT 474.800 318.300 475.600 318.400 ;
        RECT 473.200 317.700 475.600 318.300 ;
        RECT 473.200 317.600 474.000 317.700 ;
        RECT 474.800 317.600 475.600 317.700 ;
        RECT 47.600 316.300 48.400 316.400 ;
        RECT 52.400 316.300 53.200 316.400 ;
        RECT 47.600 315.700 53.200 316.300 ;
        RECT 47.600 315.600 48.400 315.700 ;
        RECT 52.400 315.600 53.200 315.700 ;
        RECT 54.000 316.300 54.800 316.400 ;
        RECT 55.600 316.300 56.400 316.400 ;
        RECT 60.400 316.300 61.200 316.400 ;
        RECT 54.000 315.700 61.200 316.300 ;
        RECT 54.000 315.600 54.800 315.700 ;
        RECT 55.600 315.600 56.400 315.700 ;
        RECT 60.400 315.600 61.200 315.700 ;
        RECT 199.600 316.300 200.400 316.400 ;
        RECT 230.000 316.300 230.800 316.400 ;
        RECT 199.600 315.700 230.800 316.300 ;
        RECT 199.600 315.600 200.400 315.700 ;
        RECT 230.000 315.600 230.800 315.700 ;
        RECT 236.400 316.300 237.200 316.400 ;
        RECT 266.800 316.300 267.600 316.400 ;
        RECT 434.800 316.300 435.600 316.400 ;
        RECT 236.400 315.700 267.600 316.300 ;
        RECT 236.400 315.600 237.200 315.700 ;
        RECT 266.800 315.600 267.600 315.700 ;
        RECT 370.900 315.700 435.600 316.300 ;
        RECT 370.900 314.400 371.500 315.700 ;
        RECT 434.800 315.600 435.600 315.700 ;
        RECT 9.200 314.300 10.000 314.400 ;
        RECT 12.400 314.300 13.200 314.400 ;
        RECT 9.200 313.700 13.200 314.300 ;
        RECT 9.200 313.600 10.000 313.700 ;
        RECT 12.400 313.600 13.200 313.700 ;
        RECT 23.600 314.300 24.400 314.400 ;
        RECT 38.000 314.300 38.800 314.400 ;
        RECT 23.600 313.700 38.800 314.300 ;
        RECT 23.600 313.600 24.400 313.700 ;
        RECT 38.000 313.600 38.800 313.700 ;
        RECT 41.200 314.300 42.000 314.400 ;
        RECT 57.200 314.300 58.000 314.400 ;
        RECT 41.200 313.700 58.000 314.300 ;
        RECT 41.200 313.600 42.000 313.700 ;
        RECT 57.200 313.600 58.000 313.700 ;
        RECT 73.200 314.300 74.000 314.400 ;
        RECT 105.200 314.300 106.000 314.400 ;
        RECT 73.200 313.700 106.000 314.300 ;
        RECT 73.200 313.600 74.000 313.700 ;
        RECT 105.200 313.600 106.000 313.700 ;
        RECT 140.400 314.300 141.200 314.400 ;
        RECT 175.600 314.300 176.400 314.400 ;
        RECT 140.400 313.700 176.400 314.300 ;
        RECT 140.400 313.600 141.200 313.700 ;
        RECT 175.600 313.600 176.400 313.700 ;
        RECT 209.200 314.300 210.000 314.400 ;
        RECT 218.800 314.300 219.600 314.400 ;
        RECT 209.200 313.700 219.600 314.300 ;
        RECT 209.200 313.600 210.000 313.700 ;
        RECT 218.800 313.600 219.600 313.700 ;
        RECT 326.000 314.300 326.800 314.400 ;
        RECT 335.600 314.300 336.400 314.400 ;
        RECT 326.000 313.700 336.400 314.300 ;
        RECT 326.000 313.600 326.800 313.700 ;
        RECT 335.600 313.600 336.400 313.700 ;
        RECT 337.200 314.300 338.000 314.400 ;
        RECT 348.400 314.300 349.200 314.400 ;
        RECT 370.800 314.300 371.600 314.400 ;
        RECT 337.200 313.700 371.600 314.300 ;
        RECT 337.200 313.600 338.000 313.700 ;
        RECT 348.400 313.600 349.200 313.700 ;
        RECT 370.800 313.600 371.600 313.700 ;
        RECT 375.600 313.600 376.400 314.400 ;
        RECT 386.800 314.300 387.600 314.400 ;
        RECT 398.000 314.300 398.800 314.400 ;
        RECT 401.200 314.300 402.000 314.400 ;
        RECT 406.000 314.300 406.800 314.400 ;
        RECT 386.800 313.700 406.800 314.300 ;
        RECT 386.800 313.600 387.600 313.700 ;
        RECT 398.000 313.600 398.800 313.700 ;
        RECT 401.200 313.600 402.000 313.700 ;
        RECT 406.000 313.600 406.800 313.700 ;
        RECT 1.200 312.300 2.000 312.400 ;
        RECT 6.000 312.300 6.800 312.400 ;
        RECT 1.200 311.700 6.800 312.300 ;
        RECT 12.500 312.300 13.100 313.600 ;
        RECT 42.800 312.300 43.600 312.400 ;
        RECT 12.500 311.700 43.600 312.300 ;
        RECT 1.200 311.600 2.000 311.700 ;
        RECT 6.000 311.600 6.800 311.700 ;
        RECT 42.800 311.600 43.600 311.700 ;
        RECT 44.400 312.300 45.200 312.400 ;
        RECT 66.800 312.300 67.600 312.400 ;
        RECT 44.400 311.700 67.600 312.300 ;
        RECT 44.400 311.600 45.200 311.700 ;
        RECT 66.800 311.600 67.600 311.700 ;
        RECT 95.600 312.300 96.400 312.400 ;
        RECT 108.400 312.300 109.200 312.400 ;
        RECT 95.600 311.700 109.200 312.300 ;
        RECT 95.600 311.600 96.400 311.700 ;
        RECT 108.400 311.600 109.200 311.700 ;
        RECT 110.000 312.300 110.800 312.400 ;
        RECT 129.200 312.300 130.000 312.400 ;
        RECT 137.200 312.300 138.000 312.400 ;
        RECT 110.000 311.700 138.000 312.300 ;
        RECT 110.000 311.600 110.800 311.700 ;
        RECT 129.200 311.600 130.000 311.700 ;
        RECT 137.200 311.600 138.000 311.700 ;
        RECT 172.400 312.300 173.200 312.400 ;
        RECT 177.200 312.300 178.000 312.400 ;
        RECT 172.400 311.700 178.000 312.300 ;
        RECT 172.400 311.600 173.200 311.700 ;
        RECT 177.200 311.600 178.000 311.700 ;
        RECT 182.000 312.300 182.800 312.400 ;
        RECT 201.200 312.300 202.000 312.400 ;
        RECT 215.600 312.300 216.400 312.400 ;
        RECT 217.200 312.300 218.000 312.400 ;
        RECT 228.400 312.300 229.200 312.400 ;
        RECT 182.000 311.700 218.000 312.300 ;
        RECT 182.000 311.600 182.800 311.700 ;
        RECT 201.200 311.600 202.000 311.700 ;
        RECT 215.600 311.600 216.400 311.700 ;
        RECT 217.200 311.600 218.000 311.700 ;
        RECT 220.500 311.700 229.200 312.300 ;
        RECT 7.600 310.300 8.400 310.400 ;
        RECT 18.800 310.300 19.600 310.400 ;
        RECT 23.600 310.300 24.400 310.400 ;
        RECT 55.600 310.300 56.400 310.400 ;
        RECT 7.600 309.700 56.400 310.300 ;
        RECT 7.600 309.600 8.400 309.700 ;
        RECT 18.800 309.600 19.600 309.700 ;
        RECT 23.600 309.600 24.400 309.700 ;
        RECT 55.600 309.600 56.400 309.700 ;
        RECT 58.800 310.300 59.600 310.400 ;
        RECT 62.000 310.300 62.800 310.400 ;
        RECT 58.800 309.700 62.800 310.300 ;
        RECT 58.800 309.600 59.600 309.700 ;
        RECT 62.000 309.600 62.800 309.700 ;
        RECT 65.200 310.300 66.000 310.400 ;
        RECT 98.800 310.300 99.600 310.400 ;
        RECT 65.200 309.700 99.600 310.300 ;
        RECT 65.200 309.600 66.000 309.700 ;
        RECT 98.800 309.600 99.600 309.700 ;
        RECT 114.800 310.300 115.600 310.400 ;
        RECT 121.200 310.300 122.000 310.400 ;
        RECT 135.600 310.300 136.400 310.400 ;
        RECT 114.800 309.700 136.400 310.300 ;
        RECT 114.800 309.600 115.600 309.700 ;
        RECT 121.200 309.600 122.000 309.700 ;
        RECT 135.600 309.600 136.400 309.700 ;
        RECT 164.400 310.300 165.200 310.400 ;
        RECT 169.200 310.300 170.000 310.400 ;
        RECT 164.400 309.700 170.000 310.300 ;
        RECT 164.400 309.600 165.200 309.700 ;
        RECT 169.200 309.600 170.000 309.700 ;
        RECT 180.400 310.300 181.200 310.400 ;
        RECT 194.800 310.300 195.600 310.400 ;
        RECT 180.400 309.700 195.600 310.300 ;
        RECT 180.400 309.600 181.200 309.700 ;
        RECT 194.800 309.600 195.600 309.700 ;
        RECT 202.800 310.300 203.600 310.400 ;
        RECT 214.000 310.300 214.800 310.400 ;
        RECT 220.500 310.300 221.100 311.700 ;
        RECT 228.400 311.600 229.200 311.700 ;
        RECT 322.800 312.300 323.600 312.400 ;
        RECT 348.400 312.300 349.200 312.400 ;
        RECT 322.800 311.700 349.200 312.300 ;
        RECT 322.800 311.600 323.600 311.700 ;
        RECT 348.400 311.600 349.200 311.700 ;
        RECT 361.200 312.300 362.000 312.400 ;
        RECT 383.600 312.300 384.400 312.400 ;
        RECT 407.600 312.300 408.400 312.400 ;
        RECT 361.200 311.700 384.400 312.300 ;
        RECT 361.200 311.600 362.000 311.700 ;
        RECT 383.600 311.600 384.400 311.700 ;
        RECT 394.900 311.700 408.400 312.300 ;
        RECT 394.900 310.400 395.500 311.700 ;
        RECT 407.600 311.600 408.400 311.700 ;
        RECT 430.000 312.300 430.800 312.400 ;
        RECT 436.400 312.300 437.200 312.400 ;
        RECT 430.000 311.700 437.200 312.300 ;
        RECT 430.000 311.600 430.800 311.700 ;
        RECT 436.400 311.600 437.200 311.700 ;
        RECT 534.000 312.300 534.800 312.400 ;
        RECT 537.200 312.300 538.000 312.400 ;
        RECT 534.000 311.700 538.000 312.300 ;
        RECT 534.000 311.600 534.800 311.700 ;
        RECT 537.200 311.600 538.000 311.700 ;
        RECT 202.800 309.700 221.100 310.300 ;
        RECT 222.000 310.300 222.800 310.400 ;
        RECT 236.400 310.300 237.200 310.400 ;
        RECT 249.200 310.300 250.000 310.400 ;
        RECT 222.000 309.700 250.000 310.300 ;
        RECT 202.800 309.600 203.600 309.700 ;
        RECT 214.000 309.600 214.800 309.700 ;
        RECT 222.000 309.600 222.800 309.700 ;
        RECT 236.400 309.600 237.200 309.700 ;
        RECT 249.200 309.600 250.000 309.700 ;
        RECT 335.600 310.300 336.400 310.400 ;
        RECT 346.800 310.300 347.600 310.400 ;
        RECT 335.600 309.700 347.600 310.300 ;
        RECT 335.600 309.600 336.400 309.700 ;
        RECT 346.800 309.600 347.600 309.700 ;
        RECT 348.400 310.300 349.200 310.400 ;
        RECT 359.600 310.300 360.400 310.400 ;
        RECT 348.400 309.700 360.400 310.300 ;
        RECT 348.400 309.600 349.200 309.700 ;
        RECT 359.600 309.600 360.400 309.700 ;
        RECT 375.600 310.300 376.400 310.400 ;
        RECT 378.800 310.300 379.600 310.400 ;
        RECT 375.600 309.700 379.600 310.300 ;
        RECT 375.600 309.600 376.400 309.700 ;
        RECT 378.800 309.600 379.600 309.700 ;
        RECT 394.800 309.600 395.600 310.400 ;
        RECT 399.600 310.300 400.400 310.400 ;
        RECT 433.200 310.300 434.000 310.400 ;
        RECT 399.600 309.700 434.000 310.300 ;
        RECT 399.600 309.600 400.400 309.700 ;
        RECT 433.200 309.600 434.000 309.700 ;
        RECT 495.600 310.300 496.400 310.400 ;
        RECT 510.000 310.300 510.800 310.400 ;
        RECT 495.600 309.700 510.800 310.300 ;
        RECT 495.600 309.600 496.400 309.700 ;
        RECT 510.000 309.600 510.800 309.700 ;
        RECT 511.600 310.300 512.400 310.400 ;
        RECT 530.800 310.300 531.600 310.400 ;
        RECT 511.600 309.700 531.600 310.300 ;
        RECT 511.600 309.600 512.400 309.700 ;
        RECT 530.800 309.600 531.600 309.700 ;
        RECT 30.000 308.300 30.800 308.400 ;
        RECT 44.400 308.300 45.200 308.400 ;
        RECT 30.000 307.700 45.200 308.300 ;
        RECT 30.000 307.600 30.800 307.700 ;
        RECT 44.400 307.600 45.200 307.700 ;
        RECT 49.200 308.300 50.000 308.400 ;
        RECT 73.200 308.300 74.000 308.400 ;
        RECT 49.200 307.700 74.000 308.300 ;
        RECT 49.200 307.600 50.000 307.700 ;
        RECT 73.200 307.600 74.000 307.700 ;
        RECT 330.800 308.300 331.600 308.400 ;
        RECT 340.400 308.300 341.200 308.400 ;
        RECT 346.800 308.300 347.600 308.400 ;
        RECT 330.800 307.700 347.600 308.300 ;
        RECT 330.800 307.600 331.600 307.700 ;
        RECT 340.400 307.600 341.200 307.700 ;
        RECT 346.800 307.600 347.600 307.700 ;
        RECT 353.200 308.300 354.000 308.400 ;
        RECT 369.200 308.300 370.000 308.400 ;
        RECT 382.000 308.300 382.800 308.400 ;
        RECT 353.200 307.700 382.800 308.300 ;
        RECT 353.200 307.600 354.000 307.700 ;
        RECT 369.200 307.600 370.000 307.700 ;
        RECT 382.000 307.600 382.800 307.700 ;
        RECT 385.200 308.300 386.000 308.400 ;
        RECT 390.000 308.300 390.800 308.400 ;
        RECT 385.200 307.700 390.800 308.300 ;
        RECT 385.200 307.600 386.000 307.700 ;
        RECT 390.000 307.600 390.800 307.700 ;
        RECT 404.400 308.300 405.200 308.400 ;
        RECT 406.000 308.300 406.800 308.400 ;
        RECT 404.400 307.700 406.800 308.300 ;
        RECT 404.400 307.600 405.200 307.700 ;
        RECT 406.000 307.600 406.800 307.700 ;
        RECT 407.600 308.300 408.400 308.400 ;
        RECT 412.400 308.300 413.200 308.400 ;
        RECT 407.600 307.700 413.200 308.300 ;
        RECT 407.600 307.600 408.400 307.700 ;
        RECT 412.400 307.600 413.200 307.700 ;
        RECT 439.600 308.300 440.400 308.400 ;
        RECT 454.000 308.300 454.800 308.400 ;
        RECT 439.600 307.700 454.800 308.300 ;
        RECT 439.600 307.600 440.400 307.700 ;
        RECT 454.000 307.600 454.800 307.700 ;
        RECT 508.400 308.300 509.200 308.400 ;
        RECT 513.200 308.300 514.000 308.400 ;
        RECT 521.200 308.300 522.000 308.400 ;
        RECT 526.000 308.300 526.800 308.400 ;
        RECT 508.400 307.700 526.800 308.300 ;
        RECT 508.400 307.600 509.200 307.700 ;
        RECT 513.200 307.600 514.000 307.700 ;
        RECT 521.200 307.600 522.000 307.700 ;
        RECT 526.000 307.600 526.800 307.700 ;
        RECT 529.200 308.300 530.000 308.400 ;
        RECT 535.600 308.300 536.400 308.400 ;
        RECT 529.200 307.700 536.400 308.300 ;
        RECT 529.200 307.600 530.000 307.700 ;
        RECT 535.600 307.600 536.400 307.700 ;
        RECT 4.400 306.300 5.200 306.400 ;
        RECT 14.000 306.300 14.800 306.400 ;
        RECT 22.000 306.300 22.800 306.400 ;
        RECT 4.400 305.700 22.800 306.300 ;
        RECT 4.400 305.600 5.200 305.700 ;
        RECT 14.000 305.600 14.800 305.700 ;
        RECT 22.000 305.600 22.800 305.700 ;
        RECT 33.200 306.300 34.000 306.400 ;
        RECT 34.800 306.300 35.600 306.400 ;
        RECT 50.800 306.300 51.600 306.400 ;
        RECT 33.200 305.700 51.600 306.300 ;
        RECT 33.200 305.600 34.000 305.700 ;
        RECT 34.800 305.600 35.600 305.700 ;
        RECT 50.800 305.600 51.600 305.700 ;
        RECT 66.800 306.300 67.600 306.400 ;
        RECT 76.400 306.300 77.200 306.400 ;
        RECT 79.600 306.300 80.400 306.400 ;
        RECT 66.800 305.700 80.400 306.300 ;
        RECT 66.800 305.600 67.600 305.700 ;
        RECT 76.400 305.600 77.200 305.700 ;
        RECT 79.600 305.600 80.400 305.700 ;
        RECT 87.600 306.300 88.400 306.400 ;
        RECT 92.400 306.300 93.200 306.400 ;
        RECT 87.600 305.700 93.200 306.300 ;
        RECT 87.600 305.600 88.400 305.700 ;
        RECT 92.400 305.600 93.200 305.700 ;
        RECT 111.600 306.300 112.400 306.400 ;
        RECT 122.800 306.300 123.600 306.400 ;
        RECT 111.600 305.700 123.600 306.300 ;
        RECT 111.600 305.600 112.400 305.700 ;
        RECT 122.800 305.600 123.600 305.700 ;
        RECT 135.600 306.300 136.400 306.400 ;
        RECT 161.200 306.300 162.000 306.400 ;
        RECT 135.600 305.700 162.000 306.300 ;
        RECT 135.600 305.600 136.400 305.700 ;
        RECT 161.200 305.600 162.000 305.700 ;
        RECT 175.600 306.300 176.400 306.400 ;
        RECT 177.200 306.300 178.000 306.400 ;
        RECT 180.400 306.300 181.200 306.400 ;
        RECT 175.600 305.700 181.200 306.300 ;
        RECT 175.600 305.600 176.400 305.700 ;
        RECT 177.200 305.600 178.000 305.700 ;
        RECT 180.400 305.600 181.200 305.700 ;
        RECT 191.600 306.300 192.400 306.400 ;
        RECT 220.400 306.300 221.200 306.400 ;
        RECT 191.600 305.700 221.200 306.300 ;
        RECT 191.600 305.600 192.400 305.700 ;
        RECT 220.400 305.600 221.200 305.700 ;
        RECT 238.000 306.300 238.800 306.400 ;
        RECT 247.600 306.300 248.400 306.400 ;
        RECT 238.000 305.700 248.400 306.300 ;
        RECT 238.000 305.600 238.800 305.700 ;
        RECT 247.600 305.600 248.400 305.700 ;
        RECT 340.400 306.300 341.200 306.400 ;
        RECT 351.600 306.300 352.400 306.400 ;
        RECT 340.400 305.700 352.400 306.300 ;
        RECT 340.400 305.600 341.200 305.700 ;
        RECT 351.600 305.600 352.400 305.700 ;
        RECT 364.400 306.300 365.200 306.400 ;
        RECT 375.600 306.300 376.400 306.400 ;
        RECT 364.400 305.700 376.400 306.300 ;
        RECT 364.400 305.600 365.200 305.700 ;
        RECT 375.600 305.600 376.400 305.700 ;
        RECT 377.200 306.300 378.000 306.400 ;
        RECT 399.600 306.300 400.400 306.400 ;
        RECT 377.200 305.700 400.400 306.300 ;
        RECT 377.200 305.600 378.000 305.700 ;
        RECT 399.600 305.600 400.400 305.700 ;
        RECT 430.000 306.300 430.800 306.400 ;
        RECT 444.400 306.300 445.200 306.400 ;
        RECT 430.000 305.700 445.200 306.300 ;
        RECT 430.000 305.600 430.800 305.700 ;
        RECT 444.400 305.600 445.200 305.700 ;
        RECT 457.200 306.300 458.000 306.400 ;
        RECT 468.400 306.300 469.200 306.400 ;
        RECT 474.800 306.300 475.600 306.400 ;
        RECT 457.200 305.700 475.600 306.300 ;
        RECT 457.200 305.600 458.000 305.700 ;
        RECT 468.400 305.600 469.200 305.700 ;
        RECT 474.800 305.600 475.600 305.700 ;
        RECT 494.000 306.300 494.800 306.400 ;
        RECT 497.200 306.300 498.000 306.400 ;
        RECT 503.600 306.300 504.400 306.400 ;
        RECT 494.000 305.700 504.400 306.300 ;
        RECT 494.000 305.600 494.800 305.700 ;
        RECT 497.200 305.600 498.000 305.700 ;
        RECT 503.600 305.600 504.400 305.700 ;
        RECT 10.800 304.300 11.600 304.400 ;
        RECT 33.200 304.300 34.000 304.400 ;
        RECT 10.800 303.700 34.000 304.300 ;
        RECT 10.800 303.600 11.600 303.700 ;
        RECT 33.200 303.600 34.000 303.700 ;
        RECT 46.000 304.300 46.800 304.400 ;
        RECT 54.000 304.300 54.800 304.400 ;
        RECT 46.000 303.700 54.800 304.300 ;
        RECT 46.000 303.600 46.800 303.700 ;
        RECT 54.000 303.600 54.800 303.700 ;
        RECT 65.200 304.300 66.000 304.400 ;
        RECT 68.400 304.300 69.200 304.400 ;
        RECT 65.200 303.700 69.200 304.300 ;
        RECT 65.200 303.600 66.000 303.700 ;
        RECT 68.400 303.600 69.200 303.700 ;
        RECT 71.600 304.300 72.400 304.400 ;
        RECT 74.800 304.300 75.600 304.400 ;
        RECT 71.600 303.700 75.600 304.300 ;
        RECT 71.600 303.600 72.400 303.700 ;
        RECT 74.800 303.600 75.600 303.700 ;
        RECT 130.800 304.300 131.600 304.400 ;
        RECT 156.400 304.300 157.200 304.400 ;
        RECT 250.800 304.300 251.600 304.400 ;
        RECT 258.800 304.300 259.600 304.400 ;
        RECT 130.800 303.700 142.700 304.300 ;
        RECT 130.800 303.600 131.600 303.700 ;
        RECT 39.600 302.300 40.400 302.400 ;
        RECT 62.000 302.300 62.800 302.400 ;
        RECT 39.600 301.700 62.800 302.300 ;
        RECT 39.600 301.600 40.400 301.700 ;
        RECT 62.000 301.600 62.800 301.700 ;
        RECT 66.800 302.300 67.600 302.400 ;
        RECT 71.600 302.300 72.400 302.400 ;
        RECT 66.800 301.700 72.400 302.300 ;
        RECT 142.100 302.300 142.700 303.700 ;
        RECT 156.400 303.700 259.600 304.300 ;
        RECT 156.400 303.600 157.200 303.700 ;
        RECT 250.800 303.600 251.600 303.700 ;
        RECT 258.800 303.600 259.600 303.700 ;
        RECT 346.800 304.300 347.600 304.400 ;
        RECT 361.200 304.300 362.000 304.400 ;
        RECT 346.800 303.700 362.000 304.300 ;
        RECT 346.800 303.600 347.600 303.700 ;
        RECT 361.200 303.600 362.000 303.700 ;
        RECT 362.800 304.300 363.600 304.400 ;
        RECT 366.000 304.300 366.800 304.400 ;
        RECT 372.400 304.300 373.200 304.400 ;
        RECT 362.800 303.700 373.200 304.300 ;
        RECT 362.800 303.600 363.600 303.700 ;
        RECT 366.000 303.600 366.800 303.700 ;
        RECT 372.400 303.600 373.200 303.700 ;
        RECT 431.600 304.300 432.400 304.400 ;
        RECT 439.600 304.300 440.400 304.400 ;
        RECT 431.600 303.700 440.400 304.300 ;
        RECT 431.600 303.600 432.400 303.700 ;
        RECT 439.600 303.600 440.400 303.700 ;
        RECT 490.800 304.300 491.600 304.400 ;
        RECT 503.600 304.300 504.400 304.400 ;
        RECT 506.800 304.300 507.600 304.400 ;
        RECT 537.200 304.300 538.000 304.400 ;
        RECT 490.800 303.700 538.000 304.300 ;
        RECT 490.800 303.600 491.600 303.700 ;
        RECT 503.600 303.600 504.400 303.700 ;
        RECT 506.800 303.600 507.600 303.700 ;
        RECT 537.200 303.600 538.000 303.700 ;
        RECT 169.200 302.300 170.000 302.400 ;
        RECT 178.800 302.300 179.600 302.400 ;
        RECT 185.200 302.300 186.000 302.400 ;
        RECT 142.100 301.700 186.000 302.300 ;
        RECT 66.800 301.600 67.600 301.700 ;
        RECT 71.600 301.600 72.400 301.700 ;
        RECT 169.200 301.600 170.000 301.700 ;
        RECT 178.800 301.600 179.600 301.700 ;
        RECT 185.200 301.600 186.000 301.700 ;
        RECT 199.600 302.300 200.400 302.400 ;
        RECT 202.800 302.300 203.600 302.400 ;
        RECT 199.600 301.700 203.600 302.300 ;
        RECT 199.600 301.600 200.400 301.700 ;
        RECT 202.800 301.600 203.600 301.700 ;
        RECT 305.200 302.300 306.000 302.400 ;
        RECT 318.000 302.300 318.800 302.400 ;
        RECT 305.200 301.700 318.800 302.300 ;
        RECT 305.200 301.600 306.000 301.700 ;
        RECT 318.000 301.600 318.800 301.700 ;
        RECT 505.200 302.300 506.000 302.400 ;
        RECT 511.600 302.300 512.400 302.400 ;
        RECT 505.200 301.700 512.400 302.300 ;
        RECT 505.200 301.600 506.000 301.700 ;
        RECT 511.600 301.600 512.400 301.700 ;
        RECT 42.800 300.300 43.600 300.400 ;
        RECT 49.200 300.300 50.000 300.400 ;
        RECT 42.800 299.700 50.000 300.300 ;
        RECT 42.800 299.600 43.600 299.700 ;
        RECT 49.200 299.600 50.000 299.700 ;
        RECT 52.400 300.300 53.200 300.400 ;
        RECT 57.200 300.300 58.000 300.400 ;
        RECT 52.400 299.700 58.000 300.300 ;
        RECT 52.400 299.600 53.200 299.700 ;
        RECT 57.200 299.600 58.000 299.700 ;
        RECT 119.600 300.300 120.400 300.400 ;
        RECT 132.400 300.300 133.200 300.400 ;
        RECT 134.000 300.300 134.800 300.400 ;
        RECT 119.600 299.700 134.800 300.300 ;
        RECT 119.600 299.600 120.400 299.700 ;
        RECT 132.400 299.600 133.200 299.700 ;
        RECT 134.000 299.600 134.800 299.700 ;
        RECT 180.400 300.300 181.200 300.400 ;
        RECT 201.200 300.300 202.000 300.400 ;
        RECT 180.400 299.700 202.000 300.300 ;
        RECT 180.400 299.600 181.200 299.700 ;
        RECT 201.200 299.600 202.000 299.700 ;
        RECT 343.600 300.300 344.400 300.400 ;
        RECT 390.000 300.300 390.800 300.400 ;
        RECT 409.200 300.300 410.000 300.400 ;
        RECT 343.600 299.700 410.000 300.300 ;
        RECT 343.600 299.600 344.400 299.700 ;
        RECT 390.000 299.600 390.800 299.700 ;
        RECT 409.200 299.600 410.000 299.700 ;
        RECT 460.400 300.300 461.200 300.400 ;
        RECT 465.200 300.300 466.000 300.400 ;
        RECT 460.400 299.700 466.000 300.300 ;
        RECT 460.400 299.600 461.200 299.700 ;
        RECT 465.200 299.600 466.000 299.700 ;
        RECT 500.400 300.300 501.200 300.400 ;
        RECT 524.400 300.300 525.200 300.400 ;
        RECT 532.400 300.300 533.200 300.400 ;
        RECT 500.400 299.700 533.200 300.300 ;
        RECT 500.400 299.600 501.200 299.700 ;
        RECT 524.400 299.600 525.200 299.700 ;
        RECT 532.400 299.600 533.200 299.700 ;
        RECT 18.800 298.300 19.600 298.400 ;
        RECT 33.200 298.300 34.000 298.400 ;
        RECT 18.800 297.700 34.000 298.300 ;
        RECT 18.800 297.600 19.600 297.700 ;
        RECT 33.200 297.600 34.000 297.700 ;
        RECT 108.400 298.300 109.200 298.400 ;
        RECT 119.600 298.300 120.400 298.400 ;
        RECT 108.400 297.700 120.400 298.300 ;
        RECT 108.400 297.600 109.200 297.700 ;
        RECT 119.600 297.600 120.400 297.700 ;
        RECT 162.800 298.300 163.600 298.400 ;
        RECT 242.800 298.300 243.600 298.400 ;
        RECT 162.800 297.700 243.600 298.300 ;
        RECT 162.800 297.600 163.600 297.700 ;
        RECT 242.800 297.600 243.600 297.700 ;
        RECT 246.000 298.300 246.800 298.400 ;
        RECT 292.400 298.300 293.200 298.400 ;
        RECT 330.800 298.300 331.600 298.400 ;
        RECT 334.000 298.300 334.800 298.400 ;
        RECT 246.000 297.700 334.800 298.300 ;
        RECT 246.000 297.600 246.800 297.700 ;
        RECT 292.400 297.600 293.200 297.700 ;
        RECT 330.800 297.600 331.600 297.700 ;
        RECT 334.000 297.600 334.800 297.700 ;
        RECT 345.200 298.300 346.000 298.400 ;
        RECT 346.800 298.300 347.600 298.400 ;
        RECT 345.200 297.700 347.600 298.300 ;
        RECT 345.200 297.600 346.000 297.700 ;
        RECT 346.800 297.600 347.600 297.700 ;
        RECT 359.600 298.300 360.400 298.400 ;
        RECT 374.000 298.300 374.800 298.400 ;
        RECT 359.600 297.700 374.800 298.300 ;
        RECT 359.600 297.600 360.400 297.700 ;
        RECT 374.000 297.600 374.800 297.700 ;
        RECT 378.800 298.300 379.600 298.400 ;
        RECT 383.600 298.300 384.400 298.400 ;
        RECT 396.400 298.300 397.200 298.400 ;
        RECT 378.800 297.700 397.200 298.300 ;
        RECT 378.800 297.600 379.600 297.700 ;
        RECT 383.600 297.600 384.400 297.700 ;
        RECT 396.400 297.600 397.200 297.700 ;
        RECT 398.000 298.300 398.800 298.400 ;
        RECT 438.000 298.300 438.800 298.400 ;
        RECT 398.000 297.700 438.800 298.300 ;
        RECT 398.000 297.600 398.800 297.700 ;
        RECT 438.000 297.600 438.800 297.700 ;
        RECT 494.000 298.300 494.800 298.400 ;
        RECT 502.000 298.300 502.800 298.400 ;
        RECT 510.000 298.300 510.800 298.400 ;
        RECT 494.000 297.700 510.800 298.300 ;
        RECT 494.000 297.600 494.800 297.700 ;
        RECT 502.000 297.600 502.800 297.700 ;
        RECT 510.000 297.600 510.800 297.700 ;
        RECT 12.400 296.300 13.200 296.400 ;
        RECT 14.000 296.300 14.800 296.400 ;
        RECT 18.800 296.300 19.600 296.400 ;
        RECT 12.400 295.700 19.600 296.300 ;
        RECT 12.400 295.600 13.200 295.700 ;
        RECT 14.000 295.600 14.800 295.700 ;
        RECT 18.800 295.600 19.600 295.700 ;
        RECT 20.400 296.300 21.200 296.400 ;
        RECT 36.400 296.300 37.200 296.400 ;
        RECT 41.200 296.300 42.000 296.400 ;
        RECT 20.400 295.700 42.000 296.300 ;
        RECT 20.400 295.600 21.200 295.700 ;
        RECT 36.400 295.600 37.200 295.700 ;
        RECT 41.200 295.600 42.000 295.700 ;
        RECT 55.600 296.300 56.400 296.400 ;
        RECT 74.800 296.300 75.600 296.400 ;
        RECT 90.800 296.300 91.600 296.400 ;
        RECT 55.600 295.700 91.600 296.300 ;
        RECT 55.600 295.600 56.400 295.700 ;
        RECT 74.800 295.600 75.600 295.700 ;
        RECT 90.800 295.600 91.600 295.700 ;
        RECT 198.000 296.300 198.800 296.400 ;
        RECT 212.400 296.300 213.200 296.400 ;
        RECT 198.000 295.700 213.200 296.300 ;
        RECT 198.000 295.600 198.800 295.700 ;
        RECT 212.400 295.600 213.200 295.700 ;
        RECT 218.800 296.300 219.600 296.400 ;
        RECT 234.800 296.300 235.600 296.400 ;
        RECT 218.800 295.700 235.600 296.300 ;
        RECT 218.800 295.600 219.600 295.700 ;
        RECT 234.800 295.600 235.600 295.700 ;
        RECT 266.800 296.300 267.600 296.400 ;
        RECT 292.400 296.300 293.200 296.400 ;
        RECT 266.800 295.700 293.200 296.300 ;
        RECT 266.800 295.600 267.600 295.700 ;
        RECT 292.400 295.600 293.200 295.700 ;
        RECT 295.600 296.300 296.400 296.400 ;
        RECT 366.000 296.300 366.800 296.400 ;
        RECT 295.600 295.700 366.800 296.300 ;
        RECT 295.600 295.600 296.400 295.700 ;
        RECT 366.000 295.600 366.800 295.700 ;
        RECT 369.200 296.300 370.000 296.400 ;
        RECT 385.200 296.300 386.000 296.400 ;
        RECT 369.200 295.700 386.000 296.300 ;
        RECT 396.500 296.300 397.100 297.600 ;
        RECT 415.600 296.300 416.400 296.400 ;
        RECT 492.400 296.300 493.200 296.400 ;
        RECT 396.500 295.700 416.400 296.300 ;
        RECT 369.200 295.600 370.000 295.700 ;
        RECT 385.200 295.600 386.000 295.700 ;
        RECT 415.600 295.600 416.400 295.700 ;
        RECT 449.300 295.700 493.200 296.300 ;
        RECT 449.300 294.400 449.900 295.700 ;
        RECT 492.400 295.600 493.200 295.700 ;
        RECT 498.800 296.300 499.600 296.400 ;
        RECT 518.000 296.300 518.800 296.400 ;
        RECT 535.600 296.300 536.400 296.400 ;
        RECT 498.800 295.700 536.400 296.300 ;
        RECT 498.800 295.600 499.600 295.700 ;
        RECT 518.000 295.600 518.800 295.700 ;
        RECT 535.600 295.600 536.400 295.700 ;
        RECT 33.200 294.300 34.000 294.400 ;
        RECT 70.000 294.300 70.800 294.400 ;
        RECT 33.200 293.700 70.800 294.300 ;
        RECT 33.200 293.600 34.000 293.700 ;
        RECT 70.000 293.600 70.800 293.700 ;
        RECT 153.200 294.300 154.000 294.400 ;
        RECT 158.000 294.300 158.800 294.400 ;
        RECT 159.600 294.300 160.400 294.400 ;
        RECT 164.400 294.300 165.200 294.400 ;
        RECT 153.200 293.700 165.200 294.300 ;
        RECT 153.200 293.600 154.000 293.700 ;
        RECT 158.000 293.600 158.800 293.700 ;
        RECT 159.600 293.600 160.400 293.700 ;
        RECT 164.400 293.600 165.200 293.700 ;
        RECT 186.800 294.300 187.600 294.400 ;
        RECT 191.600 294.300 192.400 294.400 ;
        RECT 198.000 294.300 198.800 294.400 ;
        RECT 186.800 293.700 198.800 294.300 ;
        RECT 186.800 293.600 187.600 293.700 ;
        RECT 191.600 293.600 192.400 293.700 ;
        RECT 198.000 293.600 198.800 293.700 ;
        RECT 204.400 294.300 205.200 294.400 ;
        RECT 223.600 294.300 224.400 294.400 ;
        RECT 231.600 294.300 232.400 294.400 ;
        RECT 239.600 294.300 240.400 294.400 ;
        RECT 204.400 293.700 240.400 294.300 ;
        RECT 204.400 293.600 205.200 293.700 ;
        RECT 223.600 293.600 224.400 293.700 ;
        RECT 231.600 293.600 232.400 293.700 ;
        RECT 239.600 293.600 240.400 293.700 ;
        RECT 311.600 294.300 312.400 294.400 ;
        RECT 337.200 294.300 338.000 294.400 ;
        RECT 311.600 293.700 338.000 294.300 ;
        RECT 311.600 293.600 312.400 293.700 ;
        RECT 337.200 293.600 338.000 293.700 ;
        RECT 346.800 294.300 347.600 294.400 ;
        RECT 353.200 294.300 354.000 294.400 ;
        RECT 346.800 293.700 354.000 294.300 ;
        RECT 346.800 293.600 347.600 293.700 ;
        RECT 353.200 293.600 354.000 293.700 ;
        RECT 367.600 294.300 368.400 294.400 ;
        RECT 377.200 294.300 378.000 294.400 ;
        RECT 367.600 293.700 378.000 294.300 ;
        RECT 367.600 293.600 368.400 293.700 ;
        RECT 377.200 293.600 378.000 293.700 ;
        RECT 394.800 294.300 395.600 294.400 ;
        RECT 399.600 294.300 400.400 294.400 ;
        RECT 394.800 293.700 400.400 294.300 ;
        RECT 394.800 293.600 395.600 293.700 ;
        RECT 399.600 293.600 400.400 293.700 ;
        RECT 436.400 294.300 437.200 294.400 ;
        RECT 449.200 294.300 450.000 294.400 ;
        RECT 436.400 293.700 450.000 294.300 ;
        RECT 436.400 293.600 437.200 293.700 ;
        RECT 449.200 293.600 450.000 293.700 ;
        RECT 478.000 294.300 478.800 294.400 ;
        RECT 489.200 294.300 490.000 294.400 ;
        RECT 478.000 293.700 490.000 294.300 ;
        RECT 478.000 293.600 478.800 293.700 ;
        RECT 489.200 293.600 490.000 293.700 ;
        RECT 503.600 294.300 504.400 294.400 ;
        RECT 516.400 294.300 517.200 294.400 ;
        RECT 503.600 293.700 517.200 294.300 ;
        RECT 503.600 293.600 504.400 293.700 ;
        RECT 516.400 293.600 517.200 293.700 ;
        RECT 10.800 292.300 11.600 292.400 ;
        RECT 22.000 292.300 22.800 292.400 ;
        RECT 38.000 292.300 38.800 292.400 ;
        RECT 10.800 291.700 38.800 292.300 ;
        RECT 10.800 291.600 11.600 291.700 ;
        RECT 22.000 291.600 22.800 291.700 ;
        RECT 38.000 291.600 38.800 291.700 ;
        RECT 68.400 292.300 69.200 292.400 ;
        RECT 82.800 292.300 83.600 292.400 ;
        RECT 68.400 291.700 83.600 292.300 ;
        RECT 68.400 291.600 69.200 291.700 ;
        RECT 82.800 291.600 83.600 291.700 ;
        RECT 116.400 292.300 117.200 292.400 ;
        RECT 126.000 292.300 126.800 292.400 ;
        RECT 116.400 291.700 126.800 292.300 ;
        RECT 116.400 291.600 117.200 291.700 ;
        RECT 126.000 291.600 126.800 291.700 ;
        RECT 137.200 292.300 138.000 292.400 ;
        RECT 142.000 292.300 142.800 292.400 ;
        RECT 137.200 291.700 142.800 292.300 ;
        RECT 137.200 291.600 138.000 291.700 ;
        RECT 142.000 291.600 142.800 291.700 ;
        RECT 150.000 292.300 150.800 292.400 ;
        RECT 154.800 292.300 155.600 292.400 ;
        RECT 150.000 291.700 155.600 292.300 ;
        RECT 150.000 291.600 150.800 291.700 ;
        RECT 154.800 291.600 155.600 291.700 ;
        RECT 191.600 292.300 192.400 292.400 ;
        RECT 196.400 292.300 197.200 292.400 ;
        RECT 191.600 291.700 197.200 292.300 ;
        RECT 191.600 291.600 192.400 291.700 ;
        RECT 196.400 291.600 197.200 291.700 ;
        RECT 202.800 292.300 203.600 292.400 ;
        RECT 220.400 292.300 221.200 292.400 ;
        RECT 228.400 292.300 229.200 292.400 ;
        RECT 236.400 292.300 237.200 292.400 ;
        RECT 202.800 291.700 237.200 292.300 ;
        RECT 202.800 291.600 203.600 291.700 ;
        RECT 220.400 291.600 221.200 291.700 ;
        RECT 228.400 291.600 229.200 291.700 ;
        RECT 236.400 291.600 237.200 291.700 ;
        RECT 241.200 291.600 242.000 292.400 ;
        RECT 249.200 292.300 250.000 292.400 ;
        RECT 263.600 292.300 264.400 292.400 ;
        RECT 249.200 291.700 264.400 292.300 ;
        RECT 249.200 291.600 250.000 291.700 ;
        RECT 263.600 291.600 264.400 291.700 ;
        RECT 327.600 292.300 328.400 292.400 ;
        RECT 337.200 292.300 338.000 292.400 ;
        RECT 375.600 292.300 376.400 292.400 ;
        RECT 383.600 292.300 384.400 292.400 ;
        RECT 327.600 291.700 374.700 292.300 ;
        RECT 327.600 291.600 328.400 291.700 ;
        RECT 337.200 291.600 338.000 291.700 ;
        RECT 2.800 290.300 3.600 290.400 ;
        RECT 6.000 290.300 6.800 290.400 ;
        RECT 14.000 290.300 14.800 290.400 ;
        RECT 2.800 289.700 14.800 290.300 ;
        RECT 2.800 289.600 3.600 289.700 ;
        RECT 6.000 289.600 6.800 289.700 ;
        RECT 14.000 289.600 14.800 289.700 ;
        RECT 122.800 290.300 123.600 290.400 ;
        RECT 132.400 290.300 133.200 290.400 ;
        RECT 122.800 289.700 133.200 290.300 ;
        RECT 122.800 289.600 123.600 289.700 ;
        RECT 132.400 289.600 133.200 289.700 ;
        RECT 174.000 290.300 174.800 290.400 ;
        RECT 190.000 290.300 190.800 290.400 ;
        RECT 174.000 289.700 190.800 290.300 ;
        RECT 174.000 289.600 174.800 289.700 ;
        RECT 190.000 289.600 190.800 289.700 ;
        RECT 201.200 290.300 202.000 290.400 ;
        RECT 207.600 290.300 208.400 290.400 ;
        RECT 214.000 290.300 214.800 290.400 ;
        RECT 201.200 289.700 214.800 290.300 ;
        RECT 201.200 289.600 202.000 289.700 ;
        RECT 207.600 289.600 208.400 289.700 ;
        RECT 214.000 289.600 214.800 289.700 ;
        RECT 233.200 290.300 234.000 290.400 ;
        RECT 234.800 290.300 235.600 290.400 ;
        RECT 233.200 289.700 235.600 290.300 ;
        RECT 233.200 289.600 234.000 289.700 ;
        RECT 234.800 289.600 235.600 289.700 ;
        RECT 247.600 290.300 248.400 290.400 ;
        RECT 266.800 290.300 267.600 290.400 ;
        RECT 247.600 289.700 267.600 290.300 ;
        RECT 247.600 289.600 248.400 289.700 ;
        RECT 266.800 289.600 267.600 289.700 ;
        RECT 335.600 290.300 336.400 290.400 ;
        RECT 340.400 290.300 341.200 290.400 ;
        RECT 345.200 290.300 346.000 290.400 ;
        RECT 335.600 289.700 346.000 290.300 ;
        RECT 374.100 290.300 374.700 291.700 ;
        RECT 375.600 291.700 384.400 292.300 ;
        RECT 375.600 291.600 376.400 291.700 ;
        RECT 383.600 291.600 384.400 291.700 ;
        RECT 385.200 292.300 386.000 292.400 ;
        RECT 396.400 292.300 397.200 292.400 ;
        RECT 385.200 291.700 397.200 292.300 ;
        RECT 385.200 291.600 386.000 291.700 ;
        RECT 396.400 291.600 397.200 291.700 ;
        RECT 414.000 292.300 414.800 292.400 ;
        RECT 418.800 292.300 419.600 292.400 ;
        RECT 414.000 291.700 419.600 292.300 ;
        RECT 414.000 291.600 414.800 291.700 ;
        RECT 418.800 291.600 419.600 291.700 ;
        RECT 422.000 292.300 422.800 292.400 ;
        RECT 431.600 292.300 432.400 292.400 ;
        RECT 422.000 291.700 432.400 292.300 ;
        RECT 422.000 291.600 422.800 291.700 ;
        RECT 431.600 291.600 432.400 291.700 ;
        RECT 471.600 292.300 472.400 292.400 ;
        RECT 495.600 292.300 496.400 292.400 ;
        RECT 471.600 291.700 496.400 292.300 ;
        RECT 471.600 291.600 472.400 291.700 ;
        RECT 495.600 291.600 496.400 291.700 ;
        RECT 498.800 292.300 499.600 292.400 ;
        RECT 500.400 292.300 501.200 292.400 ;
        RECT 498.800 291.700 501.200 292.300 ;
        RECT 498.800 291.600 499.600 291.700 ;
        RECT 500.400 291.600 501.200 291.700 ;
        RECT 519.600 292.300 520.400 292.400 ;
        RECT 522.800 292.300 523.600 292.400 ;
        RECT 519.600 291.700 523.600 292.300 ;
        RECT 519.600 291.600 520.400 291.700 ;
        RECT 522.800 291.600 523.600 291.700 ;
        RECT 375.600 290.300 376.400 290.400 ;
        RECT 377.200 290.300 378.000 290.400 ;
        RECT 388.400 290.300 389.200 290.400 ;
        RECT 374.100 289.700 389.200 290.300 ;
        RECT 335.600 289.600 336.400 289.700 ;
        RECT 340.400 289.600 341.200 289.700 ;
        RECT 345.200 289.600 346.000 289.700 ;
        RECT 375.600 289.600 376.400 289.700 ;
        RECT 377.200 289.600 378.000 289.700 ;
        RECT 388.400 289.600 389.200 289.700 ;
        RECT 399.600 290.300 400.400 290.400 ;
        RECT 401.200 290.300 402.000 290.400 ;
        RECT 399.600 289.700 402.000 290.300 ;
        RECT 399.600 289.600 400.400 289.700 ;
        RECT 401.200 289.600 402.000 289.700 ;
        RECT 407.600 289.600 408.400 290.400 ;
        RECT 18.800 288.300 19.600 288.400 ;
        RECT 25.200 288.300 26.000 288.400 ;
        RECT 34.800 288.300 35.600 288.400 ;
        RECT 18.800 287.700 35.600 288.300 ;
        RECT 18.800 287.600 19.600 287.700 ;
        RECT 25.200 287.600 26.000 287.700 ;
        RECT 34.800 287.600 35.600 287.700 ;
        RECT 129.200 288.300 130.000 288.400 ;
        RECT 148.400 288.300 149.200 288.400 ;
        RECT 129.200 287.700 149.200 288.300 ;
        RECT 129.200 287.600 130.000 287.700 ;
        RECT 148.400 287.600 149.200 287.700 ;
        RECT 169.200 288.300 170.000 288.400 ;
        RECT 182.000 288.300 182.800 288.400 ;
        RECT 169.200 287.700 182.800 288.300 ;
        RECT 169.200 287.600 170.000 287.700 ;
        RECT 182.000 287.600 182.800 287.700 ;
        RECT 231.600 288.300 232.400 288.400 ;
        RECT 244.400 288.300 245.200 288.400 ;
        RECT 231.600 287.700 245.200 288.300 ;
        RECT 231.600 287.600 232.400 287.700 ;
        RECT 244.400 287.600 245.200 287.700 ;
        RECT 329.200 288.300 330.000 288.400 ;
        RECT 356.400 288.300 357.200 288.400 ;
        RECT 372.400 288.300 373.200 288.400 ;
        RECT 382.000 288.300 382.800 288.400 ;
        RECT 391.600 288.300 392.400 288.400 ;
        RECT 402.800 288.300 403.600 288.400 ;
        RECT 329.200 287.700 403.600 288.300 ;
        RECT 329.200 287.600 330.000 287.700 ;
        RECT 356.400 287.600 357.200 287.700 ;
        RECT 372.400 287.600 373.200 287.700 ;
        RECT 382.000 287.600 382.800 287.700 ;
        RECT 391.600 287.600 392.400 287.700 ;
        RECT 402.800 287.600 403.600 287.700 ;
        RECT 39.600 286.300 40.400 286.400 ;
        RECT 44.400 286.300 45.200 286.400 ;
        RECT 39.600 285.700 45.200 286.300 ;
        RECT 39.600 285.600 40.400 285.700 ;
        RECT 44.400 285.600 45.200 285.700 ;
        RECT 110.000 286.300 110.800 286.400 ;
        RECT 329.300 286.300 329.900 287.600 ;
        RECT 110.000 285.700 329.900 286.300 ;
        RECT 380.400 286.300 381.200 286.400 ;
        RECT 388.400 286.300 389.200 286.400 ;
        RECT 393.200 286.300 394.000 286.400 ;
        RECT 380.400 285.700 394.000 286.300 ;
        RECT 110.000 285.600 110.800 285.700 ;
        RECT 380.400 285.600 381.200 285.700 ;
        RECT 388.400 285.600 389.200 285.700 ;
        RECT 393.200 285.600 394.000 285.700 ;
        RECT 428.400 286.300 429.200 286.400 ;
        RECT 454.000 286.300 454.800 286.400 ;
        RECT 428.400 285.700 454.800 286.300 ;
        RECT 428.400 285.600 429.200 285.700 ;
        RECT 454.000 285.600 454.800 285.700 ;
        RECT 74.800 284.300 75.600 284.400 ;
        RECT 102.000 284.300 102.800 284.400 ;
        RECT 74.800 283.700 102.800 284.300 ;
        RECT 74.800 283.600 75.600 283.700 ;
        RECT 102.000 283.600 102.800 283.700 ;
        RECT 108.400 284.300 109.200 284.400 ;
        RECT 134.000 284.300 134.800 284.400 ;
        RECT 108.400 283.700 134.800 284.300 ;
        RECT 108.400 283.600 109.200 283.700 ;
        RECT 134.000 283.600 134.800 283.700 ;
        RECT 135.600 284.300 136.400 284.400 ;
        RECT 162.800 284.300 163.600 284.400 ;
        RECT 135.600 283.700 163.600 284.300 ;
        RECT 135.600 283.600 136.400 283.700 ;
        RECT 162.800 283.600 163.600 283.700 ;
        RECT 172.400 284.300 173.200 284.400 ;
        RECT 193.200 284.300 194.000 284.400 ;
        RECT 172.400 283.700 194.000 284.300 ;
        RECT 172.400 283.600 173.200 283.700 ;
        RECT 193.200 283.600 194.000 283.700 ;
        RECT 206.000 284.300 206.800 284.400 ;
        RECT 276.400 284.300 277.200 284.400 ;
        RECT 206.000 283.700 277.200 284.300 ;
        RECT 206.000 283.600 206.800 283.700 ;
        RECT 276.400 283.600 277.200 283.700 ;
        RECT 446.000 284.300 446.800 284.400 ;
        RECT 452.400 284.300 453.200 284.400 ;
        RECT 446.000 283.700 453.200 284.300 ;
        RECT 446.000 283.600 446.800 283.700 ;
        RECT 452.400 283.600 453.200 283.700 ;
        RECT 18.800 282.300 19.600 282.400 ;
        RECT 55.600 282.300 56.400 282.400 ;
        RECT 18.800 281.700 56.400 282.300 ;
        RECT 18.800 281.600 19.600 281.700 ;
        RECT 55.600 281.600 56.400 281.700 ;
        RECT 167.600 282.300 168.400 282.400 ;
        RECT 178.800 282.300 179.600 282.400 ;
        RECT 254.000 282.300 254.800 282.400 ;
        RECT 167.600 281.700 254.800 282.300 ;
        RECT 167.600 281.600 168.400 281.700 ;
        RECT 178.800 281.600 179.600 281.700 ;
        RECT 254.000 281.600 254.800 281.700 ;
        RECT 527.600 282.300 528.400 282.400 ;
        RECT 530.800 282.300 531.600 282.400 ;
        RECT 527.600 281.700 531.600 282.300 ;
        RECT 527.600 281.600 528.400 281.700 ;
        RECT 530.800 281.600 531.600 281.700 ;
        RECT 170.800 280.300 171.600 280.400 ;
        RECT 185.200 280.300 186.000 280.400 ;
        RECT 170.800 279.700 186.000 280.300 ;
        RECT 170.800 279.600 171.600 279.700 ;
        RECT 185.200 279.600 186.000 279.700 ;
        RECT 225.200 279.600 226.000 280.400 ;
        RECT 281.200 280.300 282.000 280.400 ;
        RECT 282.800 280.300 283.600 280.400 ;
        RECT 295.600 280.300 296.400 280.400 ;
        RECT 306.800 280.300 307.600 280.400 ;
        RECT 281.200 279.700 307.600 280.300 ;
        RECT 281.200 279.600 282.000 279.700 ;
        RECT 282.800 279.600 283.600 279.700 ;
        RECT 295.600 279.600 296.400 279.700 ;
        RECT 306.800 279.600 307.600 279.700 ;
        RECT 526.000 280.300 526.800 280.400 ;
        RECT 530.800 280.300 531.600 280.400 ;
        RECT 526.000 279.700 531.600 280.300 ;
        RECT 526.000 279.600 526.800 279.700 ;
        RECT 530.800 279.600 531.600 279.700 ;
        RECT 23.600 277.600 24.400 278.400 ;
        RECT 158.000 278.300 158.800 278.400 ;
        RECT 174.000 278.300 174.800 278.400 ;
        RECT 158.000 277.700 174.800 278.300 ;
        RECT 158.000 277.600 158.800 277.700 ;
        RECT 174.000 277.600 174.800 277.700 ;
        RECT 188.400 278.300 189.200 278.400 ;
        RECT 207.600 278.300 208.400 278.400 ;
        RECT 188.400 277.700 208.400 278.300 ;
        RECT 188.400 277.600 189.200 277.700 ;
        RECT 207.600 277.600 208.400 277.700 ;
        RECT 489.200 278.300 490.000 278.400 ;
        RECT 497.200 278.300 498.000 278.400 ;
        RECT 489.200 277.700 498.000 278.300 ;
        RECT 489.200 277.600 490.000 277.700 ;
        RECT 497.200 277.600 498.000 277.700 ;
        RECT 30.000 276.300 30.800 276.400 ;
        RECT 47.600 276.300 48.400 276.400 ;
        RECT 30.000 275.700 48.400 276.300 ;
        RECT 30.000 275.600 30.800 275.700 ;
        RECT 47.600 275.600 48.400 275.700 ;
        RECT 145.200 276.300 146.000 276.400 ;
        RECT 174.000 276.300 174.800 276.400 ;
        RECT 145.200 275.700 174.800 276.300 ;
        RECT 145.200 275.600 146.000 275.700 ;
        RECT 174.000 275.600 174.800 275.700 ;
        RECT 206.000 276.300 206.800 276.400 ;
        RECT 215.600 276.300 216.400 276.400 ;
        RECT 206.000 275.700 216.400 276.300 ;
        RECT 206.000 275.600 206.800 275.700 ;
        RECT 215.600 275.600 216.400 275.700 ;
        RECT 295.600 276.300 296.400 276.400 ;
        RECT 354.800 276.300 355.600 276.400 ;
        RECT 422.000 276.300 422.800 276.400 ;
        RECT 295.600 275.700 422.800 276.300 ;
        RECT 295.600 275.600 296.400 275.700 ;
        RECT 354.800 275.600 355.600 275.700 ;
        RECT 422.000 275.600 422.800 275.700 ;
        RECT 22.000 274.300 22.800 274.400 ;
        RECT 38.000 274.300 38.800 274.400 ;
        RECT 22.000 273.700 38.800 274.300 ;
        RECT 22.000 273.600 22.800 273.700 ;
        RECT 38.000 273.600 38.800 273.700 ;
        RECT 150.000 274.300 150.800 274.400 ;
        RECT 161.200 274.300 162.000 274.400 ;
        RECT 150.000 273.700 162.000 274.300 ;
        RECT 150.000 273.600 150.800 273.700 ;
        RECT 161.200 273.600 162.000 273.700 ;
        RECT 167.600 274.300 168.400 274.400 ;
        RECT 172.400 274.300 173.200 274.400 ;
        RECT 167.600 273.700 173.200 274.300 ;
        RECT 167.600 273.600 168.400 273.700 ;
        RECT 172.400 273.600 173.200 273.700 ;
        RECT 175.600 274.300 176.400 274.400 ;
        RECT 186.800 274.300 187.600 274.400 ;
        RECT 175.600 273.700 187.600 274.300 ;
        RECT 175.600 273.600 176.400 273.700 ;
        RECT 186.800 273.600 187.600 273.700 ;
        RECT 190.000 274.300 190.800 274.400 ;
        RECT 193.200 274.300 194.000 274.400 ;
        RECT 190.000 273.700 194.000 274.300 ;
        RECT 190.000 273.600 190.800 273.700 ;
        RECT 193.200 273.600 194.000 273.700 ;
        RECT 199.600 274.300 200.400 274.400 ;
        RECT 210.800 274.300 211.600 274.400 ;
        RECT 199.600 273.700 211.600 274.300 ;
        RECT 199.600 273.600 200.400 273.700 ;
        RECT 210.800 273.600 211.600 273.700 ;
        RECT 234.800 274.300 235.600 274.400 ;
        RECT 238.000 274.300 238.800 274.400 ;
        RECT 234.800 273.700 238.800 274.300 ;
        RECT 234.800 273.600 235.600 273.700 ;
        RECT 238.000 273.600 238.800 273.700 ;
        RECT 242.800 274.300 243.600 274.400 ;
        RECT 247.600 274.300 248.400 274.400 ;
        RECT 335.600 274.300 336.400 274.400 ;
        RECT 353.200 274.300 354.000 274.400 ;
        RECT 242.800 273.700 354.000 274.300 ;
        RECT 242.800 273.600 243.600 273.700 ;
        RECT 247.600 273.600 248.400 273.700 ;
        RECT 335.600 273.600 336.400 273.700 ;
        RECT 353.200 273.600 354.000 273.700 ;
        RECT 28.400 272.300 29.200 272.400 ;
        RECT 30.000 272.300 30.800 272.400 ;
        RECT 28.400 271.700 30.800 272.300 ;
        RECT 28.400 271.600 29.200 271.700 ;
        RECT 30.000 271.600 30.800 271.700 ;
        RECT 36.400 272.300 37.200 272.400 ;
        RECT 47.600 272.300 48.400 272.400 ;
        RECT 36.400 271.700 48.400 272.300 ;
        RECT 36.400 271.600 37.200 271.700 ;
        RECT 47.600 271.600 48.400 271.700 ;
        RECT 60.400 272.300 61.200 272.400 ;
        RECT 65.200 272.300 66.000 272.400 ;
        RECT 70.000 272.300 70.800 272.400 ;
        RECT 60.400 271.700 70.800 272.300 ;
        RECT 60.400 271.600 61.200 271.700 ;
        RECT 65.200 271.600 66.000 271.700 ;
        RECT 70.000 271.600 70.800 271.700 ;
        RECT 114.800 272.300 115.600 272.400 ;
        RECT 145.200 272.300 146.000 272.400 ;
        RECT 180.400 272.300 181.200 272.400 ;
        RECT 202.800 272.300 203.600 272.400 ;
        RECT 114.800 271.700 203.600 272.300 ;
        RECT 114.800 271.600 115.600 271.700 ;
        RECT 145.200 271.600 146.000 271.700 ;
        RECT 180.400 271.600 181.200 271.700 ;
        RECT 202.800 271.600 203.600 271.700 ;
        RECT 209.200 272.300 210.000 272.400 ;
        RECT 225.200 272.300 226.000 272.400 ;
        RECT 209.200 271.700 226.000 272.300 ;
        RECT 209.200 271.600 210.000 271.700 ;
        RECT 225.200 271.600 226.000 271.700 ;
        RECT 252.400 272.300 253.200 272.400 ;
        RECT 255.600 272.300 256.400 272.400 ;
        RECT 252.400 271.700 256.400 272.300 ;
        RECT 252.400 271.600 253.200 271.700 ;
        RECT 255.600 271.600 256.400 271.700 ;
        RECT 338.800 272.300 339.600 272.400 ;
        RECT 346.800 272.300 347.600 272.400 ;
        RECT 338.800 271.700 347.600 272.300 ;
        RECT 338.800 271.600 339.600 271.700 ;
        RECT 346.800 271.600 347.600 271.700 ;
        RECT 407.600 272.300 408.400 272.400 ;
        RECT 486.000 272.300 486.800 272.400 ;
        RECT 407.600 271.700 486.800 272.300 ;
        RECT 407.600 271.600 408.400 271.700 ;
        RECT 486.000 271.600 486.800 271.700 ;
        RECT 38.000 270.300 38.800 270.400 ;
        RECT 39.600 270.300 40.400 270.400 ;
        RECT 38.000 269.700 40.400 270.300 ;
        RECT 38.000 269.600 38.800 269.700 ;
        RECT 39.600 269.600 40.400 269.700 ;
        RECT 52.400 270.300 53.200 270.400 ;
        RECT 55.600 270.300 56.400 270.400 ;
        RECT 52.400 269.700 56.400 270.300 ;
        RECT 52.400 269.600 53.200 269.700 ;
        RECT 55.600 269.600 56.400 269.700 ;
        RECT 63.600 270.300 64.400 270.400 ;
        RECT 73.200 270.300 74.000 270.400 ;
        RECT 63.600 269.700 74.000 270.300 ;
        RECT 63.600 269.600 64.400 269.700 ;
        RECT 73.200 269.600 74.000 269.700 ;
        RECT 135.600 270.300 136.400 270.400 ;
        RECT 138.800 270.300 139.600 270.400 ;
        RECT 135.600 269.700 139.600 270.300 ;
        RECT 135.600 269.600 136.400 269.700 ;
        RECT 138.800 269.600 139.600 269.700 ;
        RECT 142.000 269.600 142.800 270.400 ;
        RECT 156.400 270.300 157.200 270.400 ;
        RECT 166.000 270.300 166.800 270.400 ;
        RECT 156.400 269.700 166.800 270.300 ;
        RECT 156.400 269.600 157.200 269.700 ;
        RECT 166.000 269.600 166.800 269.700 ;
        RECT 177.200 270.300 178.000 270.400 ;
        RECT 182.000 270.300 182.800 270.400 ;
        RECT 177.200 269.700 182.800 270.300 ;
        RECT 177.200 269.600 178.000 269.700 ;
        RECT 182.000 269.600 182.800 269.700 ;
        RECT 188.400 270.300 189.200 270.400 ;
        RECT 193.200 270.300 194.000 270.400 ;
        RECT 188.400 269.700 194.000 270.300 ;
        RECT 188.400 269.600 189.200 269.700 ;
        RECT 193.200 269.600 194.000 269.700 ;
        RECT 194.800 270.300 195.600 270.400 ;
        RECT 198.000 270.300 198.800 270.400 ;
        RECT 202.800 270.300 203.600 270.400 ;
        RECT 194.800 269.700 203.600 270.300 ;
        RECT 194.800 269.600 195.600 269.700 ;
        RECT 198.000 269.600 198.800 269.700 ;
        RECT 202.800 269.600 203.600 269.700 ;
        RECT 226.800 270.300 227.600 270.400 ;
        RECT 236.400 270.300 237.200 270.400 ;
        RECT 226.800 269.700 237.200 270.300 ;
        RECT 226.800 269.600 227.600 269.700 ;
        RECT 236.400 269.600 237.200 269.700 ;
        RECT 250.800 270.300 251.600 270.400 ;
        RECT 254.000 270.300 254.800 270.400 ;
        RECT 250.800 269.700 254.800 270.300 ;
        RECT 250.800 269.600 251.600 269.700 ;
        RECT 254.000 269.600 254.800 269.700 ;
        RECT 332.400 270.300 333.200 270.400 ;
        RECT 343.600 270.300 344.400 270.400 ;
        RECT 332.400 269.700 344.400 270.300 ;
        RECT 332.400 269.600 333.200 269.700 ;
        RECT 343.600 269.600 344.400 269.700 ;
        RECT 354.800 270.300 355.600 270.400 ;
        RECT 386.800 270.300 387.600 270.400 ;
        RECT 354.800 269.700 387.600 270.300 ;
        RECT 354.800 269.600 355.600 269.700 ;
        RECT 386.800 269.600 387.600 269.700 ;
        RECT 409.200 270.300 410.000 270.400 ;
        RECT 418.800 270.300 419.600 270.400 ;
        RECT 409.200 269.700 419.600 270.300 ;
        RECT 409.200 269.600 410.000 269.700 ;
        RECT 418.800 269.600 419.600 269.700 ;
        RECT 434.800 270.300 435.600 270.400 ;
        RECT 441.200 270.300 442.000 270.400 ;
        RECT 434.800 269.700 442.000 270.300 ;
        RECT 434.800 269.600 435.600 269.700 ;
        RECT 441.200 269.600 442.000 269.700 ;
        RECT 442.800 270.300 443.600 270.400 ;
        RECT 473.200 270.300 474.000 270.400 ;
        RECT 442.800 269.700 474.000 270.300 ;
        RECT 442.800 269.600 443.600 269.700 ;
        RECT 473.200 269.600 474.000 269.700 ;
        RECT 482.800 270.300 483.600 270.400 ;
        RECT 497.200 270.300 498.000 270.400 ;
        RECT 482.800 269.700 498.000 270.300 ;
        RECT 482.800 269.600 483.600 269.700 ;
        RECT 497.200 269.600 498.000 269.700 ;
        RECT 30.000 267.600 30.800 268.400 ;
        RECT 38.000 268.300 38.800 268.400 ;
        RECT 49.200 268.300 50.000 268.400 ;
        RECT 38.000 267.700 50.000 268.300 ;
        RECT 38.000 267.600 38.800 267.700 ;
        RECT 49.200 267.600 50.000 267.700 ;
        RECT 54.000 268.300 54.800 268.400 ;
        RECT 60.400 268.300 61.200 268.400 ;
        RECT 54.000 267.700 61.200 268.300 ;
        RECT 54.000 267.600 54.800 267.700 ;
        RECT 60.400 267.600 61.200 267.700 ;
        RECT 68.400 268.300 69.200 268.400 ;
        RECT 74.800 268.300 75.600 268.400 ;
        RECT 86.000 268.300 86.800 268.400 ;
        RECT 68.400 267.700 86.800 268.300 ;
        RECT 68.400 267.600 69.200 267.700 ;
        RECT 74.800 267.600 75.600 267.700 ;
        RECT 86.000 267.600 86.800 267.700 ;
        RECT 122.800 268.300 123.600 268.400 ;
        RECT 132.400 268.300 133.200 268.400 ;
        RECT 148.400 268.300 149.200 268.400 ;
        RECT 122.800 267.700 149.200 268.300 ;
        RECT 122.800 267.600 123.600 267.700 ;
        RECT 132.400 267.600 133.200 267.700 ;
        RECT 148.400 267.600 149.200 267.700 ;
        RECT 151.600 268.300 152.400 268.400 ;
        RECT 154.800 268.300 155.600 268.400 ;
        RECT 151.600 267.700 155.600 268.300 ;
        RECT 151.600 267.600 152.400 267.700 ;
        RECT 154.800 267.600 155.600 267.700 ;
        RECT 162.800 268.300 163.600 268.400 ;
        RECT 175.600 268.300 176.400 268.400 ;
        RECT 162.800 267.700 176.400 268.300 ;
        RECT 162.800 267.600 163.600 267.700 ;
        RECT 175.600 267.600 176.400 267.700 ;
        RECT 177.200 268.300 178.000 268.400 ;
        RECT 231.600 268.300 232.400 268.400 ;
        RECT 177.200 267.700 232.400 268.300 ;
        RECT 177.200 267.600 178.000 267.700 ;
        RECT 231.600 267.600 232.400 267.700 ;
        RECT 244.400 268.300 245.200 268.400 ;
        RECT 270.000 268.300 270.800 268.400 ;
        RECT 244.400 267.700 270.800 268.300 ;
        RECT 244.400 267.600 245.200 267.700 ;
        RECT 270.000 267.600 270.800 267.700 ;
        RECT 289.200 267.600 290.000 268.400 ;
        RECT 396.400 268.300 397.200 268.400 ;
        RECT 436.400 268.300 437.200 268.400 ;
        RECT 396.400 267.700 437.200 268.300 ;
        RECT 396.400 267.600 397.200 267.700 ;
        RECT 436.400 267.600 437.200 267.700 ;
        RECT 439.600 268.300 440.400 268.400 ;
        RECT 449.200 268.300 450.000 268.400 ;
        RECT 479.600 268.300 480.400 268.400 ;
        RECT 439.600 267.700 480.400 268.300 ;
        RECT 439.600 267.600 440.400 267.700 ;
        RECT 449.200 267.600 450.000 267.700 ;
        RECT 479.600 267.600 480.400 267.700 ;
        RECT 508.400 268.300 509.200 268.400 ;
        RECT 514.800 268.300 515.600 268.400 ;
        RECT 508.400 267.700 515.600 268.300 ;
        RECT 508.400 267.600 509.200 267.700 ;
        RECT 514.800 267.600 515.600 267.700 ;
        RECT 36.400 266.300 37.200 266.400 ;
        RECT 44.400 266.300 45.200 266.400 ;
        RECT 46.000 266.300 46.800 266.400 ;
        RECT 36.400 265.700 46.800 266.300 ;
        RECT 36.400 265.600 37.200 265.700 ;
        RECT 44.400 265.600 45.200 265.700 ;
        RECT 46.000 265.600 46.800 265.700 ;
        RECT 55.600 265.600 56.400 266.400 ;
        RECT 68.400 266.300 69.200 266.400 ;
        RECT 71.600 266.300 72.400 266.400 ;
        RECT 68.400 265.700 72.400 266.300 ;
        RECT 68.400 265.600 69.200 265.700 ;
        RECT 71.600 265.600 72.400 265.700 ;
        RECT 74.800 266.300 75.600 266.400 ;
        RECT 87.600 266.300 88.400 266.400 ;
        RECT 74.800 265.700 88.400 266.300 ;
        RECT 74.800 265.600 75.600 265.700 ;
        RECT 87.600 265.600 88.400 265.700 ;
        RECT 134.000 266.300 134.800 266.400 ;
        RECT 178.800 266.300 179.600 266.400 ;
        RECT 134.000 265.700 179.600 266.300 ;
        RECT 134.000 265.600 134.800 265.700 ;
        RECT 178.800 265.600 179.600 265.700 ;
        RECT 193.200 266.300 194.000 266.400 ;
        RECT 206.000 266.300 206.800 266.400 ;
        RECT 210.800 266.300 211.600 266.400 ;
        RECT 193.200 265.700 211.600 266.300 ;
        RECT 193.200 265.600 194.000 265.700 ;
        RECT 206.000 265.600 206.800 265.700 ;
        RECT 210.800 265.600 211.600 265.700 ;
        RECT 214.000 266.300 214.800 266.400 ;
        RECT 220.400 266.300 221.200 266.400 ;
        RECT 226.800 266.300 227.600 266.400 ;
        RECT 214.000 265.700 227.600 266.300 ;
        RECT 214.000 265.600 214.800 265.700 ;
        RECT 220.400 265.600 221.200 265.700 ;
        RECT 226.800 265.600 227.600 265.700 ;
        RECT 242.800 266.300 243.600 266.400 ;
        RECT 247.600 266.300 248.400 266.400 ;
        RECT 242.800 265.700 248.400 266.300 ;
        RECT 242.800 265.600 243.600 265.700 ;
        RECT 247.600 265.600 248.400 265.700 ;
        RECT 249.200 266.300 250.000 266.400 ;
        RECT 258.800 266.300 259.600 266.400 ;
        RECT 249.200 265.700 259.600 266.300 ;
        RECT 249.200 265.600 250.000 265.700 ;
        RECT 258.800 265.600 259.600 265.700 ;
        RECT 260.400 266.300 261.200 266.400 ;
        RECT 289.200 266.300 290.000 266.400 ;
        RECT 302.000 266.300 302.800 266.400 ;
        RECT 260.400 265.700 302.800 266.300 ;
        RECT 260.400 265.600 261.200 265.700 ;
        RECT 289.200 265.600 290.000 265.700 ;
        RECT 302.000 265.600 302.800 265.700 ;
        RECT 308.400 266.300 309.200 266.400 ;
        RECT 319.600 266.300 320.400 266.400 ;
        RECT 364.400 266.300 365.200 266.400 ;
        RECT 399.600 266.300 400.400 266.400 ;
        RECT 308.400 265.700 400.400 266.300 ;
        RECT 308.400 265.600 309.200 265.700 ;
        RECT 319.600 265.600 320.400 265.700 ;
        RECT 364.400 265.600 365.200 265.700 ;
        RECT 399.600 265.600 400.400 265.700 ;
        RECT 417.200 266.300 418.000 266.400 ;
        RECT 430.000 266.300 430.800 266.400 ;
        RECT 417.200 265.700 430.800 266.300 ;
        RECT 417.200 265.600 418.000 265.700 ;
        RECT 430.000 265.600 430.800 265.700 ;
        RECT 450.800 266.300 451.600 266.400 ;
        RECT 470.000 266.300 470.800 266.400 ;
        RECT 481.200 266.300 482.000 266.400 ;
        RECT 450.800 265.700 482.000 266.300 ;
        RECT 450.800 265.600 451.600 265.700 ;
        RECT 470.000 265.600 470.800 265.700 ;
        RECT 481.200 265.600 482.000 265.700 ;
        RECT 490.800 266.300 491.600 266.400 ;
        RECT 524.400 266.300 525.200 266.400 ;
        RECT 490.800 265.700 525.200 266.300 ;
        RECT 490.800 265.600 491.600 265.700 ;
        RECT 524.400 265.600 525.200 265.700 ;
        RECT 52.400 264.300 53.200 264.400 ;
        RECT 57.200 264.300 58.000 264.400 ;
        RECT 52.400 263.700 58.000 264.300 ;
        RECT 52.400 263.600 53.200 263.700 ;
        RECT 57.200 263.600 58.000 263.700 ;
        RECT 103.600 264.300 104.400 264.400 ;
        RECT 140.400 264.300 141.200 264.400 ;
        RECT 103.600 263.700 141.200 264.300 ;
        RECT 103.600 263.600 104.400 263.700 ;
        RECT 140.400 263.600 141.200 263.700 ;
        RECT 142.000 264.300 142.800 264.400 ;
        RECT 151.600 264.300 152.400 264.400 ;
        RECT 142.000 263.700 152.400 264.300 ;
        RECT 142.000 263.600 142.800 263.700 ;
        RECT 151.600 263.600 152.400 263.700 ;
        RECT 174.000 264.300 174.800 264.400 ;
        RECT 178.800 264.300 179.600 264.400 ;
        RECT 174.000 263.700 179.600 264.300 ;
        RECT 174.000 263.600 174.800 263.700 ;
        RECT 178.800 263.600 179.600 263.700 ;
        RECT 188.400 264.300 189.200 264.400 ;
        RECT 255.600 264.300 256.400 264.400 ;
        RECT 188.400 263.700 256.400 264.300 ;
        RECT 188.400 263.600 189.200 263.700 ;
        RECT 255.600 263.600 256.400 263.700 ;
        RECT 481.200 264.300 482.000 264.400 ;
        RECT 490.800 264.300 491.600 264.400 ;
        RECT 481.200 263.700 491.600 264.300 ;
        RECT 481.200 263.600 482.000 263.700 ;
        RECT 490.800 263.600 491.600 263.700 ;
        RECT 495.600 264.300 496.400 264.400 ;
        RECT 505.200 264.300 506.000 264.400 ;
        RECT 527.600 264.300 528.400 264.400 ;
        RECT 495.600 263.700 528.400 264.300 ;
        RECT 495.600 263.600 496.400 263.700 ;
        RECT 505.200 263.600 506.000 263.700 ;
        RECT 527.600 263.600 528.400 263.700 ;
        RECT 41.200 262.300 42.000 262.400 ;
        RECT 62.000 262.300 62.800 262.400 ;
        RECT 41.200 261.700 62.800 262.300 ;
        RECT 41.200 261.600 42.000 261.700 ;
        RECT 62.000 261.600 62.800 261.700 ;
        RECT 137.200 262.300 138.000 262.400 ;
        RECT 140.400 262.300 141.200 262.400 ;
        RECT 137.200 261.700 141.200 262.300 ;
        RECT 137.200 261.600 138.000 261.700 ;
        RECT 140.400 261.600 141.200 261.700 ;
        RECT 145.200 262.300 146.000 262.400 ;
        RECT 167.600 262.300 168.400 262.400 ;
        RECT 246.000 262.300 246.800 262.400 ;
        RECT 145.200 261.700 246.800 262.300 ;
        RECT 145.200 261.600 146.000 261.700 ;
        RECT 167.600 261.600 168.400 261.700 ;
        RECT 246.000 261.600 246.800 261.700 ;
        RECT 305.200 262.300 306.000 262.400 ;
        RECT 318.000 262.300 318.800 262.400 ;
        RECT 305.200 261.700 318.800 262.300 ;
        RECT 305.200 261.600 306.000 261.700 ;
        RECT 318.000 261.600 318.800 261.700 ;
        RECT 327.600 262.300 328.400 262.400 ;
        RECT 340.400 262.300 341.200 262.400 ;
        RECT 327.600 261.700 341.200 262.300 ;
        RECT 327.600 261.600 328.400 261.700 ;
        RECT 340.400 261.600 341.200 261.700 ;
        RECT 348.400 262.300 349.200 262.400 ;
        RECT 361.200 262.300 362.000 262.400 ;
        RECT 348.400 261.700 362.000 262.300 ;
        RECT 348.400 261.600 349.200 261.700 ;
        RECT 361.200 261.600 362.000 261.700 ;
        RECT 444.400 262.300 445.200 262.400 ;
        RECT 465.200 262.300 466.000 262.400 ;
        RECT 444.400 261.700 466.000 262.300 ;
        RECT 444.400 261.600 445.200 261.700 ;
        RECT 465.200 261.600 466.000 261.700 ;
        RECT 466.800 262.300 467.600 262.400 ;
        RECT 468.400 262.300 469.200 262.400 ;
        RECT 466.800 261.700 469.200 262.300 ;
        RECT 466.800 261.600 467.600 261.700 ;
        RECT 468.400 261.600 469.200 261.700 ;
        RECT 90.800 260.300 91.600 260.400 ;
        RECT 97.200 260.300 98.000 260.400 ;
        RECT 106.800 260.300 107.600 260.400 ;
        RECT 119.600 260.300 120.400 260.400 ;
        RECT 90.800 259.700 120.400 260.300 ;
        RECT 90.800 259.600 91.600 259.700 ;
        RECT 97.200 259.600 98.000 259.700 ;
        RECT 106.800 259.600 107.600 259.700 ;
        RECT 119.600 259.600 120.400 259.700 ;
        RECT 166.000 260.300 166.800 260.400 ;
        RECT 167.600 260.300 168.400 260.400 ;
        RECT 166.000 259.700 168.400 260.300 ;
        RECT 166.000 259.600 166.800 259.700 ;
        RECT 167.600 259.600 168.400 259.700 ;
        RECT 174.000 260.300 174.800 260.400 ;
        RECT 252.400 260.300 253.200 260.400 ;
        RECT 174.000 259.700 253.200 260.300 ;
        RECT 174.000 259.600 174.800 259.700 ;
        RECT 252.400 259.600 253.200 259.700 ;
        RECT 286.000 260.300 286.800 260.400 ;
        RECT 305.200 260.300 306.000 260.400 ;
        RECT 310.000 260.300 310.800 260.400 ;
        RECT 286.000 259.700 310.800 260.300 ;
        RECT 286.000 259.600 286.800 259.700 ;
        RECT 305.200 259.600 306.000 259.700 ;
        RECT 310.000 259.600 310.800 259.700 ;
        RECT 316.400 260.300 317.200 260.400 ;
        RECT 322.800 260.300 323.600 260.400 ;
        RECT 316.400 259.700 323.600 260.300 ;
        RECT 316.400 259.600 317.200 259.700 ;
        RECT 322.800 259.600 323.600 259.700 ;
        RECT 337.200 260.300 338.000 260.400 ;
        RECT 342.000 260.300 342.800 260.400 ;
        RECT 375.600 260.300 376.400 260.400 ;
        RECT 337.200 259.700 376.400 260.300 ;
        RECT 337.200 259.600 338.000 259.700 ;
        RECT 342.000 259.600 342.800 259.700 ;
        RECT 375.600 259.600 376.400 259.700 ;
        RECT 446.000 260.300 446.800 260.400 ;
        RECT 447.600 260.300 448.400 260.400 ;
        RECT 446.000 259.700 448.400 260.300 ;
        RECT 446.000 259.600 446.800 259.700 ;
        RECT 447.600 259.600 448.400 259.700 ;
        RECT 23.600 257.600 24.400 258.400 ;
        RECT 42.800 258.300 43.600 258.400 ;
        RECT 73.200 258.300 74.000 258.400 ;
        RECT 42.800 257.700 74.000 258.300 ;
        RECT 42.800 257.600 43.600 257.700 ;
        RECT 73.200 257.600 74.000 257.700 ;
        RECT 177.200 258.300 178.000 258.400 ;
        RECT 193.200 258.300 194.000 258.400 ;
        RECT 177.200 257.700 194.000 258.300 ;
        RECT 177.200 257.600 178.000 257.700 ;
        RECT 193.200 257.600 194.000 257.700 ;
        RECT 201.200 258.300 202.000 258.400 ;
        RECT 207.600 258.300 208.400 258.400 ;
        RECT 214.000 258.300 214.800 258.400 ;
        RECT 201.200 257.700 214.800 258.300 ;
        RECT 201.200 257.600 202.000 257.700 ;
        RECT 207.600 257.600 208.400 257.700 ;
        RECT 214.000 257.600 214.800 257.700 ;
        RECT 241.200 258.300 242.000 258.400 ;
        RECT 340.400 258.300 341.200 258.400 ;
        RECT 380.400 258.300 381.200 258.400 ;
        RECT 382.000 258.300 382.800 258.400 ;
        RECT 241.200 257.700 382.800 258.300 ;
        RECT 241.200 257.600 242.000 257.700 ;
        RECT 340.400 257.600 341.200 257.700 ;
        RECT 380.400 257.600 381.200 257.700 ;
        RECT 382.000 257.600 382.800 257.700 ;
        RECT 433.200 258.300 434.000 258.400 ;
        RECT 455.600 258.300 456.400 258.400 ;
        RECT 473.200 258.300 474.000 258.400 ;
        RECT 433.200 257.700 474.000 258.300 ;
        RECT 433.200 257.600 434.000 257.700 ;
        RECT 455.600 257.600 456.400 257.700 ;
        RECT 473.200 257.600 474.000 257.700 ;
        RECT 481.200 258.300 482.000 258.400 ;
        RECT 542.000 258.300 542.800 258.400 ;
        RECT 546.800 258.300 547.600 258.400 ;
        RECT 481.200 257.700 547.600 258.300 ;
        RECT 481.200 257.600 482.000 257.700 ;
        RECT 542.000 257.600 542.800 257.700 ;
        RECT 546.800 257.600 547.600 257.700 ;
        RECT 1.200 256.300 2.000 256.400 ;
        RECT 9.200 256.300 10.000 256.400 ;
        RECT 14.000 256.300 14.800 256.400 ;
        RECT 1.200 255.700 14.800 256.300 ;
        RECT 1.200 255.600 2.000 255.700 ;
        RECT 9.200 255.600 10.000 255.700 ;
        RECT 14.000 255.600 14.800 255.700 ;
        RECT 31.600 256.300 32.400 256.400 ;
        RECT 33.200 256.300 34.000 256.400 ;
        RECT 31.600 255.700 34.000 256.300 ;
        RECT 31.600 255.600 32.400 255.700 ;
        RECT 33.200 255.600 34.000 255.700 ;
        RECT 41.200 256.300 42.000 256.400 ;
        RECT 44.400 256.300 45.200 256.400 ;
        RECT 41.200 255.700 45.200 256.300 ;
        RECT 41.200 255.600 42.000 255.700 ;
        RECT 44.400 255.600 45.200 255.700 ;
        RECT 46.000 255.600 46.800 256.400 ;
        RECT 63.600 256.300 64.400 256.400 ;
        RECT 76.400 256.300 77.200 256.400 ;
        RECT 81.200 256.300 82.000 256.400 ;
        RECT 63.600 255.700 82.000 256.300 ;
        RECT 63.600 255.600 64.400 255.700 ;
        RECT 76.400 255.600 77.200 255.700 ;
        RECT 81.200 255.600 82.000 255.700 ;
        RECT 132.400 256.300 133.200 256.400 ;
        RECT 143.600 256.300 144.400 256.400 ;
        RECT 158.000 256.300 158.800 256.400 ;
        RECT 132.400 255.700 158.800 256.300 ;
        RECT 132.400 255.600 133.200 255.700 ;
        RECT 143.600 255.600 144.400 255.700 ;
        RECT 158.000 255.600 158.800 255.700 ;
        RECT 185.200 256.300 186.000 256.400 ;
        RECT 194.800 256.300 195.600 256.400 ;
        RECT 185.200 255.700 195.600 256.300 ;
        RECT 185.200 255.600 186.000 255.700 ;
        RECT 194.800 255.600 195.600 255.700 ;
        RECT 206.000 256.300 206.800 256.400 ;
        RECT 209.200 256.300 210.000 256.400 ;
        RECT 206.000 255.700 210.000 256.300 ;
        RECT 206.000 255.600 206.800 255.700 ;
        RECT 209.200 255.600 210.000 255.700 ;
        RECT 223.600 256.300 224.400 256.400 ;
        RECT 263.600 256.300 264.400 256.400 ;
        RECT 286.000 256.300 286.800 256.400 ;
        RECT 223.600 255.700 286.800 256.300 ;
        RECT 223.600 255.600 224.400 255.700 ;
        RECT 263.600 255.600 264.400 255.700 ;
        RECT 286.000 255.600 286.800 255.700 ;
        RECT 289.200 256.300 290.000 256.400 ;
        RECT 321.200 256.300 322.000 256.400 ;
        RECT 289.200 255.700 322.000 256.300 ;
        RECT 289.200 255.600 290.000 255.700 ;
        RECT 321.200 255.600 322.000 255.700 ;
        RECT 346.800 256.300 347.600 256.400 ;
        RECT 362.800 256.300 363.600 256.400 ;
        RECT 346.800 255.700 363.600 256.300 ;
        RECT 346.800 255.600 347.600 255.700 ;
        RECT 362.800 255.600 363.600 255.700 ;
        RECT 366.000 256.300 366.800 256.400 ;
        RECT 394.800 256.300 395.600 256.400 ;
        RECT 406.000 256.300 406.800 256.400 ;
        RECT 450.800 256.300 451.600 256.400 ;
        RECT 366.000 255.700 451.600 256.300 ;
        RECT 366.000 255.600 366.800 255.700 ;
        RECT 394.800 255.600 395.600 255.700 ;
        RECT 406.000 255.600 406.800 255.700 ;
        RECT 450.800 255.600 451.600 255.700 ;
        RECT 20.400 254.300 21.200 254.400 ;
        RECT 7.700 253.700 21.200 254.300 ;
        RECT 7.700 252.400 8.300 253.700 ;
        RECT 20.400 253.600 21.200 253.700 ;
        RECT 25.200 254.300 26.000 254.400 ;
        RECT 36.400 254.300 37.200 254.400 ;
        RECT 25.200 253.700 37.200 254.300 ;
        RECT 25.200 253.600 26.000 253.700 ;
        RECT 36.400 253.600 37.200 253.700 ;
        RECT 42.800 254.300 43.600 254.400 ;
        RECT 54.000 254.300 54.800 254.400 ;
        RECT 42.800 253.700 54.800 254.300 ;
        RECT 42.800 253.600 43.600 253.700 ;
        RECT 54.000 253.600 54.800 253.700 ;
        RECT 70.000 254.300 70.800 254.400 ;
        RECT 74.800 254.300 75.600 254.400 ;
        RECT 70.000 253.700 75.600 254.300 ;
        RECT 70.000 253.600 70.800 253.700 ;
        RECT 74.800 253.600 75.600 253.700 ;
        RECT 158.000 253.600 158.800 254.400 ;
        RECT 161.200 254.300 162.000 254.400 ;
        RECT 223.600 254.300 224.400 254.400 ;
        RECT 161.200 253.700 224.400 254.300 ;
        RECT 161.200 253.600 162.000 253.700 ;
        RECT 223.600 253.600 224.400 253.700 ;
        RECT 226.800 254.300 227.600 254.400 ;
        RECT 234.800 254.300 235.600 254.400 ;
        RECT 226.800 253.700 235.600 254.300 ;
        RECT 226.800 253.600 227.600 253.700 ;
        RECT 234.800 253.600 235.600 253.700 ;
        RECT 322.800 254.300 323.600 254.400 ;
        RECT 329.200 254.300 330.000 254.400 ;
        RECT 322.800 253.700 330.000 254.300 ;
        RECT 322.800 253.600 323.600 253.700 ;
        RECT 329.200 253.600 330.000 253.700 ;
        RECT 334.000 254.300 334.800 254.400 ;
        RECT 338.800 254.300 339.600 254.400 ;
        RECT 334.000 253.700 339.600 254.300 ;
        RECT 334.000 253.600 334.800 253.700 ;
        RECT 338.800 253.600 339.600 253.700 ;
        RECT 430.000 254.300 430.800 254.400 ;
        RECT 431.600 254.300 432.400 254.400 ;
        RECT 434.800 254.300 435.600 254.400 ;
        RECT 430.000 253.700 435.600 254.300 ;
        RECT 430.000 253.600 430.800 253.700 ;
        RECT 431.600 253.600 432.400 253.700 ;
        RECT 434.800 253.600 435.600 253.700 ;
        RECT 476.400 254.300 477.200 254.400 ;
        RECT 492.400 254.300 493.200 254.400 ;
        RECT 476.400 253.700 493.200 254.300 ;
        RECT 476.400 253.600 477.200 253.700 ;
        RECT 492.400 253.600 493.200 253.700 ;
        RECT 4.400 252.300 5.200 252.400 ;
        RECT 7.600 252.300 8.400 252.400 ;
        RECT 4.400 251.700 8.400 252.300 ;
        RECT 4.400 251.600 5.200 251.700 ;
        RECT 7.600 251.600 8.400 251.700 ;
        RECT 12.400 252.300 13.200 252.400 ;
        RECT 14.000 252.300 14.800 252.400 ;
        RECT 15.600 252.300 16.400 252.400 ;
        RECT 12.400 251.700 16.400 252.300 ;
        RECT 12.400 251.600 13.200 251.700 ;
        RECT 14.000 251.600 14.800 251.700 ;
        RECT 15.600 251.600 16.400 251.700 ;
        RECT 23.600 252.300 24.400 252.400 ;
        RECT 26.800 252.300 27.600 252.400 ;
        RECT 31.600 252.300 32.400 252.400 ;
        RECT 23.600 251.700 32.400 252.300 ;
        RECT 23.600 251.600 24.400 251.700 ;
        RECT 26.800 251.600 27.600 251.700 ;
        RECT 31.600 251.600 32.400 251.700 ;
        RECT 34.800 252.300 35.600 252.400 ;
        RECT 49.200 252.300 50.000 252.400 ;
        RECT 34.800 251.700 50.000 252.300 ;
        RECT 34.800 251.600 35.600 251.700 ;
        RECT 49.200 251.600 50.000 251.700 ;
        RECT 63.600 252.300 64.400 252.400 ;
        RECT 66.800 252.300 67.600 252.400 ;
        RECT 63.600 251.700 67.600 252.300 ;
        RECT 63.600 251.600 64.400 251.700 ;
        RECT 66.800 251.600 67.600 251.700 ;
        RECT 70.000 252.300 70.800 252.400 ;
        RECT 100.400 252.300 101.200 252.400 ;
        RECT 70.000 251.700 101.200 252.300 ;
        RECT 70.000 251.600 70.800 251.700 ;
        RECT 100.400 251.600 101.200 251.700 ;
        RECT 121.200 252.300 122.000 252.400 ;
        RECT 169.200 252.300 170.000 252.400 ;
        RECT 121.200 251.700 170.000 252.300 ;
        RECT 121.200 251.600 122.000 251.700 ;
        RECT 169.200 251.600 170.000 251.700 ;
        RECT 329.200 252.300 330.000 252.400 ;
        RECT 345.200 252.300 346.000 252.400 ;
        RECT 329.200 251.700 346.000 252.300 ;
        RECT 329.200 251.600 330.000 251.700 ;
        RECT 345.200 251.600 346.000 251.700 ;
        RECT 418.800 252.300 419.600 252.400 ;
        RECT 442.800 252.300 443.600 252.400 ;
        RECT 418.800 251.700 443.600 252.300 ;
        RECT 418.800 251.600 419.600 251.700 ;
        RECT 442.800 251.600 443.600 251.700 ;
        RECT 471.600 252.300 472.400 252.400 ;
        RECT 510.000 252.300 510.800 252.400 ;
        RECT 511.600 252.300 512.400 252.400 ;
        RECT 471.600 251.700 512.400 252.300 ;
        RECT 471.600 251.600 472.400 251.700 ;
        RECT 510.000 251.600 510.800 251.700 ;
        RECT 511.600 251.600 512.400 251.700 ;
        RECT 50.800 250.300 51.600 250.400 ;
        RECT 52.400 250.300 53.200 250.400 ;
        RECT 50.800 249.700 53.200 250.300 ;
        RECT 50.800 249.600 51.600 249.700 ;
        RECT 52.400 249.600 53.200 249.700 ;
        RECT 58.800 250.300 59.600 250.400 ;
        RECT 62.000 250.300 62.800 250.400 ;
        RECT 68.400 250.300 69.200 250.400 ;
        RECT 58.800 249.700 69.200 250.300 ;
        RECT 58.800 249.600 59.600 249.700 ;
        RECT 62.000 249.600 62.800 249.700 ;
        RECT 68.400 249.600 69.200 249.700 ;
        RECT 122.800 250.300 123.600 250.400 ;
        RECT 150.000 250.300 150.800 250.400 ;
        RECT 122.800 249.700 150.800 250.300 ;
        RECT 122.800 249.600 123.600 249.700 ;
        RECT 150.000 249.600 150.800 249.700 ;
        RECT 276.400 250.300 277.200 250.400 ;
        RECT 282.800 250.300 283.600 250.400 ;
        RECT 276.400 249.700 283.600 250.300 ;
        RECT 276.400 249.600 277.200 249.700 ;
        RECT 282.800 249.600 283.600 249.700 ;
        RECT 318.000 250.300 318.800 250.400 ;
        RECT 354.800 250.300 355.600 250.400 ;
        RECT 318.000 249.700 355.600 250.300 ;
        RECT 318.000 249.600 318.800 249.700 ;
        RECT 354.800 249.600 355.600 249.700 ;
        RECT 422.000 250.300 422.800 250.400 ;
        RECT 468.400 250.300 469.200 250.400 ;
        RECT 422.000 249.700 469.200 250.300 ;
        RECT 422.000 249.600 422.800 249.700 ;
        RECT 468.400 249.600 469.200 249.700 ;
        RECT 470.000 250.300 470.800 250.400 ;
        RECT 474.800 250.300 475.600 250.400 ;
        RECT 470.000 249.700 475.600 250.300 ;
        RECT 470.000 249.600 470.800 249.700 ;
        RECT 474.800 249.600 475.600 249.700 ;
        RECT 10.800 248.300 11.600 248.400 ;
        RECT 38.000 248.300 38.800 248.400 ;
        RECT 10.800 247.700 38.800 248.300 ;
        RECT 10.800 247.600 11.600 247.700 ;
        RECT 38.000 247.600 38.800 247.700 ;
        RECT 46.000 248.300 46.800 248.400 ;
        RECT 65.200 248.300 66.000 248.400 ;
        RECT 46.000 247.700 66.000 248.300 ;
        RECT 46.000 247.600 46.800 247.700 ;
        RECT 65.200 247.600 66.000 247.700 ;
        RECT 110.000 248.300 110.800 248.400 ;
        RECT 114.800 248.300 115.600 248.400 ;
        RECT 134.000 248.300 134.800 248.400 ;
        RECT 140.400 248.300 141.200 248.400 ;
        RECT 158.000 248.300 158.800 248.400 ;
        RECT 182.000 248.300 182.800 248.400 ;
        RECT 110.000 247.700 182.800 248.300 ;
        RECT 110.000 247.600 110.800 247.700 ;
        RECT 114.800 247.600 115.600 247.700 ;
        RECT 134.000 247.600 134.800 247.700 ;
        RECT 140.400 247.600 141.200 247.700 ;
        RECT 158.000 247.600 158.800 247.700 ;
        RECT 182.000 247.600 182.800 247.700 ;
        RECT 345.200 248.300 346.000 248.400 ;
        RECT 346.800 248.300 347.600 248.400 ;
        RECT 345.200 247.700 347.600 248.300 ;
        RECT 345.200 247.600 346.000 247.700 ;
        RECT 346.800 247.600 347.600 247.700 ;
        RECT 18.800 246.300 19.600 246.400 ;
        RECT 20.400 246.300 21.200 246.400 ;
        RECT 18.800 245.700 21.200 246.300 ;
        RECT 18.800 245.600 19.600 245.700 ;
        RECT 20.400 245.600 21.200 245.700 ;
        RECT 30.000 246.300 30.800 246.400 ;
        RECT 39.600 246.300 40.400 246.400 ;
        RECT 30.000 245.700 40.400 246.300 ;
        RECT 30.000 245.600 30.800 245.700 ;
        RECT 39.600 245.600 40.400 245.700 ;
        RECT 41.200 246.300 42.000 246.400 ;
        RECT 47.600 246.300 48.400 246.400 ;
        RECT 41.200 245.700 48.400 246.300 ;
        RECT 41.200 245.600 42.000 245.700 ;
        RECT 47.600 245.600 48.400 245.700 ;
        RECT 57.200 246.300 58.000 246.400 ;
        RECT 58.800 246.300 59.600 246.400 ;
        RECT 62.000 246.300 62.800 246.400 ;
        RECT 76.400 246.300 77.200 246.400 ;
        RECT 57.200 245.700 77.200 246.300 ;
        RECT 57.200 245.600 58.000 245.700 ;
        RECT 58.800 245.600 59.600 245.700 ;
        RECT 62.000 245.600 62.800 245.700 ;
        RECT 76.400 245.600 77.200 245.700 ;
        RECT 135.600 246.300 136.400 246.400 ;
        RECT 146.800 246.300 147.600 246.400 ;
        RECT 135.600 245.700 147.600 246.300 ;
        RECT 135.600 245.600 136.400 245.700 ;
        RECT 146.800 245.600 147.600 245.700 ;
        RECT 431.600 246.300 432.400 246.400 ;
        RECT 450.800 246.300 451.600 246.400 ;
        RECT 431.600 245.700 451.600 246.300 ;
        RECT 431.600 245.600 432.400 245.700 ;
        RECT 450.800 245.600 451.600 245.700 ;
        RECT 418.800 244.300 419.600 244.400 ;
        RECT 478.000 244.300 478.800 244.400 ;
        RECT 482.800 244.300 483.600 244.400 ;
        RECT 516.400 244.300 517.200 244.400 ;
        RECT 530.800 244.300 531.600 244.400 ;
        RECT 418.800 243.700 531.600 244.300 ;
        RECT 418.800 243.600 419.600 243.700 ;
        RECT 478.000 243.600 478.800 243.700 ;
        RECT 482.800 243.600 483.600 243.700 ;
        RECT 516.400 243.600 517.200 243.700 ;
        RECT 530.800 243.600 531.600 243.700 ;
        RECT 543.600 244.300 544.400 244.400 ;
        RECT 548.400 244.300 549.200 244.400 ;
        RECT 543.600 243.700 549.200 244.300 ;
        RECT 543.600 243.600 544.400 243.700 ;
        RECT 548.400 243.600 549.200 243.700 ;
        RECT 46.000 242.300 46.800 242.400 ;
        RECT 49.200 242.300 50.000 242.400 ;
        RECT 46.000 241.700 50.000 242.300 ;
        RECT 46.000 241.600 46.800 241.700 ;
        RECT 49.200 241.600 50.000 241.700 ;
        RECT 151.600 242.300 152.400 242.400 ;
        RECT 154.800 242.300 155.600 242.400 ;
        RECT 151.600 241.700 155.600 242.300 ;
        RECT 151.600 241.600 152.400 241.700 ;
        RECT 154.800 241.600 155.600 241.700 ;
        RECT 212.400 242.300 213.200 242.400 ;
        RECT 241.200 242.300 242.000 242.400 ;
        RECT 212.400 241.700 242.000 242.300 ;
        RECT 212.400 241.600 213.200 241.700 ;
        RECT 241.200 241.600 242.000 241.700 ;
        RECT 257.200 242.300 258.000 242.400 ;
        RECT 263.600 242.300 264.400 242.400 ;
        RECT 257.200 241.700 264.400 242.300 ;
        RECT 257.200 241.600 258.000 241.700 ;
        RECT 263.600 241.600 264.400 241.700 ;
        RECT 266.800 242.300 267.600 242.400 ;
        RECT 356.400 242.300 357.200 242.400 ;
        RECT 266.800 241.700 357.200 242.300 ;
        RECT 266.800 241.600 267.600 241.700 ;
        RECT 356.400 241.600 357.200 241.700 ;
        RECT 433.200 242.300 434.000 242.400 ;
        RECT 441.200 242.300 442.000 242.400 ;
        RECT 433.200 241.700 442.000 242.300 ;
        RECT 433.200 241.600 434.000 241.700 ;
        RECT 441.200 241.600 442.000 241.700 ;
        RECT 49.200 240.300 50.000 240.400 ;
        RECT 73.200 240.300 74.000 240.400 ;
        RECT 103.600 240.300 104.400 240.400 ;
        RECT 49.200 239.700 104.400 240.300 ;
        RECT 49.200 239.600 50.000 239.700 ;
        RECT 73.200 239.600 74.000 239.700 ;
        RECT 103.600 239.600 104.400 239.700 ;
        RECT 308.400 240.300 309.200 240.400 ;
        RECT 359.600 240.300 360.400 240.400 ;
        RECT 308.400 239.700 360.400 240.300 ;
        RECT 308.400 239.600 309.200 239.700 ;
        RECT 359.600 239.600 360.400 239.700 ;
        RECT 438.000 240.300 438.800 240.400 ;
        RECT 441.200 240.300 442.000 240.400 ;
        RECT 438.000 239.700 442.000 240.300 ;
        RECT 438.000 239.600 438.800 239.700 ;
        RECT 441.200 239.600 442.000 239.700 ;
        RECT 39.600 238.300 40.400 238.400 ;
        RECT 70.000 238.300 70.800 238.400 ;
        RECT 74.800 238.300 75.600 238.400 ;
        RECT 39.600 237.700 75.600 238.300 ;
        RECT 39.600 237.600 40.400 237.700 ;
        RECT 70.000 237.600 70.800 237.700 ;
        RECT 74.800 237.600 75.600 237.700 ;
        RECT 102.000 238.300 102.800 238.400 ;
        RECT 206.000 238.300 206.800 238.400 ;
        RECT 102.000 237.700 206.800 238.300 ;
        RECT 102.000 237.600 102.800 237.700 ;
        RECT 206.000 237.600 206.800 237.700 ;
        RECT 302.000 238.300 302.800 238.400 ;
        RECT 305.200 238.300 306.000 238.400 ;
        RECT 302.000 237.700 306.000 238.300 ;
        RECT 302.000 237.600 302.800 237.700 ;
        RECT 305.200 237.600 306.000 237.700 ;
        RECT 420.400 238.300 421.200 238.400 ;
        RECT 444.400 238.300 445.200 238.400 ;
        RECT 420.400 237.700 445.200 238.300 ;
        RECT 420.400 237.600 421.200 237.700 ;
        RECT 444.400 237.600 445.200 237.700 ;
        RECT 455.600 238.300 456.400 238.400 ;
        RECT 458.800 238.300 459.600 238.400 ;
        RECT 455.600 237.700 459.600 238.300 ;
        RECT 455.600 237.600 456.400 237.700 ;
        RECT 458.800 237.600 459.600 237.700 ;
        RECT 38.000 236.300 38.800 236.400 ;
        RECT 50.800 236.300 51.600 236.400 ;
        RECT 38.000 235.700 51.600 236.300 ;
        RECT 38.000 235.600 38.800 235.700 ;
        RECT 50.800 235.600 51.600 235.700 ;
        RECT 52.400 236.300 53.200 236.400 ;
        RECT 100.400 236.300 101.200 236.400 ;
        RECT 52.400 235.700 101.200 236.300 ;
        RECT 52.400 235.600 53.200 235.700 ;
        RECT 100.400 235.600 101.200 235.700 ;
        RECT 183.600 236.300 184.400 236.400 ;
        RECT 330.800 236.300 331.600 236.400 ;
        RECT 351.600 236.300 352.400 236.400 ;
        RECT 183.600 235.700 352.400 236.300 ;
        RECT 183.600 235.600 184.400 235.700 ;
        RECT 330.800 235.600 331.600 235.700 ;
        RECT 351.600 235.600 352.400 235.700 ;
        RECT 361.200 236.300 362.000 236.400 ;
        RECT 366.000 236.300 366.800 236.400 ;
        RECT 361.200 235.700 366.800 236.300 ;
        RECT 361.200 235.600 362.000 235.700 ;
        RECT 366.000 235.600 366.800 235.700 ;
        RECT 38.000 234.300 38.800 234.400 ;
        RECT 60.400 234.300 61.200 234.400 ;
        RECT 68.400 234.300 69.200 234.400 ;
        RECT 73.200 234.300 74.000 234.400 ;
        RECT 38.000 233.700 74.000 234.300 ;
        RECT 38.000 233.600 38.800 233.700 ;
        RECT 60.400 233.600 61.200 233.700 ;
        RECT 68.400 233.600 69.200 233.700 ;
        RECT 73.200 233.600 74.000 233.700 ;
        RECT 78.000 234.300 78.800 234.400 ;
        RECT 84.400 234.300 85.200 234.400 ;
        RECT 87.600 234.300 88.400 234.400 ;
        RECT 78.000 233.700 88.400 234.300 ;
        RECT 78.000 233.600 78.800 233.700 ;
        RECT 84.400 233.600 85.200 233.700 ;
        RECT 87.600 233.600 88.400 233.700 ;
        RECT 150.000 234.300 150.800 234.400 ;
        RECT 161.200 234.300 162.000 234.400 ;
        RECT 150.000 233.700 162.000 234.300 ;
        RECT 150.000 233.600 150.800 233.700 ;
        RECT 161.200 233.600 162.000 233.700 ;
        RECT 177.200 234.300 178.000 234.400 ;
        RECT 180.400 234.300 181.200 234.400 ;
        RECT 188.400 234.300 189.200 234.400 ;
        RECT 194.800 234.300 195.600 234.400 ;
        RECT 249.200 234.300 250.000 234.400 ;
        RECT 177.200 233.700 250.000 234.300 ;
        RECT 177.200 233.600 178.000 233.700 ;
        RECT 180.400 233.600 181.200 233.700 ;
        RECT 188.400 233.600 189.200 233.700 ;
        RECT 194.800 233.600 195.600 233.700 ;
        RECT 249.200 233.600 250.000 233.700 ;
        RECT 431.600 234.300 432.400 234.400 ;
        RECT 439.600 234.300 440.400 234.400 ;
        RECT 460.400 234.300 461.200 234.400 ;
        RECT 466.800 234.300 467.600 234.400 ;
        RECT 431.600 233.700 467.600 234.300 ;
        RECT 431.600 233.600 432.400 233.700 ;
        RECT 439.600 233.600 440.400 233.700 ;
        RECT 460.400 233.600 461.200 233.700 ;
        RECT 466.800 233.600 467.600 233.700 ;
        RECT 22.000 232.300 22.800 232.400 ;
        RECT 44.400 232.300 45.200 232.400 ;
        RECT 22.000 231.700 45.200 232.300 ;
        RECT 22.000 231.600 22.800 231.700 ;
        RECT 44.400 231.600 45.200 231.700 ;
        RECT 71.600 232.300 72.400 232.400 ;
        RECT 82.800 232.300 83.600 232.400 ;
        RECT 71.600 231.700 83.600 232.300 ;
        RECT 71.600 231.600 72.400 231.700 ;
        RECT 82.800 231.600 83.600 231.700 ;
        RECT 145.200 232.300 146.000 232.400 ;
        RECT 153.200 232.300 154.000 232.400 ;
        RECT 145.200 231.700 154.000 232.300 ;
        RECT 145.200 231.600 146.000 231.700 ;
        RECT 153.200 231.600 154.000 231.700 ;
        RECT 158.000 232.300 158.800 232.400 ;
        RECT 162.800 232.300 163.600 232.400 ;
        RECT 158.000 231.700 163.600 232.300 ;
        RECT 158.000 231.600 158.800 231.700 ;
        RECT 162.800 231.600 163.600 231.700 ;
        RECT 166.000 232.300 166.800 232.400 ;
        RECT 167.600 232.300 168.400 232.400 ;
        RECT 170.800 232.300 171.600 232.400 ;
        RECT 166.000 231.700 171.600 232.300 ;
        RECT 166.000 231.600 166.800 231.700 ;
        RECT 167.600 231.600 168.400 231.700 ;
        RECT 170.800 231.600 171.600 231.700 ;
        RECT 177.200 232.300 178.000 232.400 ;
        RECT 178.800 232.300 179.600 232.400 ;
        RECT 191.600 232.300 192.400 232.400 ;
        RECT 177.200 231.700 192.400 232.300 ;
        RECT 177.200 231.600 178.000 231.700 ;
        RECT 178.800 231.600 179.600 231.700 ;
        RECT 191.600 231.600 192.400 231.700 ;
        RECT 202.800 232.300 203.600 232.400 ;
        RECT 209.200 232.300 210.000 232.400 ;
        RECT 202.800 231.700 210.000 232.300 ;
        RECT 202.800 231.600 203.600 231.700 ;
        RECT 209.200 231.600 210.000 231.700 ;
        RECT 276.400 232.300 277.200 232.400 ;
        RECT 311.600 232.300 312.400 232.400 ;
        RECT 276.400 231.700 312.400 232.300 ;
        RECT 276.400 231.600 277.200 231.700 ;
        RECT 311.600 231.600 312.400 231.700 ;
        RECT 330.800 232.300 331.600 232.400 ;
        RECT 337.200 232.300 338.000 232.400 ;
        RECT 330.800 231.700 338.000 232.300 ;
        RECT 330.800 231.600 331.600 231.700 ;
        RECT 337.200 231.600 338.000 231.700 ;
        RECT 359.600 232.300 360.400 232.400 ;
        RECT 367.600 232.300 368.400 232.400 ;
        RECT 359.600 231.700 368.400 232.300 ;
        RECT 359.600 231.600 360.400 231.700 ;
        RECT 367.600 231.600 368.400 231.700 ;
        RECT 370.800 232.300 371.600 232.400 ;
        RECT 415.600 232.300 416.400 232.400 ;
        RECT 418.800 232.300 419.600 232.400 ;
        RECT 370.800 231.700 419.600 232.300 ;
        RECT 370.800 231.600 371.600 231.700 ;
        RECT 415.600 231.600 416.400 231.700 ;
        RECT 418.800 231.600 419.600 231.700 ;
        RECT 428.400 232.300 429.200 232.400 ;
        RECT 441.200 232.300 442.000 232.400 ;
        RECT 446.000 232.300 446.800 232.400 ;
        RECT 457.200 232.300 458.000 232.400 ;
        RECT 463.600 232.300 464.400 232.400 ;
        RECT 428.400 231.700 464.400 232.300 ;
        RECT 428.400 231.600 429.200 231.700 ;
        RECT 441.200 231.600 442.000 231.700 ;
        RECT 446.000 231.600 446.800 231.700 ;
        RECT 457.200 231.600 458.000 231.700 ;
        RECT 463.600 231.600 464.400 231.700 ;
        RECT 465.200 232.300 466.000 232.400 ;
        RECT 476.400 232.300 477.200 232.400 ;
        RECT 465.200 231.700 477.200 232.300 ;
        RECT 465.200 231.600 466.000 231.700 ;
        RECT 476.400 231.600 477.200 231.700 ;
        RECT 478.000 232.300 478.800 232.400 ;
        RECT 487.600 232.300 488.400 232.400 ;
        RECT 478.000 231.700 488.400 232.300 ;
        RECT 478.000 231.600 478.800 231.700 ;
        RECT 487.600 231.600 488.400 231.700 ;
        RECT 4.400 230.300 5.200 230.400 ;
        RECT 36.400 230.300 37.200 230.400 ;
        RECT 4.400 229.700 37.200 230.300 ;
        RECT 4.400 229.600 5.200 229.700 ;
        RECT 36.400 229.600 37.200 229.700 ;
        RECT 46.000 230.300 46.800 230.400 ;
        RECT 47.600 230.300 48.400 230.400 ;
        RECT 46.000 229.700 48.400 230.300 ;
        RECT 46.000 229.600 46.800 229.700 ;
        RECT 47.600 229.600 48.400 229.700 ;
        RECT 60.400 230.300 61.200 230.400 ;
        RECT 65.200 230.300 66.000 230.400 ;
        RECT 60.400 229.700 66.000 230.300 ;
        RECT 60.400 229.600 61.200 229.700 ;
        RECT 65.200 229.600 66.000 229.700 ;
        RECT 79.600 230.300 80.400 230.400 ;
        RECT 86.000 230.300 86.800 230.400 ;
        RECT 92.400 230.300 93.200 230.400 ;
        RECT 105.200 230.300 106.000 230.400 ;
        RECT 79.600 229.700 106.000 230.300 ;
        RECT 79.600 229.600 80.400 229.700 ;
        RECT 86.000 229.600 86.800 229.700 ;
        RECT 92.400 229.600 93.200 229.700 ;
        RECT 105.200 229.600 106.000 229.700 ;
        RECT 159.600 230.300 160.400 230.400 ;
        RECT 169.200 230.300 170.000 230.400 ;
        RECT 159.600 229.700 170.000 230.300 ;
        RECT 159.600 229.600 160.400 229.700 ;
        RECT 169.200 229.600 170.000 229.700 ;
        RECT 191.600 230.300 192.400 230.400 ;
        RECT 199.600 230.300 200.400 230.400 ;
        RECT 191.600 229.700 200.400 230.300 ;
        RECT 191.600 229.600 192.400 229.700 ;
        RECT 199.600 229.600 200.400 229.700 ;
        RECT 234.800 230.300 235.600 230.400 ;
        RECT 249.200 230.300 250.000 230.400 ;
        RECT 234.800 229.700 250.000 230.300 ;
        RECT 234.800 229.600 235.600 229.700 ;
        RECT 249.200 229.600 250.000 229.700 ;
        RECT 270.000 230.300 270.800 230.400 ;
        RECT 276.400 230.300 277.200 230.400 ;
        RECT 270.000 229.700 277.200 230.300 ;
        RECT 270.000 229.600 270.800 229.700 ;
        RECT 276.400 229.600 277.200 229.700 ;
        RECT 321.200 230.300 322.000 230.400 ;
        RECT 327.600 230.300 328.400 230.400 ;
        RECT 332.400 230.300 333.200 230.400 ;
        RECT 338.800 230.300 339.600 230.400 ;
        RECT 356.400 230.300 357.200 230.400 ;
        RECT 366.000 230.300 366.800 230.400 ;
        RECT 321.200 229.700 366.800 230.300 ;
        RECT 321.200 229.600 322.000 229.700 ;
        RECT 327.600 229.600 328.400 229.700 ;
        RECT 332.400 229.600 333.200 229.700 ;
        RECT 338.800 229.600 339.600 229.700 ;
        RECT 356.400 229.600 357.200 229.700 ;
        RECT 366.000 229.600 366.800 229.700 ;
        RECT 377.200 230.300 378.000 230.400 ;
        RECT 430.000 230.300 430.800 230.400 ;
        RECT 436.400 230.300 437.200 230.400 ;
        RECT 377.200 229.700 429.100 230.300 ;
        RECT 377.200 229.600 378.000 229.700 ;
        RECT 18.800 228.300 19.600 228.400 ;
        RECT 39.600 228.300 40.400 228.400 ;
        RECT 50.800 228.300 51.600 228.400 ;
        RECT 18.800 227.700 22.700 228.300 ;
        RECT 18.800 227.600 19.600 227.700 ;
        RECT 22.100 226.400 22.700 227.700 ;
        RECT 39.600 227.700 51.600 228.300 ;
        RECT 39.600 227.600 40.400 227.700 ;
        RECT 50.800 227.600 51.600 227.700 ;
        RECT 62.000 228.300 62.800 228.400 ;
        RECT 102.000 228.300 102.800 228.400 ;
        RECT 62.000 227.700 102.800 228.300 ;
        RECT 62.000 227.600 62.800 227.700 ;
        RECT 102.000 227.600 102.800 227.700 ;
        RECT 132.400 228.300 133.200 228.400 ;
        RECT 138.800 228.300 139.600 228.400 ;
        RECT 158.000 228.300 158.800 228.400 ;
        RECT 166.000 228.300 166.800 228.400 ;
        RECT 174.000 228.300 174.800 228.400 ;
        RECT 198.000 228.300 198.800 228.400 ;
        RECT 212.400 228.300 213.200 228.400 ;
        RECT 132.400 227.700 213.200 228.300 ;
        RECT 132.400 227.600 133.200 227.700 ;
        RECT 138.800 227.600 139.600 227.700 ;
        RECT 158.000 227.600 158.800 227.700 ;
        RECT 166.000 227.600 166.800 227.700 ;
        RECT 174.000 227.600 174.800 227.700 ;
        RECT 198.000 227.600 198.800 227.700 ;
        RECT 212.400 227.600 213.200 227.700 ;
        RECT 260.400 227.600 261.200 228.400 ;
        RECT 282.800 228.300 283.600 228.400 ;
        RECT 319.600 228.300 320.400 228.400 ;
        RECT 322.800 228.300 323.600 228.400 ;
        RECT 282.800 227.700 323.600 228.300 ;
        RECT 282.800 227.600 283.600 227.700 ;
        RECT 319.600 227.600 320.400 227.700 ;
        RECT 322.800 227.600 323.600 227.700 ;
        RECT 324.400 228.300 325.200 228.400 ;
        RECT 332.400 228.300 333.200 228.400 ;
        RECT 324.400 227.700 333.200 228.300 ;
        RECT 324.400 227.600 325.200 227.700 ;
        RECT 332.400 227.600 333.200 227.700 ;
        RECT 334.000 228.300 334.800 228.400 ;
        RECT 337.200 228.300 338.000 228.400 ;
        RECT 343.600 228.300 344.400 228.400 ;
        RECT 334.000 227.700 344.400 228.300 ;
        RECT 334.000 227.600 334.800 227.700 ;
        RECT 337.200 227.600 338.000 227.700 ;
        RECT 343.600 227.600 344.400 227.700 ;
        RECT 353.200 228.300 354.000 228.400 ;
        RECT 370.800 228.300 371.600 228.400 ;
        RECT 353.200 227.700 371.600 228.300 ;
        RECT 353.200 227.600 354.000 227.700 ;
        RECT 370.800 227.600 371.600 227.700 ;
        RECT 398.000 228.300 398.800 228.400 ;
        RECT 418.800 228.300 419.600 228.400 ;
        RECT 398.000 227.700 419.600 228.300 ;
        RECT 428.500 228.300 429.100 229.700 ;
        RECT 430.000 229.700 437.200 230.300 ;
        RECT 430.000 229.600 430.800 229.700 ;
        RECT 436.400 229.600 437.200 229.700 ;
        RECT 455.600 230.300 456.400 230.400 ;
        RECT 479.600 230.300 480.400 230.400 ;
        RECT 455.600 229.700 480.400 230.300 ;
        RECT 455.600 229.600 456.400 229.700 ;
        RECT 479.600 229.600 480.400 229.700 ;
        RECT 484.400 230.300 485.200 230.400 ;
        RECT 516.400 230.300 517.200 230.400 ;
        RECT 484.400 229.700 517.200 230.300 ;
        RECT 484.400 229.600 485.200 229.700 ;
        RECT 516.400 229.600 517.200 229.700 ;
        RECT 431.600 228.300 432.400 228.400 ;
        RECT 434.800 228.300 435.600 228.400 ;
        RECT 428.500 227.700 435.600 228.300 ;
        RECT 398.000 227.600 398.800 227.700 ;
        RECT 418.800 227.600 419.600 227.700 ;
        RECT 431.600 227.600 432.400 227.700 ;
        RECT 434.800 227.600 435.600 227.700 ;
        RECT 450.800 228.300 451.600 228.400 ;
        RECT 450.800 227.700 457.900 228.300 ;
        RECT 450.800 227.600 451.600 227.700 ;
        RECT 18.800 226.300 19.600 226.400 ;
        RECT 20.400 226.300 21.200 226.400 ;
        RECT 18.800 225.700 21.200 226.300 ;
        RECT 18.800 225.600 19.600 225.700 ;
        RECT 20.400 225.600 21.200 225.700 ;
        RECT 22.000 225.600 22.800 226.400 ;
        RECT 33.200 226.300 34.000 226.400 ;
        RECT 39.700 226.300 40.300 227.600 ;
        RECT 457.300 226.400 457.900 227.700 ;
        RECT 458.800 227.600 459.600 228.400 ;
        RECT 460.400 228.300 461.200 228.400 ;
        RECT 470.000 228.300 470.800 228.400 ;
        RECT 460.400 227.700 470.800 228.300 ;
        RECT 460.400 227.600 461.200 227.700 ;
        RECT 470.000 227.600 470.800 227.700 ;
        RECT 471.600 228.300 472.400 228.400 ;
        RECT 473.200 228.300 474.000 228.400 ;
        RECT 471.600 227.700 474.000 228.300 ;
        RECT 471.600 227.600 472.400 227.700 ;
        RECT 473.200 227.600 474.000 227.700 ;
        RECT 474.800 228.300 475.600 228.400 ;
        RECT 497.200 228.300 498.000 228.400 ;
        RECT 474.800 227.700 498.000 228.300 ;
        RECT 474.800 227.600 475.600 227.700 ;
        RECT 497.200 227.600 498.000 227.700 ;
        RECT 33.200 225.700 40.300 226.300 ;
        RECT 54.000 226.300 54.800 226.400 ;
        RECT 62.000 226.300 62.800 226.400 ;
        RECT 54.000 225.700 62.800 226.300 ;
        RECT 33.200 225.600 34.000 225.700 ;
        RECT 54.000 225.600 54.800 225.700 ;
        RECT 62.000 225.600 62.800 225.700 ;
        RECT 145.200 226.300 146.000 226.400 ;
        RECT 178.800 226.300 179.600 226.400 ;
        RECT 145.200 225.700 179.600 226.300 ;
        RECT 145.200 225.600 146.000 225.700 ;
        RECT 178.800 225.600 179.600 225.700 ;
        RECT 204.400 226.300 205.200 226.400 ;
        RECT 225.200 226.300 226.000 226.400 ;
        RECT 204.400 225.700 226.000 226.300 ;
        RECT 204.400 225.600 205.200 225.700 ;
        RECT 225.200 225.600 226.000 225.700 ;
        RECT 244.400 226.300 245.200 226.400 ;
        RECT 276.400 226.300 277.200 226.400 ;
        RECT 244.400 225.700 277.200 226.300 ;
        RECT 244.400 225.600 245.200 225.700 ;
        RECT 276.400 225.600 277.200 225.700 ;
        RECT 305.200 226.300 306.000 226.400 ;
        RECT 329.200 226.300 330.000 226.400 ;
        RECT 305.200 225.700 330.000 226.300 ;
        RECT 305.200 225.600 306.000 225.700 ;
        RECT 329.200 225.600 330.000 225.700 ;
        RECT 378.800 226.300 379.600 226.400 ;
        RECT 412.400 226.300 413.200 226.400 ;
        RECT 378.800 225.700 413.200 226.300 ;
        RECT 378.800 225.600 379.600 225.700 ;
        RECT 412.400 225.600 413.200 225.700 ;
        RECT 417.200 226.300 418.000 226.400 ;
        RECT 433.200 226.300 434.000 226.400 ;
        RECT 417.200 225.700 434.000 226.300 ;
        RECT 417.200 225.600 418.000 225.700 ;
        RECT 433.200 225.600 434.000 225.700 ;
        RECT 457.200 226.300 458.000 226.400 ;
        RECT 479.600 226.300 480.400 226.400 ;
        RECT 457.200 225.700 480.400 226.300 ;
        RECT 457.200 225.600 458.000 225.700 ;
        RECT 479.600 225.600 480.400 225.700 ;
        RECT 495.600 226.300 496.400 226.400 ;
        RECT 513.200 226.300 514.000 226.400 ;
        RECT 495.600 225.700 514.000 226.300 ;
        RECT 495.600 225.600 496.400 225.700 ;
        RECT 513.200 225.600 514.000 225.700 ;
        RECT 522.800 226.300 523.600 226.400 ;
        RECT 526.000 226.300 526.800 226.400 ;
        RECT 522.800 225.700 526.800 226.300 ;
        RECT 522.800 225.600 523.600 225.700 ;
        RECT 526.000 225.600 526.800 225.700 ;
        RECT 537.200 226.300 538.000 226.400 ;
        RECT 542.000 226.300 542.800 226.400 ;
        RECT 546.800 226.300 547.600 226.400 ;
        RECT 537.200 225.700 547.600 226.300 ;
        RECT 537.200 225.600 538.000 225.700 ;
        RECT 542.000 225.600 542.800 225.700 ;
        RECT 546.800 225.600 547.600 225.700 ;
        RECT 30.000 224.300 30.800 224.400 ;
        RECT 79.600 224.300 80.400 224.400 ;
        RECT 30.000 223.700 80.400 224.300 ;
        RECT 30.000 223.600 30.800 223.700 ;
        RECT 79.600 223.600 80.400 223.700 ;
        RECT 86.000 224.300 86.800 224.400 ;
        RECT 97.200 224.300 98.000 224.400 ;
        RECT 86.000 223.700 98.000 224.300 ;
        RECT 86.000 223.600 86.800 223.700 ;
        RECT 97.200 223.600 98.000 223.700 ;
        RECT 113.200 224.300 114.000 224.400 ;
        RECT 124.400 224.300 125.200 224.400 ;
        RECT 113.200 223.700 125.200 224.300 ;
        RECT 113.200 223.600 114.000 223.700 ;
        RECT 124.400 223.600 125.200 223.700 ;
        RECT 164.400 224.300 165.200 224.400 ;
        RECT 169.200 224.300 170.000 224.400 ;
        RECT 172.400 224.300 173.200 224.400 ;
        RECT 164.400 223.700 173.200 224.300 ;
        RECT 164.400 223.600 165.200 223.700 ;
        RECT 169.200 223.600 170.000 223.700 ;
        RECT 172.400 223.600 173.200 223.700 ;
        RECT 175.600 224.300 176.400 224.400 ;
        RECT 186.800 224.300 187.600 224.400 ;
        RECT 175.600 223.700 187.600 224.300 ;
        RECT 175.600 223.600 176.400 223.700 ;
        RECT 186.800 223.600 187.600 223.700 ;
        RECT 374.000 224.300 374.800 224.400 ;
        RECT 378.800 224.300 379.600 224.400 ;
        RECT 374.000 223.700 379.600 224.300 ;
        RECT 374.000 223.600 374.800 223.700 ;
        RECT 378.800 223.600 379.600 223.700 ;
        RECT 385.200 224.300 386.000 224.400 ;
        RECT 410.800 224.300 411.600 224.400 ;
        RECT 385.200 223.700 411.600 224.300 ;
        RECT 385.200 223.600 386.000 223.700 ;
        RECT 410.800 223.600 411.600 223.700 ;
        RECT 412.400 224.300 413.200 224.400 ;
        RECT 423.600 224.300 424.400 224.400 ;
        RECT 438.000 224.300 438.800 224.400 ;
        RECT 470.000 224.300 470.800 224.400 ;
        RECT 473.200 224.300 474.000 224.400 ;
        RECT 474.800 224.300 475.600 224.400 ;
        RECT 537.200 224.300 538.000 224.400 ;
        RECT 412.400 223.700 538.000 224.300 ;
        RECT 412.400 223.600 413.200 223.700 ;
        RECT 423.600 223.600 424.400 223.700 ;
        RECT 438.000 223.600 438.800 223.700 ;
        RECT 470.000 223.600 470.800 223.700 ;
        RECT 473.200 223.600 474.000 223.700 ;
        RECT 474.800 223.600 475.600 223.700 ;
        RECT 537.200 223.600 538.000 223.700 ;
        RECT 6.000 222.300 6.800 222.400 ;
        RECT 42.800 222.300 43.600 222.400 ;
        RECT 6.000 221.700 43.600 222.300 ;
        RECT 6.000 221.600 6.800 221.700 ;
        RECT 42.800 221.600 43.600 221.700 ;
        RECT 159.600 222.300 160.400 222.400 ;
        RECT 162.800 222.300 163.600 222.400 ;
        RECT 178.800 222.300 179.600 222.400 ;
        RECT 185.200 222.300 186.000 222.400 ;
        RECT 159.600 221.700 186.000 222.300 ;
        RECT 159.600 221.600 160.400 221.700 ;
        RECT 162.800 221.600 163.600 221.700 ;
        RECT 178.800 221.600 179.600 221.700 ;
        RECT 185.200 221.600 186.000 221.700 ;
        RECT 196.400 222.300 197.200 222.400 ;
        RECT 220.400 222.300 221.200 222.400 ;
        RECT 196.400 221.700 221.200 222.300 ;
        RECT 196.400 221.600 197.200 221.700 ;
        RECT 220.400 221.600 221.200 221.700 ;
        RECT 284.400 222.300 285.200 222.400 ;
        RECT 302.000 222.300 302.800 222.400 ;
        RECT 308.400 222.300 309.200 222.400 ;
        RECT 319.600 222.300 320.400 222.400 ;
        RECT 284.400 221.700 320.400 222.300 ;
        RECT 284.400 221.600 285.200 221.700 ;
        RECT 302.000 221.600 302.800 221.700 ;
        RECT 308.400 221.600 309.200 221.700 ;
        RECT 319.600 221.600 320.400 221.700 ;
        RECT 322.800 222.300 323.600 222.400 ;
        RECT 390.000 222.300 390.800 222.400 ;
        RECT 322.800 221.700 390.800 222.300 ;
        RECT 322.800 221.600 323.600 221.700 ;
        RECT 390.000 221.600 390.800 221.700 ;
        RECT 402.800 222.300 403.600 222.400 ;
        RECT 414.000 222.300 414.800 222.400 ;
        RECT 402.800 221.700 414.800 222.300 ;
        RECT 402.800 221.600 403.600 221.700 ;
        RECT 414.000 221.600 414.800 221.700 ;
        RECT 433.200 222.300 434.000 222.400 ;
        RECT 452.400 222.300 453.200 222.400 ;
        RECT 433.200 221.700 453.200 222.300 ;
        RECT 433.200 221.600 434.000 221.700 ;
        RECT 452.400 221.600 453.200 221.700 ;
        RECT 458.800 222.300 459.600 222.400 ;
        RECT 490.800 222.300 491.600 222.400 ;
        RECT 458.800 221.700 491.600 222.300 ;
        RECT 458.800 221.600 459.600 221.700 ;
        RECT 490.800 221.600 491.600 221.700 ;
        RECT 508.400 222.300 509.200 222.400 ;
        RECT 522.800 222.300 523.600 222.400 ;
        RECT 508.400 221.700 523.600 222.300 ;
        RECT 508.400 221.600 509.200 221.700 ;
        RECT 522.800 221.600 523.600 221.700 ;
        RECT 22.000 220.300 22.800 220.400 ;
        RECT 28.400 220.300 29.200 220.400 ;
        RECT 31.600 220.300 32.400 220.400 ;
        RECT 55.600 220.300 56.400 220.400 ;
        RECT 22.000 219.700 56.400 220.300 ;
        RECT 22.000 219.600 22.800 219.700 ;
        RECT 28.400 219.600 29.200 219.700 ;
        RECT 31.600 219.600 32.400 219.700 ;
        RECT 55.600 219.600 56.400 219.700 ;
        RECT 146.800 220.300 147.600 220.400 ;
        RECT 167.600 220.300 168.400 220.400 ;
        RECT 199.600 220.300 200.400 220.400 ;
        RECT 146.800 219.700 200.400 220.300 ;
        RECT 146.800 219.600 147.600 219.700 ;
        RECT 167.600 219.600 168.400 219.700 ;
        RECT 199.600 219.600 200.400 219.700 ;
        RECT 226.800 220.300 227.600 220.400 ;
        RECT 238.000 220.300 238.800 220.400 ;
        RECT 226.800 219.700 238.800 220.300 ;
        RECT 226.800 219.600 227.600 219.700 ;
        RECT 238.000 219.600 238.800 219.700 ;
        RECT 257.200 220.300 258.000 220.400 ;
        RECT 263.600 220.300 264.400 220.400 ;
        RECT 257.200 219.700 264.400 220.300 ;
        RECT 257.200 219.600 258.000 219.700 ;
        RECT 263.600 219.600 264.400 219.700 ;
        RECT 289.200 220.300 290.000 220.400 ;
        RECT 326.000 220.300 326.800 220.400 ;
        RECT 337.200 220.300 338.000 220.400 ;
        RECT 532.400 220.300 533.200 220.400 ;
        RECT 289.200 219.700 338.000 220.300 ;
        RECT 289.200 219.600 290.000 219.700 ;
        RECT 326.000 219.600 326.800 219.700 ;
        RECT 337.200 219.600 338.000 219.700 ;
        RECT 495.700 219.700 533.200 220.300 ;
        RECT 15.600 218.300 16.400 218.400 ;
        RECT 65.200 218.300 66.000 218.400 ;
        RECT 68.400 218.300 69.200 218.400 ;
        RECT 15.600 217.700 69.200 218.300 ;
        RECT 15.600 217.600 16.400 217.700 ;
        RECT 65.200 217.600 66.000 217.700 ;
        RECT 68.400 217.600 69.200 217.700 ;
        RECT 78.000 218.300 78.800 218.400 ;
        RECT 95.600 218.300 96.400 218.400 ;
        RECT 78.000 217.700 96.400 218.300 ;
        RECT 78.000 217.600 78.800 217.700 ;
        RECT 95.600 217.600 96.400 217.700 ;
        RECT 135.600 218.300 136.400 218.400 ;
        RECT 250.800 218.300 251.600 218.400 ;
        RECT 135.600 217.700 251.600 218.300 ;
        RECT 135.600 217.600 136.400 217.700 ;
        RECT 250.800 217.600 251.600 217.700 ;
        RECT 255.600 218.300 256.400 218.400 ;
        RECT 342.000 218.300 342.800 218.400 ;
        RECT 255.600 217.700 342.800 218.300 ;
        RECT 255.600 217.600 256.400 217.700 ;
        RECT 342.000 217.600 342.800 217.700 ;
        RECT 343.600 218.300 344.400 218.400 ;
        RECT 354.800 218.300 355.600 218.400 ;
        RECT 370.800 218.300 371.600 218.400 ;
        RECT 343.600 217.700 371.600 218.300 ;
        RECT 343.600 217.600 344.400 217.700 ;
        RECT 354.800 217.600 355.600 217.700 ;
        RECT 370.800 217.600 371.600 217.700 ;
        RECT 375.600 218.300 376.400 218.400 ;
        RECT 388.400 218.300 389.200 218.400 ;
        RECT 375.600 217.700 389.200 218.300 ;
        RECT 375.600 217.600 376.400 217.700 ;
        RECT 388.400 217.600 389.200 217.700 ;
        RECT 399.600 218.300 400.400 218.400 ;
        RECT 412.400 218.300 413.200 218.400 ;
        RECT 399.600 217.700 413.200 218.300 ;
        RECT 399.600 217.600 400.400 217.700 ;
        RECT 412.400 217.600 413.200 217.700 ;
        RECT 434.800 218.300 435.600 218.400 ;
        RECT 449.200 218.300 450.000 218.400 ;
        RECT 495.700 218.300 496.300 219.700 ;
        RECT 532.400 219.600 533.200 219.700 ;
        RECT 434.800 217.700 496.300 218.300 ;
        RECT 500.400 218.300 501.200 218.400 ;
        RECT 514.800 218.300 515.600 218.400 ;
        RECT 500.400 217.700 515.600 218.300 ;
        RECT 434.800 217.600 435.600 217.700 ;
        RECT 449.200 217.600 450.000 217.700 ;
        RECT 500.400 217.600 501.200 217.700 ;
        RECT 514.800 217.600 515.600 217.700 ;
        RECT 7.600 216.300 8.400 216.400 ;
        RECT 17.200 216.300 18.000 216.400 ;
        RECT 26.800 216.300 27.600 216.400 ;
        RECT 7.600 215.700 27.600 216.300 ;
        RECT 7.600 215.600 8.400 215.700 ;
        RECT 17.200 215.600 18.000 215.700 ;
        RECT 26.800 215.600 27.600 215.700 ;
        RECT 30.000 216.300 30.800 216.400 ;
        RECT 38.000 216.300 38.800 216.400 ;
        RECT 30.000 215.700 38.800 216.300 ;
        RECT 30.000 215.600 30.800 215.700 ;
        RECT 38.000 215.600 38.800 215.700 ;
        RECT 183.600 216.300 184.400 216.400 ;
        RECT 194.800 216.300 195.600 216.400 ;
        RECT 183.600 215.700 195.600 216.300 ;
        RECT 183.600 215.600 184.400 215.700 ;
        RECT 194.800 215.600 195.600 215.700 ;
        RECT 201.200 216.300 202.000 216.400 ;
        RECT 222.000 216.300 222.800 216.400 ;
        RECT 201.200 215.700 222.800 216.300 ;
        RECT 201.200 215.600 202.000 215.700 ;
        RECT 222.000 215.600 222.800 215.700 ;
        RECT 223.600 216.300 224.400 216.400 ;
        RECT 233.200 216.300 234.000 216.400 ;
        RECT 223.600 215.700 234.000 216.300 ;
        RECT 223.600 215.600 224.400 215.700 ;
        RECT 233.200 215.600 234.000 215.700 ;
        RECT 292.400 216.300 293.200 216.400 ;
        RECT 326.000 216.300 326.800 216.400 ;
        RECT 334.000 216.300 334.800 216.400 ;
        RECT 292.400 215.700 334.800 216.300 ;
        RECT 292.400 215.600 293.200 215.700 ;
        RECT 326.000 215.600 326.800 215.700 ;
        RECT 334.000 215.600 334.800 215.700 ;
        RECT 337.200 216.300 338.000 216.400 ;
        RECT 396.400 216.300 397.200 216.400 ;
        RECT 407.600 216.300 408.400 216.400 ;
        RECT 337.200 215.700 397.200 216.300 ;
        RECT 337.200 215.600 338.000 215.700 ;
        RECT 396.400 215.600 397.200 215.700 ;
        RECT 399.700 215.700 408.400 216.300 ;
        RECT 9.200 214.300 10.000 214.400 ;
        RECT 15.600 214.300 16.400 214.400 ;
        RECT 18.800 214.300 19.600 214.400 ;
        RECT 9.200 213.700 19.600 214.300 ;
        RECT 9.200 213.600 10.000 213.700 ;
        RECT 15.600 213.600 16.400 213.700 ;
        RECT 18.800 213.600 19.600 213.700 ;
        RECT 36.400 214.300 37.200 214.400 ;
        RECT 39.600 214.300 40.400 214.400 ;
        RECT 36.400 213.700 40.400 214.300 ;
        RECT 36.400 213.600 37.200 213.700 ;
        RECT 39.600 213.600 40.400 213.700 ;
        RECT 63.600 214.300 64.400 214.400 ;
        RECT 89.200 214.300 90.000 214.400 ;
        RECT 63.600 213.700 90.000 214.300 ;
        RECT 63.600 213.600 64.400 213.700 ;
        RECT 89.200 213.600 90.000 213.700 ;
        RECT 92.400 214.300 93.200 214.400 ;
        RECT 97.200 214.300 98.000 214.400 ;
        RECT 92.400 213.700 98.000 214.300 ;
        RECT 92.400 213.600 93.200 213.700 ;
        RECT 97.200 213.600 98.000 213.700 ;
        RECT 129.200 214.300 130.000 214.400 ;
        RECT 158.000 214.300 158.800 214.400 ;
        RECT 129.200 213.700 158.800 214.300 ;
        RECT 129.200 213.600 130.000 213.700 ;
        RECT 158.000 213.600 158.800 213.700 ;
        RECT 159.600 214.300 160.400 214.400 ;
        RECT 169.200 214.300 170.000 214.400 ;
        RECT 188.400 214.300 189.200 214.400 ;
        RECT 196.400 214.300 197.200 214.400 ;
        RECT 159.600 213.700 170.000 214.300 ;
        RECT 159.600 213.600 160.400 213.700 ;
        RECT 169.200 213.600 170.000 213.700 ;
        RECT 180.500 213.700 197.200 214.300 ;
        RECT 180.500 212.400 181.100 213.700 ;
        RECT 188.400 213.600 189.200 213.700 ;
        RECT 196.400 213.600 197.200 213.700 ;
        RECT 199.600 214.300 200.400 214.400 ;
        RECT 209.200 214.300 210.000 214.400 ;
        RECT 199.600 213.700 210.000 214.300 ;
        RECT 199.600 213.600 200.400 213.700 ;
        RECT 209.200 213.600 210.000 213.700 ;
        RECT 220.400 214.300 221.200 214.400 ;
        RECT 286.000 214.300 286.800 214.400 ;
        RECT 220.400 213.700 286.800 214.300 ;
        RECT 220.400 213.600 221.200 213.700 ;
        RECT 286.000 213.600 286.800 213.700 ;
        RECT 311.600 214.300 312.400 214.400 ;
        RECT 332.400 214.300 333.200 214.400 ;
        RECT 311.600 213.700 333.200 214.300 ;
        RECT 311.600 213.600 312.400 213.700 ;
        RECT 332.400 213.600 333.200 213.700 ;
        RECT 380.400 214.300 381.200 214.400 ;
        RECT 385.200 214.300 386.000 214.400 ;
        RECT 380.400 213.700 386.000 214.300 ;
        RECT 380.400 213.600 381.200 213.700 ;
        RECT 385.200 213.600 386.000 213.700 ;
        RECT 394.800 214.300 395.600 214.400 ;
        RECT 399.700 214.300 400.300 215.700 ;
        RECT 407.600 215.600 408.400 215.700 ;
        RECT 410.800 215.600 411.600 216.400 ;
        RECT 436.400 216.300 437.200 216.400 ;
        RECT 444.400 216.300 445.200 216.400 ;
        RECT 436.400 215.700 445.200 216.300 ;
        RECT 436.400 215.600 437.200 215.700 ;
        RECT 444.400 215.600 445.200 215.700 ;
        RECT 446.000 216.300 446.800 216.400 ;
        RECT 447.600 216.300 448.400 216.400 ;
        RECT 446.000 215.700 448.400 216.300 ;
        RECT 446.000 215.600 446.800 215.700 ;
        RECT 447.600 215.600 448.400 215.700 ;
        RECT 513.200 216.300 514.000 216.400 ;
        RECT 530.800 216.300 531.600 216.400 ;
        RECT 513.200 215.700 531.600 216.300 ;
        RECT 513.200 215.600 514.000 215.700 ;
        RECT 530.800 215.600 531.600 215.700 ;
        RECT 394.800 213.700 400.300 214.300 ;
        RECT 401.200 214.300 402.000 214.400 ;
        RECT 452.400 214.300 453.200 214.400 ;
        RECT 401.200 213.700 453.200 214.300 ;
        RECT 394.800 213.600 395.600 213.700 ;
        RECT 401.200 213.600 402.000 213.700 ;
        RECT 452.400 213.600 453.200 213.700 ;
        RECT 454.000 214.300 454.800 214.400 ;
        RECT 455.600 214.300 456.400 214.400 ;
        RECT 454.000 213.700 456.400 214.300 ;
        RECT 454.000 213.600 454.800 213.700 ;
        RECT 455.600 213.600 456.400 213.700 ;
        RECT 462.000 214.300 462.800 214.400 ;
        RECT 527.600 214.300 528.400 214.400 ;
        RECT 542.000 214.300 542.800 214.400 ;
        RECT 462.000 213.700 465.900 214.300 ;
        RECT 462.000 213.600 462.800 213.700 ;
        RECT 465.300 212.400 465.900 213.700 ;
        RECT 527.600 213.700 542.800 214.300 ;
        RECT 527.600 213.600 528.400 213.700 ;
        RECT 542.000 213.600 542.800 213.700 ;
        RECT 17.200 212.300 18.000 212.400 ;
        RECT 34.800 212.300 35.600 212.400 ;
        RECT 17.200 211.700 35.600 212.300 ;
        RECT 17.200 211.600 18.000 211.700 ;
        RECT 34.800 211.600 35.600 211.700 ;
        RECT 39.600 212.300 40.400 212.400 ;
        RECT 44.400 212.300 45.200 212.400 ;
        RECT 39.600 211.700 45.200 212.300 ;
        RECT 39.600 211.600 40.400 211.700 ;
        RECT 44.400 211.600 45.200 211.700 ;
        RECT 47.600 212.300 48.400 212.400 ;
        RECT 76.400 212.300 77.200 212.400 ;
        RECT 47.600 211.700 77.200 212.300 ;
        RECT 47.600 211.600 48.400 211.700 ;
        RECT 76.400 211.600 77.200 211.700 ;
        RECT 87.600 212.300 88.400 212.400 ;
        RECT 92.400 212.300 93.200 212.400 ;
        RECT 87.600 211.700 93.200 212.300 ;
        RECT 87.600 211.600 88.400 211.700 ;
        RECT 92.400 211.600 93.200 211.700 ;
        RECT 154.800 212.300 155.600 212.400 ;
        RECT 161.200 212.300 162.000 212.400 ;
        RECT 180.400 212.300 181.200 212.400 ;
        RECT 154.800 211.700 181.200 212.300 ;
        RECT 154.800 211.600 155.600 211.700 ;
        RECT 161.200 211.600 162.000 211.700 ;
        RECT 180.400 211.600 181.200 211.700 ;
        RECT 183.600 212.300 184.400 212.400 ;
        RECT 191.600 212.300 192.400 212.400 ;
        RECT 183.600 211.700 192.400 212.300 ;
        RECT 183.600 211.600 184.400 211.700 ;
        RECT 191.600 211.600 192.400 211.700 ;
        RECT 198.000 212.300 198.800 212.400 ;
        RECT 204.400 212.300 205.200 212.400 ;
        RECT 198.000 211.700 205.200 212.300 ;
        RECT 198.000 211.600 198.800 211.700 ;
        RECT 204.400 211.600 205.200 211.700 ;
        RECT 222.000 212.300 222.800 212.400 ;
        RECT 246.000 212.300 246.800 212.400 ;
        RECT 222.000 211.700 246.800 212.300 ;
        RECT 222.000 211.600 222.800 211.700 ;
        RECT 246.000 211.600 246.800 211.700 ;
        RECT 276.400 212.300 277.200 212.400 ;
        RECT 318.000 212.300 318.800 212.400 ;
        RECT 276.400 211.700 318.800 212.300 ;
        RECT 276.400 211.600 277.200 211.700 ;
        RECT 318.000 211.600 318.800 211.700 ;
        RECT 330.800 212.300 331.600 212.400 ;
        RECT 335.600 212.300 336.400 212.400 ;
        RECT 330.800 211.700 336.400 212.300 ;
        RECT 330.800 211.600 331.600 211.700 ;
        RECT 335.600 211.600 336.400 211.700 ;
        RECT 367.600 212.300 368.400 212.400 ;
        RECT 372.400 212.300 373.200 212.400 ;
        RECT 391.600 212.300 392.400 212.400 ;
        RECT 398.000 212.300 398.800 212.400 ;
        RECT 367.600 211.700 398.800 212.300 ;
        RECT 367.600 211.600 368.400 211.700 ;
        RECT 372.400 211.600 373.200 211.700 ;
        RECT 391.600 211.600 392.400 211.700 ;
        RECT 398.000 211.600 398.800 211.700 ;
        RECT 409.200 212.300 410.000 212.400 ;
        RECT 415.600 212.300 416.400 212.400 ;
        RECT 409.200 211.700 416.400 212.300 ;
        RECT 409.200 211.600 410.000 211.700 ;
        RECT 415.600 211.600 416.400 211.700 ;
        RECT 434.800 212.300 435.600 212.400 ;
        RECT 463.600 212.300 464.400 212.400 ;
        RECT 434.800 211.700 464.400 212.300 ;
        RECT 434.800 211.600 435.600 211.700 ;
        RECT 463.600 211.600 464.400 211.700 ;
        RECT 465.200 211.600 466.000 212.400 ;
        RECT 471.600 212.300 472.400 212.400 ;
        RECT 478.000 212.300 478.800 212.400 ;
        RECT 487.600 212.300 488.400 212.400 ;
        RECT 471.600 211.700 488.400 212.300 ;
        RECT 471.600 211.600 472.400 211.700 ;
        RECT 478.000 211.600 478.800 211.700 ;
        RECT 487.600 211.600 488.400 211.700 ;
        RECT 497.200 212.300 498.000 212.400 ;
        RECT 506.800 212.300 507.600 212.400 ;
        RECT 518.000 212.300 518.800 212.400 ;
        RECT 497.200 211.700 518.800 212.300 ;
        RECT 497.200 211.600 498.000 211.700 ;
        RECT 506.800 211.600 507.600 211.700 ;
        RECT 518.000 211.600 518.800 211.700 ;
        RECT 535.600 212.300 536.400 212.400 ;
        RECT 540.400 212.300 541.200 212.400 ;
        RECT 535.600 211.700 541.200 212.300 ;
        RECT 535.600 211.600 536.400 211.700 ;
        RECT 540.400 211.600 541.200 211.700 ;
        RECT 26.800 210.300 27.600 210.400 ;
        RECT 38.000 210.300 38.800 210.400 ;
        RECT 26.800 209.700 38.800 210.300 ;
        RECT 26.800 209.600 27.600 209.700 ;
        RECT 38.000 209.600 38.800 209.700 ;
        RECT 46.000 210.300 46.800 210.400 ;
        RECT 52.400 210.300 53.200 210.400 ;
        RECT 46.000 209.700 53.200 210.300 ;
        RECT 46.000 209.600 46.800 209.700 ;
        RECT 52.400 209.600 53.200 209.700 ;
        RECT 71.600 210.300 72.400 210.400 ;
        RECT 81.200 210.300 82.000 210.400 ;
        RECT 71.600 209.700 82.000 210.300 ;
        RECT 71.600 209.600 72.400 209.700 ;
        RECT 81.200 209.600 82.000 209.700 ;
        RECT 100.400 210.300 101.200 210.400 ;
        RECT 108.400 210.300 109.200 210.400 ;
        RECT 100.400 209.700 109.200 210.300 ;
        RECT 100.400 209.600 101.200 209.700 ;
        RECT 108.400 209.600 109.200 209.700 ;
        RECT 151.600 210.300 152.400 210.400 ;
        RECT 166.000 210.300 166.800 210.400 ;
        RECT 151.600 209.700 166.800 210.300 ;
        RECT 151.600 209.600 152.400 209.700 ;
        RECT 166.000 209.600 166.800 209.700 ;
        RECT 206.000 210.300 206.800 210.400 ;
        RECT 217.200 210.300 218.000 210.400 ;
        RECT 206.000 209.700 218.000 210.300 ;
        RECT 206.000 209.600 206.800 209.700 ;
        RECT 217.200 209.600 218.000 209.700 ;
        RECT 225.200 210.300 226.000 210.400 ;
        RECT 239.600 210.300 240.400 210.400 ;
        RECT 225.200 209.700 240.400 210.300 ;
        RECT 225.200 209.600 226.000 209.700 ;
        RECT 239.600 209.600 240.400 209.700 ;
        RECT 241.200 210.300 242.000 210.400 ;
        RECT 266.800 210.300 267.600 210.400 ;
        RECT 241.200 209.700 267.600 210.300 ;
        RECT 241.200 209.600 242.000 209.700 ;
        RECT 266.800 209.600 267.600 209.700 ;
        RECT 346.800 210.300 347.600 210.400 ;
        RECT 350.000 210.300 350.800 210.400 ;
        RECT 346.800 209.700 350.800 210.300 ;
        RECT 346.800 209.600 347.600 209.700 ;
        RECT 350.000 209.600 350.800 209.700 ;
        RECT 358.000 210.300 358.800 210.400 ;
        RECT 375.600 210.300 376.400 210.400 ;
        RECT 358.000 209.700 376.400 210.300 ;
        RECT 358.000 209.600 358.800 209.700 ;
        RECT 375.600 209.600 376.400 209.700 ;
        RECT 382.000 210.300 382.800 210.400 ;
        RECT 412.400 210.300 413.200 210.400 ;
        RECT 382.000 209.700 413.200 210.300 ;
        RECT 382.000 209.600 382.800 209.700 ;
        RECT 412.400 209.600 413.200 209.700 ;
        RECT 428.400 210.300 429.200 210.400 ;
        RECT 447.600 210.300 448.400 210.400 ;
        RECT 428.400 209.700 448.400 210.300 ;
        RECT 428.400 209.600 429.200 209.700 ;
        RECT 447.600 209.600 448.400 209.700 ;
        RECT 449.200 210.300 450.000 210.400 ;
        RECT 474.800 210.300 475.600 210.400 ;
        RECT 449.200 209.700 475.600 210.300 ;
        RECT 449.200 209.600 450.000 209.700 ;
        RECT 474.800 209.600 475.600 209.700 ;
        RECT 12.400 208.300 13.200 208.400 ;
        RECT 25.200 208.300 26.000 208.400 ;
        RECT 12.400 207.700 26.000 208.300 ;
        RECT 12.400 207.600 13.200 207.700 ;
        RECT 25.200 207.600 26.000 207.700 ;
        RECT 42.800 208.300 43.600 208.400 ;
        RECT 62.000 208.300 62.800 208.400 ;
        RECT 42.800 207.700 62.800 208.300 ;
        RECT 42.800 207.600 43.600 207.700 ;
        RECT 62.000 207.600 62.800 207.700 ;
        RECT 68.400 208.300 69.200 208.400 ;
        RECT 105.200 208.300 106.000 208.400 ;
        RECT 68.400 207.700 106.000 208.300 ;
        RECT 68.400 207.600 69.200 207.700 ;
        RECT 105.200 207.600 106.000 207.700 ;
        RECT 191.600 208.300 192.400 208.400 ;
        RECT 202.800 208.300 203.600 208.400 ;
        RECT 191.600 207.700 203.600 208.300 ;
        RECT 191.600 207.600 192.400 207.700 ;
        RECT 202.800 207.600 203.600 207.700 ;
        RECT 228.400 208.300 229.200 208.400 ;
        RECT 233.200 208.300 234.000 208.400 ;
        RECT 228.400 207.700 234.000 208.300 ;
        RECT 228.400 207.600 229.200 207.700 ;
        RECT 233.200 207.600 234.000 207.700 ;
        RECT 239.600 208.300 240.400 208.400 ;
        RECT 242.800 208.300 243.600 208.400 ;
        RECT 239.600 207.700 243.600 208.300 ;
        RECT 239.600 207.600 240.400 207.700 ;
        RECT 242.800 207.600 243.600 207.700 ;
        RECT 364.400 208.300 365.200 208.400 ;
        RECT 370.800 208.300 371.600 208.400 ;
        RECT 375.600 208.300 376.400 208.400 ;
        RECT 380.400 208.300 381.200 208.400 ;
        RECT 364.400 207.700 381.200 208.300 ;
        RECT 364.400 207.600 365.200 207.700 ;
        RECT 370.800 207.600 371.600 207.700 ;
        RECT 375.600 207.600 376.400 207.700 ;
        RECT 380.400 207.600 381.200 207.700 ;
        RECT 382.000 208.300 382.800 208.400 ;
        RECT 402.800 208.300 403.600 208.400 ;
        RECT 382.000 207.700 403.600 208.300 ;
        RECT 382.000 207.600 382.800 207.700 ;
        RECT 402.800 207.600 403.600 207.700 ;
        RECT 407.600 208.300 408.400 208.400 ;
        RECT 410.800 208.300 411.600 208.400 ;
        RECT 407.600 207.700 411.600 208.300 ;
        RECT 407.600 207.600 408.400 207.700 ;
        RECT 410.800 207.600 411.600 207.700 ;
        RECT 414.000 208.300 414.800 208.400 ;
        RECT 444.400 208.300 445.200 208.400 ;
        RECT 414.000 207.700 445.200 208.300 ;
        RECT 414.000 207.600 414.800 207.700 ;
        RECT 444.400 207.600 445.200 207.700 ;
        RECT 446.000 208.300 446.800 208.400 ;
        RECT 449.200 208.300 450.000 208.400 ;
        RECT 446.000 207.700 450.000 208.300 ;
        RECT 446.000 207.600 446.800 207.700 ;
        RECT 449.200 207.600 450.000 207.700 ;
        RECT 23.600 206.300 24.400 206.400 ;
        RECT 42.800 206.300 43.600 206.400 ;
        RECT 23.600 205.700 43.600 206.300 ;
        RECT 23.600 205.600 24.400 205.700 ;
        RECT 42.800 205.600 43.600 205.700 ;
        RECT 44.400 206.300 45.200 206.400 ;
        RECT 63.600 206.300 64.400 206.400 ;
        RECT 44.400 205.700 64.400 206.300 ;
        RECT 44.400 205.600 45.200 205.700 ;
        RECT 63.600 205.600 64.400 205.700 ;
        RECT 225.200 206.300 226.000 206.400 ;
        RECT 228.400 206.300 229.200 206.400 ;
        RECT 225.200 205.700 229.200 206.300 ;
        RECT 225.200 205.600 226.000 205.700 ;
        RECT 228.400 205.600 229.200 205.700 ;
        RECT 231.600 206.300 232.400 206.400 ;
        RECT 234.800 206.300 235.600 206.400 ;
        RECT 231.600 205.700 235.600 206.300 ;
        RECT 231.600 205.600 232.400 205.700 ;
        RECT 234.800 205.600 235.600 205.700 ;
        RECT 247.600 206.300 248.400 206.400 ;
        RECT 255.600 206.300 256.400 206.400 ;
        RECT 247.600 205.700 256.400 206.300 ;
        RECT 247.600 205.600 248.400 205.700 ;
        RECT 255.600 205.600 256.400 205.700 ;
        RECT 380.400 206.300 381.200 206.400 ;
        RECT 404.400 206.300 405.200 206.400 ;
        RECT 417.200 206.300 418.000 206.400 ;
        RECT 455.600 206.300 456.400 206.400 ;
        RECT 478.000 206.300 478.800 206.400 ;
        RECT 489.200 206.300 490.000 206.400 ;
        RECT 380.400 205.700 490.000 206.300 ;
        RECT 380.400 205.600 381.200 205.700 ;
        RECT 404.400 205.600 405.200 205.700 ;
        RECT 417.200 205.600 418.000 205.700 ;
        RECT 455.600 205.600 456.400 205.700 ;
        RECT 478.000 205.600 478.800 205.700 ;
        RECT 489.200 205.600 490.000 205.700 ;
        RECT 38.000 204.300 38.800 204.400 ;
        RECT 74.800 204.300 75.600 204.400 ;
        RECT 38.000 203.700 75.600 204.300 ;
        RECT 38.000 203.600 38.800 203.700 ;
        RECT 74.800 203.600 75.600 203.700 ;
        RECT 214.000 204.300 214.800 204.400 ;
        RECT 250.800 204.300 251.600 204.400 ;
        RECT 292.400 204.300 293.200 204.400 ;
        RECT 214.000 203.700 293.200 204.300 ;
        RECT 214.000 203.600 214.800 203.700 ;
        RECT 250.800 203.600 251.600 203.700 ;
        RECT 292.400 203.600 293.200 203.700 ;
        RECT 369.200 204.300 370.000 204.400 ;
        RECT 399.600 204.300 400.400 204.400 ;
        RECT 369.200 203.700 400.400 204.300 ;
        RECT 369.200 203.600 370.000 203.700 ;
        RECT 399.600 203.600 400.400 203.700 ;
        RECT 441.200 204.300 442.000 204.400 ;
        RECT 458.800 204.300 459.600 204.400 ;
        RECT 522.800 204.300 523.600 204.400 ;
        RECT 441.200 203.700 523.600 204.300 ;
        RECT 441.200 203.600 442.000 203.700 ;
        RECT 458.800 203.600 459.600 203.700 ;
        RECT 522.800 203.600 523.600 203.700 ;
        RECT 42.800 202.300 43.600 202.400 ;
        RECT 50.800 202.300 51.600 202.400 ;
        RECT 42.800 201.700 51.600 202.300 ;
        RECT 42.800 201.600 43.600 201.700 ;
        RECT 50.800 201.600 51.600 201.700 ;
        RECT 60.400 202.300 61.200 202.400 ;
        RECT 63.600 202.300 64.400 202.400 ;
        RECT 60.400 201.700 64.400 202.300 ;
        RECT 60.400 201.600 61.200 201.700 ;
        RECT 63.600 201.600 64.400 201.700 ;
        RECT 258.800 202.300 259.600 202.400 ;
        RECT 260.400 202.300 261.200 202.400 ;
        RECT 258.800 201.700 261.200 202.300 ;
        RECT 258.800 201.600 259.600 201.700 ;
        RECT 260.400 201.600 261.200 201.700 ;
        RECT 388.400 202.300 389.200 202.400 ;
        RECT 414.000 202.300 414.800 202.400 ;
        RECT 388.400 201.700 414.800 202.300 ;
        RECT 388.400 201.600 389.200 201.700 ;
        RECT 414.000 201.600 414.800 201.700 ;
        RECT 460.400 202.300 461.200 202.400 ;
        RECT 462.000 202.300 462.800 202.400 ;
        RECT 460.400 201.700 462.800 202.300 ;
        RECT 460.400 201.600 461.200 201.700 ;
        RECT 462.000 201.600 462.800 201.700 ;
        RECT 518.000 202.300 518.800 202.400 ;
        RECT 522.800 202.300 523.600 202.400 ;
        RECT 518.000 201.700 523.600 202.300 ;
        RECT 518.000 201.600 518.800 201.700 ;
        RECT 522.800 201.600 523.600 201.700 ;
        RECT 33.200 200.300 34.000 200.400 ;
        RECT 62.000 200.300 62.800 200.400 ;
        RECT 33.200 199.700 62.800 200.300 ;
        RECT 33.200 199.600 34.000 199.700 ;
        RECT 62.000 199.600 62.800 199.700 ;
        RECT 63.600 200.300 64.400 200.400 ;
        RECT 70.000 200.300 70.800 200.400 ;
        RECT 63.600 199.700 70.800 200.300 ;
        RECT 63.600 199.600 64.400 199.700 ;
        RECT 70.000 199.600 70.800 199.700 ;
        RECT 73.200 200.300 74.000 200.400 ;
        RECT 94.000 200.300 94.800 200.400 ;
        RECT 73.200 199.700 94.800 200.300 ;
        RECT 73.200 199.600 74.000 199.700 ;
        RECT 94.000 199.600 94.800 199.700 ;
        RECT 98.800 200.300 99.600 200.400 ;
        RECT 100.400 200.300 101.200 200.400 ;
        RECT 98.800 199.700 101.200 200.300 ;
        RECT 98.800 199.600 99.600 199.700 ;
        RECT 100.400 199.600 101.200 199.700 ;
        RECT 150.000 200.300 150.800 200.400 ;
        RECT 175.600 200.300 176.400 200.400 ;
        RECT 150.000 199.700 176.400 200.300 ;
        RECT 150.000 199.600 150.800 199.700 ;
        RECT 175.600 199.600 176.400 199.700 ;
        RECT 342.000 200.300 342.800 200.400 ;
        RECT 348.400 200.300 349.200 200.400 ;
        RECT 342.000 199.700 349.200 200.300 ;
        RECT 342.000 199.600 342.800 199.700 ;
        RECT 348.400 199.600 349.200 199.700 ;
        RECT 394.800 200.300 395.600 200.400 ;
        RECT 410.800 200.300 411.600 200.400 ;
        RECT 394.800 199.700 411.600 200.300 ;
        RECT 394.800 199.600 395.600 199.700 ;
        RECT 410.800 199.600 411.600 199.700 ;
        RECT 442.800 200.300 443.600 200.400 ;
        RECT 465.200 200.300 466.000 200.400 ;
        RECT 442.800 199.700 466.000 200.300 ;
        RECT 442.800 199.600 443.600 199.700 ;
        RECT 465.200 199.600 466.000 199.700 ;
        RECT 481.200 200.300 482.000 200.400 ;
        RECT 500.400 200.300 501.200 200.400 ;
        RECT 481.200 199.700 501.200 200.300 ;
        RECT 481.200 199.600 482.000 199.700 ;
        RECT 500.400 199.600 501.200 199.700 ;
        RECT 49.200 198.300 50.000 198.400 ;
        RECT 57.200 198.300 58.000 198.400 ;
        RECT 82.800 198.300 83.600 198.400 ;
        RECT 49.200 197.700 83.600 198.300 ;
        RECT 49.200 197.600 50.000 197.700 ;
        RECT 57.200 197.600 58.000 197.700 ;
        RECT 82.800 197.600 83.600 197.700 ;
        RECT 98.800 198.300 99.600 198.400 ;
        RECT 110.000 198.300 110.800 198.400 ;
        RECT 98.800 197.700 110.800 198.300 ;
        RECT 98.800 197.600 99.600 197.700 ;
        RECT 110.000 197.600 110.800 197.700 ;
        RECT 180.400 198.300 181.200 198.400 ;
        RECT 183.600 198.300 184.400 198.400 ;
        RECT 180.400 197.700 184.400 198.300 ;
        RECT 180.400 197.600 181.200 197.700 ;
        RECT 183.600 197.600 184.400 197.700 ;
        RECT 378.800 198.300 379.600 198.400 ;
        RECT 418.800 198.300 419.600 198.400 ;
        RECT 378.800 197.700 419.600 198.300 ;
        RECT 378.800 197.600 379.600 197.700 ;
        RECT 418.800 197.600 419.600 197.700 ;
        RECT 468.400 198.300 469.200 198.400 ;
        RECT 489.200 198.300 490.000 198.400 ;
        RECT 468.400 197.700 490.000 198.300 ;
        RECT 468.400 197.600 469.200 197.700 ;
        RECT 489.200 197.600 490.000 197.700 ;
        RECT 31.600 196.300 32.400 196.400 ;
        RECT 54.000 196.300 54.800 196.400 ;
        RECT 31.600 195.700 54.800 196.300 ;
        RECT 31.600 195.600 32.400 195.700 ;
        RECT 54.000 195.600 54.800 195.700 ;
        RECT 95.600 196.300 96.400 196.400 ;
        RECT 98.800 196.300 99.600 196.400 ;
        RECT 95.600 195.700 99.600 196.300 ;
        RECT 95.600 195.600 96.400 195.700 ;
        RECT 98.800 195.600 99.600 195.700 ;
        RECT 142.000 196.300 142.800 196.400 ;
        RECT 295.600 196.300 296.400 196.400 ;
        RECT 142.000 195.700 296.400 196.300 ;
        RECT 142.000 195.600 142.800 195.700 ;
        RECT 295.600 195.600 296.400 195.700 ;
        RECT 334.000 196.300 334.800 196.400 ;
        RECT 458.800 196.300 459.600 196.400 ;
        RECT 334.000 195.700 459.600 196.300 ;
        RECT 334.000 195.600 334.800 195.700 ;
        RECT 458.800 195.600 459.600 195.700 ;
        RECT 31.600 194.300 32.400 194.400 ;
        RECT 33.200 194.300 34.000 194.400 ;
        RECT 31.600 193.700 34.000 194.300 ;
        RECT 31.600 193.600 32.400 193.700 ;
        RECT 33.200 193.600 34.000 193.700 ;
        RECT 46.000 194.300 46.800 194.400 ;
        RECT 52.400 194.300 53.200 194.400 ;
        RECT 46.000 193.700 53.200 194.300 ;
        RECT 46.000 193.600 46.800 193.700 ;
        RECT 52.400 193.600 53.200 193.700 ;
        RECT 218.800 194.300 219.600 194.400 ;
        RECT 225.200 194.300 226.000 194.400 ;
        RECT 218.800 193.700 226.000 194.300 ;
        RECT 218.800 193.600 219.600 193.700 ;
        RECT 225.200 193.600 226.000 193.700 ;
        RECT 228.400 194.300 229.200 194.400 ;
        RECT 337.200 194.300 338.000 194.400 ;
        RECT 228.400 193.700 338.000 194.300 ;
        RECT 228.400 193.600 229.200 193.700 ;
        RECT 337.200 193.600 338.000 193.700 ;
        RECT 353.200 194.300 354.000 194.400 ;
        RECT 390.000 194.300 390.800 194.400 ;
        RECT 353.200 193.700 390.800 194.300 ;
        RECT 353.200 193.600 354.000 193.700 ;
        RECT 390.000 193.600 390.800 193.700 ;
        RECT 391.600 194.300 392.400 194.400 ;
        RECT 394.800 194.300 395.600 194.400 ;
        RECT 391.600 193.700 395.600 194.300 ;
        RECT 391.600 193.600 392.400 193.700 ;
        RECT 394.800 193.600 395.600 193.700 ;
        RECT 401.200 194.300 402.000 194.400 ;
        RECT 407.600 194.300 408.400 194.400 ;
        RECT 401.200 193.700 408.400 194.300 ;
        RECT 401.200 193.600 402.000 193.700 ;
        RECT 407.600 193.600 408.400 193.700 ;
        RECT 412.400 194.300 413.200 194.400 ;
        RECT 415.600 194.300 416.400 194.400 ;
        RECT 412.400 193.700 416.400 194.300 ;
        RECT 412.400 193.600 413.200 193.700 ;
        RECT 415.600 193.600 416.400 193.700 ;
        RECT 418.800 194.300 419.600 194.400 ;
        RECT 418.800 193.700 433.900 194.300 ;
        RECT 418.800 193.600 419.600 193.700 ;
        RECT 433.300 192.400 433.900 193.700 ;
        RECT 436.400 193.600 437.200 194.400 ;
        RECT 446.000 194.300 446.800 194.400 ;
        RECT 460.400 194.300 461.200 194.400 ;
        RECT 463.600 194.300 464.400 194.400 ;
        RECT 446.000 193.700 464.400 194.300 ;
        RECT 446.000 193.600 446.800 193.700 ;
        RECT 460.400 193.600 461.200 193.700 ;
        RECT 463.600 193.600 464.400 193.700 ;
        RECT 6.000 192.300 6.800 192.400 ;
        RECT 10.800 192.300 11.600 192.400 ;
        RECT 6.000 191.700 11.600 192.300 ;
        RECT 6.000 191.600 6.800 191.700 ;
        RECT 10.800 191.600 11.600 191.700 ;
        RECT 34.800 192.300 35.600 192.400 ;
        RECT 58.800 192.300 59.600 192.400 ;
        RECT 66.800 192.300 67.600 192.400 ;
        RECT 34.800 191.700 67.600 192.300 ;
        RECT 34.800 191.600 35.600 191.700 ;
        RECT 58.800 191.600 59.600 191.700 ;
        RECT 66.800 191.600 67.600 191.700 ;
        RECT 90.800 192.300 91.600 192.400 ;
        RECT 129.200 192.300 130.000 192.400 ;
        RECT 148.400 192.300 149.200 192.400 ;
        RECT 90.800 191.700 149.200 192.300 ;
        RECT 90.800 191.600 91.600 191.700 ;
        RECT 129.200 191.600 130.000 191.700 ;
        RECT 148.400 191.600 149.200 191.700 ;
        RECT 228.400 192.300 229.200 192.400 ;
        RECT 231.600 192.300 232.400 192.400 ;
        RECT 247.600 192.300 248.400 192.400 ;
        RECT 282.800 192.300 283.600 192.400 ;
        RECT 228.400 191.700 283.600 192.300 ;
        RECT 228.400 191.600 229.200 191.700 ;
        RECT 231.600 191.600 232.400 191.700 ;
        RECT 247.600 191.600 248.400 191.700 ;
        RECT 282.800 191.600 283.600 191.700 ;
        RECT 377.200 192.300 378.000 192.400 ;
        RECT 401.200 192.300 402.000 192.400 ;
        RECT 377.200 191.700 402.000 192.300 ;
        RECT 377.200 191.600 378.000 191.700 ;
        RECT 401.200 191.600 402.000 191.700 ;
        RECT 410.800 192.300 411.600 192.400 ;
        RECT 414.000 192.300 414.800 192.400 ;
        RECT 423.600 192.300 424.400 192.400 ;
        RECT 410.800 191.700 424.400 192.300 ;
        RECT 410.800 191.600 411.600 191.700 ;
        RECT 414.000 191.600 414.800 191.700 ;
        RECT 423.600 191.600 424.400 191.700 ;
        RECT 433.200 192.300 434.000 192.400 ;
        RECT 436.400 192.300 437.200 192.400 ;
        RECT 433.200 191.700 437.200 192.300 ;
        RECT 433.200 191.600 434.000 191.700 ;
        RECT 436.400 191.600 437.200 191.700 ;
        RECT 500.400 192.300 501.200 192.400 ;
        RECT 516.400 192.300 517.200 192.400 ;
        RECT 500.400 191.700 517.200 192.300 ;
        RECT 500.400 191.600 501.200 191.700 ;
        RECT 516.400 191.600 517.200 191.700 ;
        RECT 519.600 192.300 520.400 192.400 ;
        RECT 532.400 192.300 533.200 192.400 ;
        RECT 546.800 192.300 547.600 192.400 ;
        RECT 519.600 191.700 547.600 192.300 ;
        RECT 519.600 191.600 520.400 191.700 ;
        RECT 532.400 191.600 533.200 191.700 ;
        RECT 546.800 191.600 547.600 191.700 ;
        RECT 4.400 190.300 5.200 190.400 ;
        RECT 6.000 190.300 6.800 190.400 ;
        RECT 22.000 190.300 22.800 190.400 ;
        RECT 4.400 189.700 22.800 190.300 ;
        RECT 4.400 189.600 5.200 189.700 ;
        RECT 6.000 189.600 6.800 189.700 ;
        RECT 22.000 189.600 22.800 189.700 ;
        RECT 49.200 190.300 50.000 190.400 ;
        RECT 81.200 190.300 82.000 190.400 ;
        RECT 49.200 189.700 82.000 190.300 ;
        RECT 49.200 189.600 50.000 189.700 ;
        RECT 81.200 189.600 82.000 189.700 ;
        RECT 175.600 190.300 176.400 190.400 ;
        RECT 191.600 190.300 192.400 190.400 ;
        RECT 175.600 189.700 192.400 190.300 ;
        RECT 175.600 189.600 176.400 189.700 ;
        RECT 191.600 189.600 192.400 189.700 ;
        RECT 218.800 190.300 219.600 190.400 ;
        RECT 223.600 190.300 224.400 190.400 ;
        RECT 218.800 189.700 224.400 190.300 ;
        RECT 218.800 189.600 219.600 189.700 ;
        RECT 223.600 189.600 224.400 189.700 ;
        RECT 234.800 190.300 235.600 190.400 ;
        RECT 252.400 190.300 253.200 190.400 ;
        RECT 268.400 190.300 269.200 190.400 ;
        RECT 234.800 189.700 269.200 190.300 ;
        RECT 234.800 189.600 235.600 189.700 ;
        RECT 252.400 189.600 253.200 189.700 ;
        RECT 268.400 189.600 269.200 189.700 ;
        RECT 337.200 190.300 338.000 190.400 ;
        RECT 375.600 190.300 376.400 190.400 ;
        RECT 378.800 190.300 379.600 190.400 ;
        RECT 337.200 189.700 379.600 190.300 ;
        RECT 337.200 189.600 338.000 189.700 ;
        RECT 375.600 189.600 376.400 189.700 ;
        RECT 378.800 189.600 379.600 189.700 ;
        RECT 388.400 190.300 389.200 190.400 ;
        RECT 398.000 190.300 398.800 190.400 ;
        RECT 388.400 189.700 398.800 190.300 ;
        RECT 388.400 189.600 389.200 189.700 ;
        RECT 398.000 189.600 398.800 189.700 ;
        RECT 404.400 190.300 405.200 190.400 ;
        RECT 434.800 190.300 435.600 190.400 ;
        RECT 404.400 189.700 435.600 190.300 ;
        RECT 404.400 189.600 405.200 189.700 ;
        RECT 434.800 189.600 435.600 189.700 ;
        RECT 465.200 189.600 466.000 190.400 ;
        RECT 466.800 190.300 467.600 190.400 ;
        RECT 481.200 190.300 482.000 190.400 ;
        RECT 466.800 189.700 482.000 190.300 ;
        RECT 466.800 189.600 467.600 189.700 ;
        RECT 481.200 189.600 482.000 189.700 ;
        RECT 503.600 190.300 504.400 190.400 ;
        RECT 511.600 190.300 512.400 190.400 ;
        RECT 503.600 189.700 512.400 190.300 ;
        RECT 503.600 189.600 504.400 189.700 ;
        RECT 511.600 189.600 512.400 189.700 ;
        RECT 513.200 190.300 514.000 190.400 ;
        RECT 550.000 190.300 550.800 190.400 ;
        RECT 513.200 189.700 550.800 190.300 ;
        RECT 513.200 189.600 514.000 189.700 ;
        RECT 550.000 189.600 550.800 189.700 ;
        RECT 1.200 188.300 2.000 188.400 ;
        RECT 17.200 188.300 18.000 188.400 ;
        RECT 1.200 187.700 18.000 188.300 ;
        RECT 1.200 187.600 2.000 187.700 ;
        RECT 17.200 187.600 18.000 187.700 ;
        RECT 26.800 188.300 27.600 188.400 ;
        RECT 34.800 188.300 35.600 188.400 ;
        RECT 26.800 187.700 35.600 188.300 ;
        RECT 26.800 187.600 27.600 187.700 ;
        RECT 34.800 187.600 35.600 187.700 ;
        RECT 65.200 188.300 66.000 188.400 ;
        RECT 79.600 188.300 80.400 188.400 ;
        RECT 65.200 187.700 80.400 188.300 ;
        RECT 65.200 187.600 66.000 187.700 ;
        RECT 79.600 187.600 80.400 187.700 ;
        RECT 122.800 188.300 123.600 188.400 ;
        RECT 132.400 188.300 133.200 188.400 ;
        RECT 122.800 187.700 133.200 188.300 ;
        RECT 122.800 187.600 123.600 187.700 ;
        RECT 132.400 187.600 133.200 187.700 ;
        RECT 218.800 188.300 219.600 188.400 ;
        RECT 230.000 188.300 230.800 188.400 ;
        RECT 238.000 188.300 238.800 188.400 ;
        RECT 218.800 187.700 238.800 188.300 ;
        RECT 218.800 187.600 219.600 187.700 ;
        RECT 230.000 187.600 230.800 187.700 ;
        RECT 238.000 187.600 238.800 187.700 ;
        RECT 266.800 188.300 267.600 188.400 ;
        RECT 287.600 188.300 288.400 188.400 ;
        RECT 266.800 187.700 288.400 188.300 ;
        RECT 266.800 187.600 267.600 187.700 ;
        RECT 287.600 187.600 288.400 187.700 ;
        RECT 345.200 188.300 346.000 188.400 ;
        RECT 359.600 188.300 360.400 188.400 ;
        RECT 345.200 187.700 360.400 188.300 ;
        RECT 345.200 187.600 346.000 187.700 ;
        RECT 359.600 187.600 360.400 187.700 ;
        RECT 386.800 188.300 387.600 188.400 ;
        RECT 399.600 188.300 400.400 188.400 ;
        RECT 386.800 187.700 400.400 188.300 ;
        RECT 386.800 187.600 387.600 187.700 ;
        RECT 399.600 187.600 400.400 187.700 ;
        RECT 401.200 188.300 402.000 188.400 ;
        RECT 410.800 188.300 411.600 188.400 ;
        RECT 433.200 188.300 434.000 188.400 ;
        RECT 447.600 188.300 448.400 188.400 ;
        RECT 401.200 187.700 409.900 188.300 ;
        RECT 401.200 187.600 402.000 187.700 ;
        RECT 9.200 186.300 10.000 186.400 ;
        RECT 14.000 186.300 14.800 186.400 ;
        RECT 22.000 186.300 22.800 186.400 ;
        RECT 30.000 186.300 30.800 186.400 ;
        RECT 9.200 185.700 30.800 186.300 ;
        RECT 9.200 185.600 10.000 185.700 ;
        RECT 14.000 185.600 14.800 185.700 ;
        RECT 22.000 185.600 22.800 185.700 ;
        RECT 30.000 185.600 30.800 185.700 ;
        RECT 44.400 186.300 45.200 186.400 ;
        RECT 47.600 186.300 48.400 186.400 ;
        RECT 44.400 185.700 48.400 186.300 ;
        RECT 44.400 185.600 45.200 185.700 ;
        RECT 47.600 185.600 48.400 185.700 ;
        RECT 49.200 186.300 50.000 186.400 ;
        RECT 57.200 186.300 58.000 186.400 ;
        RECT 92.400 186.300 93.200 186.400 ;
        RECT 49.200 185.700 93.200 186.300 ;
        RECT 49.200 185.600 50.000 185.700 ;
        RECT 57.200 185.600 58.000 185.700 ;
        RECT 92.400 185.600 93.200 185.700 ;
        RECT 159.600 186.300 160.400 186.400 ;
        RECT 167.600 186.300 168.400 186.400 ;
        RECT 159.600 185.700 168.400 186.300 ;
        RECT 159.600 185.600 160.400 185.700 ;
        RECT 167.600 185.600 168.400 185.700 ;
        RECT 222.000 186.300 222.800 186.400 ;
        RECT 230.000 186.300 230.800 186.400 ;
        RECT 222.000 185.700 230.800 186.300 ;
        RECT 222.000 185.600 222.800 185.700 ;
        RECT 230.000 185.600 230.800 185.700 ;
        RECT 249.200 186.300 250.000 186.400 ;
        RECT 262.000 186.300 262.800 186.400 ;
        RECT 249.200 185.700 262.800 186.300 ;
        RECT 249.200 185.600 250.000 185.700 ;
        RECT 262.000 185.600 262.800 185.700 ;
        RECT 335.600 186.300 336.400 186.400 ;
        RECT 338.800 186.300 339.600 186.400 ;
        RECT 342.000 186.300 342.800 186.400 ;
        RECT 343.600 186.300 344.400 186.400 ;
        RECT 359.600 186.300 360.400 186.400 ;
        RECT 380.400 186.300 381.200 186.400 ;
        RECT 335.600 185.700 381.200 186.300 ;
        RECT 335.600 185.600 336.400 185.700 ;
        RECT 338.800 185.600 339.600 185.700 ;
        RECT 342.000 185.600 342.800 185.700 ;
        RECT 343.600 185.600 344.400 185.700 ;
        RECT 359.600 185.600 360.400 185.700 ;
        RECT 380.400 185.600 381.200 185.700 ;
        RECT 385.200 186.300 386.000 186.400 ;
        RECT 394.800 186.300 395.600 186.400 ;
        RECT 385.200 185.700 395.600 186.300 ;
        RECT 409.300 186.300 409.900 187.700 ;
        RECT 410.800 187.700 448.400 188.300 ;
        RECT 410.800 187.600 411.600 187.700 ;
        RECT 433.200 187.600 434.000 187.700 ;
        RECT 447.600 187.600 448.400 187.700 ;
        RECT 458.800 188.300 459.600 188.400 ;
        RECT 462.000 188.300 462.800 188.400 ;
        RECT 458.800 187.700 462.800 188.300 ;
        RECT 458.800 187.600 459.600 187.700 ;
        RECT 462.000 187.600 462.800 187.700 ;
        RECT 474.800 188.300 475.600 188.400 ;
        RECT 498.800 188.300 499.600 188.400 ;
        RECT 505.200 188.300 506.000 188.400 ;
        RECT 474.800 187.700 506.000 188.300 ;
        RECT 474.800 187.600 475.600 187.700 ;
        RECT 498.800 187.600 499.600 187.700 ;
        RECT 505.200 187.600 506.000 187.700 ;
        RECT 514.800 188.300 515.600 188.400 ;
        RECT 518.000 188.300 518.800 188.400 ;
        RECT 538.800 188.300 539.600 188.400 ;
        RECT 514.800 187.700 539.600 188.300 ;
        RECT 514.800 187.600 515.600 187.700 ;
        RECT 518.000 187.600 518.800 187.700 ;
        RECT 538.800 187.600 539.600 187.700 ;
        RECT 412.400 186.300 413.200 186.400 ;
        RECT 409.300 185.700 413.200 186.300 ;
        RECT 385.200 185.600 386.000 185.700 ;
        RECT 394.800 185.600 395.600 185.700 ;
        RECT 412.400 185.600 413.200 185.700 ;
        RECT 431.600 186.300 432.400 186.400 ;
        RECT 500.400 186.300 501.200 186.400 ;
        RECT 431.600 185.700 501.200 186.300 ;
        RECT 431.600 185.600 432.400 185.700 ;
        RECT 500.400 185.600 501.200 185.700 ;
        RECT 52.400 183.600 53.200 184.400 ;
        RECT 223.600 184.300 224.400 184.400 ;
        RECT 268.400 184.300 269.200 184.400 ;
        RECT 223.600 183.700 269.200 184.300 ;
        RECT 223.600 183.600 224.400 183.700 ;
        RECT 268.400 183.600 269.200 183.700 ;
        RECT 362.800 184.300 363.600 184.400 ;
        RECT 380.400 184.300 381.200 184.400 ;
        RECT 434.800 184.300 435.600 184.400 ;
        RECT 486.000 184.300 486.800 184.400 ;
        RECT 362.800 183.700 486.800 184.300 ;
        RECT 362.800 183.600 363.600 183.700 ;
        RECT 380.400 183.600 381.200 183.700 ;
        RECT 434.800 183.600 435.600 183.700 ;
        RECT 486.000 183.600 486.800 183.700 ;
        RECT 521.200 184.300 522.000 184.400 ;
        RECT 542.000 184.300 542.800 184.400 ;
        RECT 521.200 183.700 542.800 184.300 ;
        RECT 521.200 183.600 522.000 183.700 ;
        RECT 542.000 183.600 542.800 183.700 ;
        RECT 26.800 182.300 27.600 182.400 ;
        RECT 28.400 182.300 29.200 182.400 ;
        RECT 26.800 181.700 29.200 182.300 ;
        RECT 26.800 181.600 27.600 181.700 ;
        RECT 28.400 181.600 29.200 181.700 ;
        RECT 52.400 182.300 53.200 182.400 ;
        RECT 55.600 182.300 56.400 182.400 ;
        RECT 52.400 181.700 56.400 182.300 ;
        RECT 52.400 181.600 53.200 181.700 ;
        RECT 55.600 181.600 56.400 181.700 ;
        RECT 174.000 182.300 174.800 182.400 ;
        RECT 212.400 182.300 213.200 182.400 ;
        RECT 174.000 181.700 213.200 182.300 ;
        RECT 174.000 181.600 174.800 181.700 ;
        RECT 212.400 181.600 213.200 181.700 ;
        RECT 226.800 182.300 227.600 182.400 ;
        RECT 270.000 182.300 270.800 182.400 ;
        RECT 226.800 181.700 270.800 182.300 ;
        RECT 226.800 181.600 227.600 181.700 ;
        RECT 270.000 181.600 270.800 181.700 ;
        RECT 297.200 182.300 298.000 182.400 ;
        RECT 324.400 182.300 325.200 182.400 ;
        RECT 332.400 182.300 333.200 182.400 ;
        RECT 353.200 182.300 354.000 182.400 ;
        RECT 388.400 182.300 389.200 182.400 ;
        RECT 447.600 182.300 448.400 182.400 ;
        RECT 454.000 182.300 454.800 182.400 ;
        RECT 478.000 182.300 478.800 182.400 ;
        RECT 297.200 181.700 478.800 182.300 ;
        RECT 297.200 181.600 298.000 181.700 ;
        RECT 324.400 181.600 325.200 181.700 ;
        RECT 332.400 181.600 333.200 181.700 ;
        RECT 353.200 181.600 354.000 181.700 ;
        RECT 388.400 181.600 389.200 181.700 ;
        RECT 447.600 181.600 448.400 181.700 ;
        RECT 454.000 181.600 454.800 181.700 ;
        RECT 478.000 181.600 478.800 181.700 ;
        RECT 487.600 182.300 488.400 182.400 ;
        RECT 508.400 182.300 509.200 182.400 ;
        RECT 487.600 181.700 509.200 182.300 ;
        RECT 487.600 181.600 488.400 181.700 ;
        RECT 508.400 181.600 509.200 181.700 ;
        RECT 511.600 182.300 512.400 182.400 ;
        RECT 527.600 182.300 528.400 182.400 ;
        RECT 511.600 181.700 528.400 182.300 ;
        RECT 511.600 181.600 512.400 181.700 ;
        RECT 527.600 181.600 528.400 181.700 ;
        RECT 20.400 180.300 21.200 180.400 ;
        RECT 28.400 180.300 29.200 180.400 ;
        RECT 54.000 180.300 54.800 180.400 ;
        RECT 20.400 179.700 54.800 180.300 ;
        RECT 20.400 179.600 21.200 179.700 ;
        RECT 28.400 179.600 29.200 179.700 ;
        RECT 54.000 179.600 54.800 179.700 ;
        RECT 233.200 180.300 234.000 180.400 ;
        RECT 260.400 180.300 261.200 180.400 ;
        RECT 233.200 179.700 261.200 180.300 ;
        RECT 233.200 179.600 234.000 179.700 ;
        RECT 260.400 179.600 261.200 179.700 ;
        RECT 332.400 180.300 333.200 180.400 ;
        RECT 410.800 180.300 411.600 180.400 ;
        RECT 332.400 179.700 411.600 180.300 ;
        RECT 332.400 179.600 333.200 179.700 ;
        RECT 410.800 179.600 411.600 179.700 ;
        RECT 417.200 180.300 418.000 180.400 ;
        RECT 431.600 180.300 432.400 180.400 ;
        RECT 417.200 179.700 432.400 180.300 ;
        RECT 417.200 179.600 418.000 179.700 ;
        RECT 431.600 179.600 432.400 179.700 ;
        RECT 468.400 180.300 469.200 180.400 ;
        RECT 476.400 180.300 477.200 180.400 ;
        RECT 468.400 179.700 477.200 180.300 ;
        RECT 468.400 179.600 469.200 179.700 ;
        RECT 476.400 179.600 477.200 179.700 ;
        RECT 478.000 180.300 478.800 180.400 ;
        RECT 481.200 180.300 482.000 180.400 ;
        RECT 478.000 179.700 482.000 180.300 ;
        RECT 478.000 179.600 478.800 179.700 ;
        RECT 481.200 179.600 482.000 179.700 ;
        RECT 538.800 180.300 539.600 180.400 ;
        RECT 545.200 180.300 546.000 180.400 ;
        RECT 538.800 179.700 546.000 180.300 ;
        RECT 538.800 179.600 539.600 179.700 ;
        RECT 545.200 179.600 546.000 179.700 ;
        RECT 23.600 178.300 24.400 178.400 ;
        RECT 57.200 178.300 58.000 178.400 ;
        RECT 23.600 177.700 58.000 178.300 ;
        RECT 23.600 177.600 24.400 177.700 ;
        RECT 57.200 177.600 58.000 177.700 ;
        RECT 73.200 178.300 74.000 178.400 ;
        RECT 82.800 178.300 83.600 178.400 ;
        RECT 119.600 178.300 120.400 178.400 ;
        RECT 134.000 178.300 134.800 178.400 ;
        RECT 73.200 177.700 134.800 178.300 ;
        RECT 73.200 177.600 74.000 177.700 ;
        RECT 82.800 177.600 83.600 177.700 ;
        RECT 119.600 177.600 120.400 177.700 ;
        RECT 134.000 177.600 134.800 177.700 ;
        RECT 244.400 178.300 245.200 178.400 ;
        RECT 271.600 178.300 272.400 178.400 ;
        RECT 314.800 178.300 315.600 178.400 ;
        RECT 244.400 177.700 267.500 178.300 ;
        RECT 244.400 177.600 245.200 177.700 ;
        RECT 266.900 176.400 267.500 177.700 ;
        RECT 271.600 177.700 315.600 178.300 ;
        RECT 271.600 177.600 272.400 177.700 ;
        RECT 314.800 177.600 315.600 177.700 ;
        RECT 322.800 178.300 323.600 178.400 ;
        RECT 342.000 178.300 342.800 178.400 ;
        RECT 322.800 177.700 342.800 178.300 ;
        RECT 322.800 177.600 323.600 177.700 ;
        RECT 342.000 177.600 342.800 177.700 ;
        RECT 350.000 178.300 350.800 178.400 ;
        RECT 354.800 178.300 355.600 178.400 ;
        RECT 350.000 177.700 355.600 178.300 ;
        RECT 350.000 177.600 350.800 177.700 ;
        RECT 354.800 177.600 355.600 177.700 ;
        RECT 359.600 178.300 360.400 178.400 ;
        RECT 362.800 178.300 363.600 178.400 ;
        RECT 359.600 177.700 363.600 178.300 ;
        RECT 359.600 177.600 360.400 177.700 ;
        RECT 362.800 177.600 363.600 177.700 ;
        RECT 367.600 178.300 368.400 178.400 ;
        RECT 370.800 178.300 371.600 178.400 ;
        RECT 367.600 177.700 371.600 178.300 ;
        RECT 367.600 177.600 368.400 177.700 ;
        RECT 370.800 177.600 371.600 177.700 ;
        RECT 391.600 178.300 392.400 178.400 ;
        RECT 401.200 178.300 402.000 178.400 ;
        RECT 446.000 178.300 446.800 178.400 ;
        RECT 391.600 177.700 446.800 178.300 ;
        RECT 391.600 177.600 392.400 177.700 ;
        RECT 401.200 177.600 402.000 177.700 ;
        RECT 446.000 177.600 446.800 177.700 ;
        RECT 4.400 176.300 5.200 176.400 ;
        RECT 9.200 176.300 10.000 176.400 ;
        RECT 4.400 175.700 10.000 176.300 ;
        RECT 4.400 175.600 5.200 175.700 ;
        RECT 9.200 175.600 10.000 175.700 ;
        RECT 10.800 176.300 11.600 176.400 ;
        RECT 22.000 176.300 22.800 176.400 ;
        RECT 38.000 176.300 38.800 176.400 ;
        RECT 10.800 175.700 38.800 176.300 ;
        RECT 10.800 175.600 11.600 175.700 ;
        RECT 22.000 175.600 22.800 175.700 ;
        RECT 38.000 175.600 38.800 175.700 ;
        RECT 42.800 176.300 43.600 176.400 ;
        RECT 76.400 176.300 77.200 176.400 ;
        RECT 42.800 175.700 77.200 176.300 ;
        RECT 42.800 175.600 43.600 175.700 ;
        RECT 76.400 175.600 77.200 175.700 ;
        RECT 86.000 176.300 86.800 176.400 ;
        RECT 90.800 176.300 91.600 176.400 ;
        RECT 86.000 175.700 91.600 176.300 ;
        RECT 86.000 175.600 86.800 175.700 ;
        RECT 90.800 175.600 91.600 175.700 ;
        RECT 164.400 176.300 165.200 176.400 ;
        RECT 193.200 176.300 194.000 176.400 ;
        RECT 164.400 175.700 194.000 176.300 ;
        RECT 164.400 175.600 165.200 175.700 ;
        RECT 193.200 175.600 194.000 175.700 ;
        RECT 199.600 176.300 200.400 176.400 ;
        RECT 228.400 176.300 229.200 176.400 ;
        RECT 199.600 175.700 229.200 176.300 ;
        RECT 199.600 175.600 200.400 175.700 ;
        RECT 228.400 175.600 229.200 175.700 ;
        RECT 244.400 176.300 245.200 176.400 ;
        RECT 247.600 176.300 248.400 176.400 ;
        RECT 244.400 175.700 248.400 176.300 ;
        RECT 244.400 175.600 245.200 175.700 ;
        RECT 247.600 175.600 248.400 175.700 ;
        RECT 266.800 176.300 267.600 176.400 ;
        RECT 290.800 176.300 291.600 176.400 ;
        RECT 266.800 175.700 291.600 176.300 ;
        RECT 266.800 175.600 267.600 175.700 ;
        RECT 290.800 175.600 291.600 175.700 ;
        RECT 303.600 176.300 304.400 176.400 ;
        RECT 334.000 176.300 334.800 176.400 ;
        RECT 303.600 175.700 334.800 176.300 ;
        RECT 303.600 175.600 304.400 175.700 ;
        RECT 334.000 175.600 334.800 175.700 ;
        RECT 348.400 176.300 349.200 176.400 ;
        RECT 353.200 176.300 354.000 176.400 ;
        RECT 348.400 175.700 354.000 176.300 ;
        RECT 348.400 175.600 349.200 175.700 ;
        RECT 353.200 175.600 354.000 175.700 ;
        RECT 460.400 176.300 461.200 176.400 ;
        RECT 468.400 176.300 469.200 176.400 ;
        RECT 460.400 175.700 469.200 176.300 ;
        RECT 460.400 175.600 461.200 175.700 ;
        RECT 468.400 175.600 469.200 175.700 ;
        RECT 470.000 176.300 470.800 176.400 ;
        RECT 486.000 176.300 486.800 176.400 ;
        RECT 470.000 175.700 486.800 176.300 ;
        RECT 470.000 175.600 470.800 175.700 ;
        RECT 486.000 175.600 486.800 175.700 ;
        RECT 497.200 176.300 498.000 176.400 ;
        RECT 502.000 176.300 502.800 176.400 ;
        RECT 497.200 175.700 502.800 176.300 ;
        RECT 497.200 175.600 498.000 175.700 ;
        RECT 502.000 175.600 502.800 175.700 ;
        RECT 20.400 174.300 21.200 174.400 ;
        RECT 30.000 174.300 30.800 174.400 ;
        RECT 20.400 173.700 30.800 174.300 ;
        RECT 20.400 173.600 21.200 173.700 ;
        RECT 30.000 173.600 30.800 173.700 ;
        RECT 36.400 174.300 37.200 174.400 ;
        RECT 42.800 174.300 43.600 174.400 ;
        RECT 36.400 173.700 43.600 174.300 ;
        RECT 36.400 173.600 37.200 173.700 ;
        RECT 42.800 173.600 43.600 173.700 ;
        RECT 94.000 174.300 94.800 174.400 ;
        RECT 100.400 174.300 101.200 174.400 ;
        RECT 94.000 173.700 101.200 174.300 ;
        RECT 94.000 173.600 94.800 173.700 ;
        RECT 100.400 173.600 101.200 173.700 ;
        RECT 105.200 174.300 106.000 174.400 ;
        RECT 137.200 174.300 138.000 174.400 ;
        RECT 105.200 173.700 138.000 174.300 ;
        RECT 105.200 173.600 106.000 173.700 ;
        RECT 137.200 173.600 138.000 173.700 ;
        RECT 178.800 174.300 179.600 174.400 ;
        RECT 186.800 174.300 187.600 174.400 ;
        RECT 178.800 173.700 187.600 174.300 ;
        RECT 178.800 173.600 179.600 173.700 ;
        RECT 186.800 173.600 187.600 173.700 ;
        RECT 222.000 174.300 222.800 174.400 ;
        RECT 238.000 174.300 238.800 174.400 ;
        RECT 222.000 173.700 238.800 174.300 ;
        RECT 222.000 173.600 222.800 173.700 ;
        RECT 238.000 173.600 238.800 173.700 ;
        RECT 246.000 174.300 246.800 174.400 ;
        RECT 257.200 174.300 258.000 174.400 ;
        RECT 246.000 173.700 258.000 174.300 ;
        RECT 246.000 173.600 246.800 173.700 ;
        RECT 257.200 173.600 258.000 173.700 ;
        RECT 265.200 174.300 266.000 174.400 ;
        RECT 273.200 174.300 274.000 174.400 ;
        RECT 265.200 173.700 274.000 174.300 ;
        RECT 265.200 173.600 266.000 173.700 ;
        RECT 273.200 173.600 274.000 173.700 ;
        RECT 282.800 174.300 283.600 174.400 ;
        RECT 289.200 174.300 290.000 174.400 ;
        RECT 282.800 173.700 290.000 174.300 ;
        RECT 282.800 173.600 283.600 173.700 ;
        RECT 289.200 173.600 290.000 173.700 ;
        RECT 302.000 174.300 302.800 174.400 ;
        RECT 356.400 174.300 357.200 174.400 ;
        RECT 302.000 173.700 357.200 174.300 ;
        RECT 302.000 173.600 302.800 173.700 ;
        RECT 356.400 173.600 357.200 173.700 ;
        RECT 401.200 174.300 402.000 174.400 ;
        RECT 404.400 174.300 405.200 174.400 ;
        RECT 401.200 173.700 405.200 174.300 ;
        RECT 401.200 173.600 402.000 173.700 ;
        RECT 404.400 173.600 405.200 173.700 ;
        RECT 463.600 174.300 464.400 174.400 ;
        RECT 471.600 174.300 472.400 174.400 ;
        RECT 463.600 173.700 472.400 174.300 ;
        RECT 463.600 173.600 464.400 173.700 ;
        RECT 471.600 173.600 472.400 173.700 ;
        RECT 478.000 174.300 478.800 174.400 ;
        RECT 502.000 174.300 502.800 174.400 ;
        RECT 505.200 174.300 506.000 174.400 ;
        RECT 478.000 173.700 506.000 174.300 ;
        RECT 478.000 173.600 478.800 173.700 ;
        RECT 502.000 173.600 502.800 173.700 ;
        RECT 505.200 173.600 506.000 173.700 ;
        RECT 506.800 174.300 507.600 174.400 ;
        RECT 513.200 174.300 514.000 174.400 ;
        RECT 506.800 173.700 514.000 174.300 ;
        RECT 506.800 173.600 507.600 173.700 ;
        RECT 513.200 173.600 514.000 173.700 ;
        RECT 9.200 172.300 10.000 172.400 ;
        RECT 33.200 172.300 34.000 172.400 ;
        RECT 46.000 172.300 46.800 172.400 ;
        RECT 9.200 171.700 46.800 172.300 ;
        RECT 9.200 171.600 10.000 171.700 ;
        RECT 33.200 171.600 34.000 171.700 ;
        RECT 46.000 171.600 46.800 171.700 ;
        RECT 97.200 172.300 98.000 172.400 ;
        RECT 106.800 172.300 107.600 172.400 ;
        RECT 97.200 171.700 107.600 172.300 ;
        RECT 97.200 171.600 98.000 171.700 ;
        RECT 106.800 171.600 107.600 171.700 ;
        RECT 164.400 172.300 165.200 172.400 ;
        RECT 167.600 172.300 168.400 172.400 ;
        RECT 218.800 172.300 219.600 172.400 ;
        RECT 238.000 172.300 238.800 172.400 ;
        RECT 164.400 171.700 238.800 172.300 ;
        RECT 164.400 171.600 165.200 171.700 ;
        RECT 167.600 171.600 168.400 171.700 ;
        RECT 218.800 171.600 219.600 171.700 ;
        RECT 238.000 171.600 238.800 171.700 ;
        RECT 241.200 172.300 242.000 172.400 ;
        RECT 252.400 172.300 253.200 172.400 ;
        RECT 241.200 171.700 253.200 172.300 ;
        RECT 241.200 171.600 242.000 171.700 ;
        RECT 252.400 171.600 253.200 171.700 ;
        RECT 262.000 172.300 262.800 172.400 ;
        RECT 270.000 172.300 270.800 172.400 ;
        RECT 284.400 172.300 285.200 172.400 ;
        RECT 262.000 171.700 285.200 172.300 ;
        RECT 262.000 171.600 262.800 171.700 ;
        RECT 270.000 171.600 270.800 171.700 ;
        RECT 284.400 171.600 285.200 171.700 ;
        RECT 406.000 172.300 406.800 172.400 ;
        RECT 410.800 172.300 411.600 172.400 ;
        RECT 406.000 171.700 411.600 172.300 ;
        RECT 406.000 171.600 406.800 171.700 ;
        RECT 410.800 171.600 411.600 171.700 ;
        RECT 505.200 172.300 506.000 172.400 ;
        RECT 510.000 172.300 510.800 172.400 ;
        RECT 505.200 171.700 510.800 172.300 ;
        RECT 505.200 171.600 506.000 171.700 ;
        RECT 510.000 171.600 510.800 171.700 ;
        RECT 522.800 172.300 523.600 172.400 ;
        RECT 526.000 172.300 526.800 172.400 ;
        RECT 522.800 171.700 526.800 172.300 ;
        RECT 522.800 171.600 523.600 171.700 ;
        RECT 526.000 171.600 526.800 171.700 ;
        RECT 15.600 170.300 16.400 170.400 ;
        RECT 49.200 170.300 50.000 170.400 ;
        RECT 15.600 169.700 50.000 170.300 ;
        RECT 15.600 169.600 16.400 169.700 ;
        RECT 49.200 169.600 50.000 169.700 ;
        RECT 146.800 170.300 147.600 170.400 ;
        RECT 153.200 170.300 154.000 170.400 ;
        RECT 146.800 169.700 154.000 170.300 ;
        RECT 146.800 169.600 147.600 169.700 ;
        RECT 153.200 169.600 154.000 169.700 ;
        RECT 196.400 170.300 197.200 170.400 ;
        RECT 199.600 170.300 200.400 170.400 ;
        RECT 241.300 170.300 241.900 171.600 ;
        RECT 196.400 169.700 241.900 170.300 ;
        RECT 250.800 170.300 251.600 170.400 ;
        RECT 257.200 170.300 258.000 170.400 ;
        RECT 250.800 169.700 258.000 170.300 ;
        RECT 196.400 169.600 197.200 169.700 ;
        RECT 199.600 169.600 200.400 169.700 ;
        RECT 250.800 169.600 251.600 169.700 ;
        RECT 257.200 169.600 258.000 169.700 ;
        RECT 287.600 170.300 288.400 170.400 ;
        RECT 292.400 170.300 293.200 170.400 ;
        RECT 287.600 169.700 293.200 170.300 ;
        RECT 287.600 169.600 288.400 169.700 ;
        RECT 292.400 169.600 293.200 169.700 ;
        RECT 308.400 170.300 309.200 170.400 ;
        RECT 329.200 170.300 330.000 170.400 ;
        RECT 308.400 169.700 330.000 170.300 ;
        RECT 308.400 169.600 309.200 169.700 ;
        RECT 329.200 169.600 330.000 169.700 ;
        RECT 42.800 167.600 43.600 168.400 ;
        RECT 87.600 168.300 88.400 168.400 ;
        RECT 95.600 168.300 96.400 168.400 ;
        RECT 87.600 167.700 96.400 168.300 ;
        RECT 87.600 167.600 88.400 167.700 ;
        RECT 95.600 167.600 96.400 167.700 ;
        RECT 230.000 168.300 230.800 168.400 ;
        RECT 265.200 168.300 266.000 168.400 ;
        RECT 286.000 168.300 286.800 168.400 ;
        RECT 230.000 167.700 286.800 168.300 ;
        RECT 230.000 167.600 230.800 167.700 ;
        RECT 265.200 167.600 266.000 167.700 ;
        RECT 286.000 167.600 286.800 167.700 ;
        RECT 398.000 168.300 398.800 168.400 ;
        RECT 402.800 168.300 403.600 168.400 ;
        RECT 398.000 167.700 403.600 168.300 ;
        RECT 398.000 167.600 398.800 167.700 ;
        RECT 402.800 167.600 403.600 167.700 ;
        RECT 479.600 168.300 480.400 168.400 ;
        RECT 484.400 168.300 485.200 168.400 ;
        RECT 479.600 167.700 485.200 168.300 ;
        RECT 479.600 167.600 480.400 167.700 ;
        RECT 484.400 167.600 485.200 167.700 ;
        RECT 486.000 168.300 486.800 168.400 ;
        RECT 489.200 168.300 490.000 168.400 ;
        RECT 494.000 168.300 494.800 168.400 ;
        RECT 486.000 167.700 494.800 168.300 ;
        RECT 486.000 167.600 486.800 167.700 ;
        RECT 489.200 167.600 490.000 167.700 ;
        RECT 494.000 167.600 494.800 167.700 ;
        RECT 30.000 166.300 30.800 166.400 ;
        RECT 41.200 166.300 42.000 166.400 ;
        RECT 30.000 165.700 42.000 166.300 ;
        RECT 30.000 165.600 30.800 165.700 ;
        RECT 41.200 165.600 42.000 165.700 ;
        RECT 234.800 166.300 235.600 166.400 ;
        RECT 258.800 166.300 259.600 166.400 ;
        RECT 234.800 165.700 259.600 166.300 ;
        RECT 234.800 165.600 235.600 165.700 ;
        RECT 258.800 165.600 259.600 165.700 ;
        RECT 334.000 166.300 334.800 166.400 ;
        RECT 398.000 166.300 398.800 166.400 ;
        RECT 466.800 166.300 467.600 166.400 ;
        RECT 334.000 165.700 397.100 166.300 ;
        RECT 334.000 165.600 334.800 165.700 ;
        RECT 28.400 164.300 29.200 164.400 ;
        RECT 34.800 164.300 35.600 164.400 ;
        RECT 58.800 164.300 59.600 164.400 ;
        RECT 28.400 163.700 59.600 164.300 ;
        RECT 28.400 163.600 29.200 163.700 ;
        RECT 34.800 163.600 35.600 163.700 ;
        RECT 58.800 163.600 59.600 163.700 ;
        RECT 218.800 164.300 219.600 164.400 ;
        RECT 236.400 164.300 237.200 164.400 ;
        RECT 218.800 163.700 237.200 164.300 ;
        RECT 218.800 163.600 219.600 163.700 ;
        RECT 236.400 163.600 237.200 163.700 ;
        RECT 238.000 164.300 238.800 164.400 ;
        RECT 311.600 164.300 312.400 164.400 ;
        RECT 238.000 163.700 312.400 164.300 ;
        RECT 396.500 164.300 397.100 165.700 ;
        RECT 398.000 165.700 467.600 166.300 ;
        RECT 398.000 165.600 398.800 165.700 ;
        RECT 466.800 165.600 467.600 165.700 ;
        RECT 468.400 166.300 469.200 166.400 ;
        RECT 474.800 166.300 475.600 166.400 ;
        RECT 468.400 165.700 475.600 166.300 ;
        RECT 468.400 165.600 469.200 165.700 ;
        RECT 474.800 165.600 475.600 165.700 ;
        RECT 497.200 165.600 498.000 166.400 ;
        RECT 503.600 166.300 504.400 166.400 ;
        RECT 510.000 166.300 510.800 166.400 ;
        RECT 503.600 165.700 510.800 166.300 ;
        RECT 503.600 165.600 504.400 165.700 ;
        RECT 510.000 165.600 510.800 165.700 ;
        RECT 399.600 164.300 400.400 164.400 ;
        RECT 396.500 163.700 400.400 164.300 ;
        RECT 238.000 163.600 238.800 163.700 ;
        RECT 311.600 163.600 312.400 163.700 ;
        RECT 399.600 163.600 400.400 163.700 ;
        RECT 407.600 164.300 408.400 164.400 ;
        RECT 502.000 164.300 502.800 164.400 ;
        RECT 508.400 164.300 509.200 164.400 ;
        RECT 407.600 163.700 459.500 164.300 ;
        RECT 407.600 163.600 408.400 163.700 ;
        RECT 44.400 162.300 45.200 162.400 ;
        RECT 57.200 162.300 58.000 162.400 ;
        RECT 90.800 162.300 91.600 162.400 ;
        RECT 44.400 161.700 91.600 162.300 ;
        RECT 44.400 161.600 45.200 161.700 ;
        RECT 57.200 161.600 58.000 161.700 ;
        RECT 90.800 161.600 91.600 161.700 ;
        RECT 220.400 162.300 221.200 162.400 ;
        RECT 242.800 162.300 243.600 162.400 ;
        RECT 246.000 162.300 246.800 162.400 ;
        RECT 220.400 161.700 246.800 162.300 ;
        RECT 220.400 161.600 221.200 161.700 ;
        RECT 242.800 161.600 243.600 161.700 ;
        RECT 246.000 161.600 246.800 161.700 ;
        RECT 390.000 162.300 390.800 162.400 ;
        RECT 396.400 162.300 397.200 162.400 ;
        RECT 390.000 161.700 397.200 162.300 ;
        RECT 458.900 162.300 459.500 163.700 ;
        RECT 502.000 163.700 509.200 164.300 ;
        RECT 502.000 163.600 502.800 163.700 ;
        RECT 508.400 163.600 509.200 163.700 ;
        RECT 511.600 162.300 512.400 162.400 ;
        RECT 458.900 161.700 512.400 162.300 ;
        RECT 390.000 161.600 390.800 161.700 ;
        RECT 396.400 161.600 397.200 161.700 ;
        RECT 511.600 161.600 512.400 161.700 ;
        RECT 49.200 159.600 50.000 160.400 ;
        RECT 356.400 160.300 357.200 160.400 ;
        RECT 406.000 160.300 406.800 160.400 ;
        RECT 356.400 159.700 406.800 160.300 ;
        RECT 356.400 159.600 357.200 159.700 ;
        RECT 406.000 159.600 406.800 159.700 ;
        RECT 452.400 160.300 453.200 160.400 ;
        RECT 462.000 160.300 462.800 160.400 ;
        RECT 452.400 159.700 462.800 160.300 ;
        RECT 452.400 159.600 453.200 159.700 ;
        RECT 462.000 159.600 462.800 159.700 ;
        RECT 465.200 160.300 466.000 160.400 ;
        RECT 495.600 160.300 496.400 160.400 ;
        RECT 465.200 159.700 496.400 160.300 ;
        RECT 465.200 159.600 466.000 159.700 ;
        RECT 495.600 159.600 496.400 159.700 ;
        RECT 4.400 158.300 5.200 158.400 ;
        RECT 119.600 158.300 120.400 158.400 ;
        RECT 4.400 157.700 120.400 158.300 ;
        RECT 4.400 157.600 5.200 157.700 ;
        RECT 119.600 157.600 120.400 157.700 ;
        RECT 239.600 158.300 240.400 158.400 ;
        RECT 241.200 158.300 242.000 158.400 ;
        RECT 290.800 158.300 291.600 158.400 ;
        RECT 239.600 157.700 291.600 158.300 ;
        RECT 239.600 157.600 240.400 157.700 ;
        RECT 241.200 157.600 242.000 157.700 ;
        RECT 290.800 157.600 291.600 157.700 ;
        RECT 351.600 158.300 352.400 158.400 ;
        RECT 372.400 158.300 373.200 158.400 ;
        RECT 351.600 157.700 373.200 158.300 ;
        RECT 351.600 157.600 352.400 157.700 ;
        RECT 372.400 157.600 373.200 157.700 ;
        RECT 380.400 158.300 381.200 158.400 ;
        RECT 398.000 158.300 398.800 158.400 ;
        RECT 463.600 158.300 464.400 158.400 ;
        RECT 481.200 158.300 482.000 158.400 ;
        RECT 380.400 157.700 398.800 158.300 ;
        RECT 380.400 157.600 381.200 157.700 ;
        RECT 398.000 157.600 398.800 157.700 ;
        RECT 415.700 157.700 482.000 158.300 ;
        RECT 42.800 156.300 43.600 156.400 ;
        RECT 63.600 156.300 64.400 156.400 ;
        RECT 42.800 155.700 64.400 156.300 ;
        RECT 42.800 155.600 43.600 155.700 ;
        RECT 63.600 155.600 64.400 155.700 ;
        RECT 103.600 156.300 104.400 156.400 ;
        RECT 108.400 156.300 109.200 156.400 ;
        RECT 103.600 155.700 109.200 156.300 ;
        RECT 103.600 155.600 104.400 155.700 ;
        RECT 108.400 155.600 109.200 155.700 ;
        RECT 110.000 156.300 110.800 156.400 ;
        RECT 121.200 156.300 122.000 156.400 ;
        RECT 145.200 156.300 146.000 156.400 ;
        RECT 110.000 155.700 146.000 156.300 ;
        RECT 110.000 155.600 110.800 155.700 ;
        RECT 121.200 155.600 122.000 155.700 ;
        RECT 145.200 155.600 146.000 155.700 ;
        RECT 337.200 156.300 338.000 156.400 ;
        RECT 375.600 156.300 376.400 156.400 ;
        RECT 337.200 155.700 376.400 156.300 ;
        RECT 337.200 155.600 338.000 155.700 ;
        RECT 375.600 155.600 376.400 155.700 ;
        RECT 378.800 156.300 379.600 156.400 ;
        RECT 415.700 156.300 416.300 157.700 ;
        RECT 463.600 157.600 464.400 157.700 ;
        RECT 481.200 157.600 482.000 157.700 ;
        RECT 378.800 155.700 416.300 156.300 ;
        RECT 417.200 156.300 418.000 156.400 ;
        RECT 433.200 156.300 434.000 156.400 ;
        RECT 458.800 156.300 459.600 156.400 ;
        RECT 487.600 156.300 488.400 156.400 ;
        RECT 417.200 155.700 488.400 156.300 ;
        RECT 378.800 155.600 379.600 155.700 ;
        RECT 417.200 155.600 418.000 155.700 ;
        RECT 433.200 155.600 434.000 155.700 ;
        RECT 458.800 155.600 459.600 155.700 ;
        RECT 487.600 155.600 488.400 155.700 ;
        RECT 7.600 154.300 8.400 154.400 ;
        RECT 25.200 154.300 26.000 154.400 ;
        RECT 7.600 153.700 26.000 154.300 ;
        RECT 7.600 153.600 8.400 153.700 ;
        RECT 25.200 153.600 26.000 153.700 ;
        RECT 36.400 154.300 37.200 154.400 ;
        RECT 42.800 154.300 43.600 154.400 ;
        RECT 44.400 154.300 45.200 154.400 ;
        RECT 36.400 153.700 45.200 154.300 ;
        RECT 36.400 153.600 37.200 153.700 ;
        RECT 42.800 153.600 43.600 153.700 ;
        RECT 44.400 153.600 45.200 153.700 ;
        RECT 50.800 154.300 51.600 154.400 ;
        RECT 60.400 154.300 61.200 154.400 ;
        RECT 50.800 153.700 61.200 154.300 ;
        RECT 50.800 153.600 51.600 153.700 ;
        RECT 60.400 153.600 61.200 153.700 ;
        RECT 81.200 154.300 82.000 154.400 ;
        RECT 114.800 154.300 115.600 154.400 ;
        RECT 81.200 153.700 115.600 154.300 ;
        RECT 81.200 153.600 82.000 153.700 ;
        RECT 114.800 153.600 115.600 153.700 ;
        RECT 255.600 154.300 256.400 154.400 ;
        RECT 271.600 154.300 272.400 154.400 ;
        RECT 279.600 154.300 280.400 154.400 ;
        RECT 255.600 153.700 280.400 154.300 ;
        RECT 255.600 153.600 256.400 153.700 ;
        RECT 271.600 153.600 272.400 153.700 ;
        RECT 279.600 153.600 280.400 153.700 ;
        RECT 334.000 154.300 334.800 154.400 ;
        RECT 369.200 154.300 370.000 154.400 ;
        RECT 334.000 153.700 370.000 154.300 ;
        RECT 334.000 153.600 334.800 153.700 ;
        RECT 369.200 153.600 370.000 153.700 ;
        RECT 394.800 154.300 395.600 154.400 ;
        RECT 398.000 154.300 398.800 154.400 ;
        RECT 404.400 154.300 405.200 154.400 ;
        RECT 394.800 153.700 405.200 154.300 ;
        RECT 394.800 153.600 395.600 153.700 ;
        RECT 398.000 153.600 398.800 153.700 ;
        RECT 404.400 153.600 405.200 153.700 ;
        RECT 407.600 154.300 408.400 154.400 ;
        RECT 455.600 154.300 456.400 154.400 ;
        RECT 407.600 153.700 456.400 154.300 ;
        RECT 407.600 153.600 408.400 153.700 ;
        RECT 455.600 153.600 456.400 153.700 ;
        RECT 463.600 154.300 464.400 154.400 ;
        RECT 487.600 154.300 488.400 154.400 ;
        RECT 494.000 154.300 494.800 154.400 ;
        RECT 463.600 153.700 472.300 154.300 ;
        RECT 463.600 153.600 464.400 153.700 ;
        RECT 471.700 152.400 472.300 153.700 ;
        RECT 487.600 153.700 494.800 154.300 ;
        RECT 487.600 153.600 488.400 153.700 ;
        RECT 494.000 153.600 494.800 153.700 ;
        RECT 498.800 154.300 499.600 154.400 ;
        RECT 506.800 154.300 507.600 154.400 ;
        RECT 511.600 154.300 512.400 154.400 ;
        RECT 498.800 153.700 512.400 154.300 ;
        RECT 498.800 153.600 499.600 153.700 ;
        RECT 506.800 153.600 507.600 153.700 ;
        RECT 511.600 153.600 512.400 153.700 ;
        RECT 516.400 154.300 517.200 154.400 ;
        RECT 519.600 154.300 520.400 154.400 ;
        RECT 516.400 153.700 520.400 154.300 ;
        RECT 516.400 153.600 517.200 153.700 ;
        RECT 519.600 153.600 520.400 153.700 ;
        RECT 2.800 152.300 3.600 152.400 ;
        RECT 4.400 152.300 5.200 152.400 ;
        RECT 6.000 152.300 6.800 152.400 ;
        RECT 2.800 151.700 6.800 152.300 ;
        RECT 2.800 151.600 3.600 151.700 ;
        RECT 4.400 151.600 5.200 151.700 ;
        RECT 6.000 151.600 6.800 151.700 ;
        RECT 14.000 152.300 14.800 152.400 ;
        RECT 18.800 152.300 19.600 152.400 ;
        RECT 36.400 152.300 37.200 152.400 ;
        RECT 14.000 151.700 37.200 152.300 ;
        RECT 14.000 151.600 14.800 151.700 ;
        RECT 18.800 151.600 19.600 151.700 ;
        RECT 36.400 151.600 37.200 151.700 ;
        RECT 52.400 152.300 53.200 152.400 ;
        RECT 65.200 152.300 66.000 152.400 ;
        RECT 102.000 152.300 102.800 152.400 ;
        RECT 106.800 152.300 107.600 152.400 ;
        RECT 52.400 151.700 107.600 152.300 ;
        RECT 52.400 151.600 53.200 151.700 ;
        RECT 65.200 151.600 66.000 151.700 ;
        RECT 102.000 151.600 102.800 151.700 ;
        RECT 106.800 151.600 107.600 151.700 ;
        RECT 183.600 152.300 184.400 152.400 ;
        RECT 188.400 152.300 189.200 152.400 ;
        RECT 183.600 151.700 189.200 152.300 ;
        RECT 183.600 151.600 184.400 151.700 ;
        RECT 188.400 151.600 189.200 151.700 ;
        RECT 201.200 152.300 202.000 152.400 ;
        RECT 215.600 152.300 216.400 152.400 ;
        RECT 303.600 152.300 304.400 152.400 ;
        RECT 201.200 151.700 304.400 152.300 ;
        RECT 201.200 151.600 202.000 151.700 ;
        RECT 215.600 151.600 216.400 151.700 ;
        RECT 303.600 151.600 304.400 151.700 ;
        RECT 329.200 152.300 330.000 152.400 ;
        RECT 340.400 152.300 341.200 152.400 ;
        RECT 329.200 151.700 341.200 152.300 ;
        RECT 329.200 151.600 330.000 151.700 ;
        RECT 340.400 151.600 341.200 151.700 ;
        RECT 345.200 152.300 346.000 152.400 ;
        RECT 351.600 152.300 352.400 152.400 ;
        RECT 362.800 152.300 363.600 152.400 ;
        RECT 345.200 151.700 363.600 152.300 ;
        RECT 345.200 151.600 346.000 151.700 ;
        RECT 351.600 151.600 352.400 151.700 ;
        RECT 362.800 151.600 363.600 151.700 ;
        RECT 370.800 152.300 371.600 152.400 ;
        RECT 382.000 152.300 382.800 152.400 ;
        RECT 388.400 152.300 389.200 152.400 ;
        RECT 370.800 151.700 389.200 152.300 ;
        RECT 370.800 151.600 371.600 151.700 ;
        RECT 382.000 151.600 382.800 151.700 ;
        RECT 388.400 151.600 389.200 151.700 ;
        RECT 396.400 152.300 397.200 152.400 ;
        RECT 409.200 152.300 410.000 152.400 ;
        RECT 396.400 151.700 410.000 152.300 ;
        RECT 396.400 151.600 397.200 151.700 ;
        RECT 409.200 151.600 410.000 151.700 ;
        RECT 414.000 152.300 414.800 152.400 ;
        RECT 423.600 152.300 424.400 152.400 ;
        RECT 414.000 151.700 424.400 152.300 ;
        RECT 414.000 151.600 414.800 151.700 ;
        RECT 423.600 151.600 424.400 151.700 ;
        RECT 446.000 152.300 446.800 152.400 ;
        RECT 454.000 152.300 454.800 152.400 ;
        RECT 446.000 151.700 454.800 152.300 ;
        RECT 446.000 151.600 446.800 151.700 ;
        RECT 454.000 151.600 454.800 151.700 ;
        RECT 471.600 152.300 472.400 152.400 ;
        RECT 479.600 152.300 480.400 152.400 ;
        RECT 508.400 152.300 509.200 152.400 ;
        RECT 471.600 151.700 480.400 152.300 ;
        RECT 471.600 151.600 472.400 151.700 ;
        RECT 479.600 151.600 480.400 151.700 ;
        RECT 487.700 151.700 509.200 152.300 ;
        RECT 487.700 150.400 488.300 151.700 ;
        RECT 508.400 151.600 509.200 151.700 ;
        RECT 510.000 152.300 510.800 152.400 ;
        RECT 545.200 152.300 546.000 152.400 ;
        RECT 510.000 151.700 546.000 152.300 ;
        RECT 510.000 151.600 510.800 151.700 ;
        RECT 545.200 151.600 546.000 151.700 ;
        RECT 7.600 150.300 8.400 150.400 ;
        RECT 17.200 150.300 18.000 150.400 ;
        RECT 28.400 150.300 29.200 150.400 ;
        RECT 7.600 149.700 29.200 150.300 ;
        RECT 7.600 149.600 8.400 149.700 ;
        RECT 17.200 149.600 18.000 149.700 ;
        RECT 28.400 149.600 29.200 149.700 ;
        RECT 119.600 150.300 120.400 150.400 ;
        RECT 135.600 150.300 136.400 150.400 ;
        RECT 119.600 149.700 136.400 150.300 ;
        RECT 119.600 149.600 120.400 149.700 ;
        RECT 135.600 149.600 136.400 149.700 ;
        RECT 175.600 150.300 176.400 150.400 ;
        RECT 193.200 150.300 194.000 150.400 ;
        RECT 204.400 150.300 205.200 150.400 ;
        RECT 207.600 150.300 208.400 150.400 ;
        RECT 175.600 149.700 208.400 150.300 ;
        RECT 175.600 149.600 176.400 149.700 ;
        RECT 193.200 149.600 194.000 149.700 ;
        RECT 204.400 149.600 205.200 149.700 ;
        RECT 207.600 149.600 208.400 149.700 ;
        RECT 222.000 150.300 222.800 150.400 ;
        RECT 225.200 150.300 226.000 150.400 ;
        RECT 222.000 149.700 226.000 150.300 ;
        RECT 222.000 149.600 222.800 149.700 ;
        RECT 225.200 149.600 226.000 149.700 ;
        RECT 260.400 150.300 261.200 150.400 ;
        RECT 270.000 150.300 270.800 150.400 ;
        RECT 281.200 150.300 282.000 150.400 ;
        RECT 260.400 149.700 282.000 150.300 ;
        RECT 260.400 149.600 261.200 149.700 ;
        RECT 270.000 149.600 270.800 149.700 ;
        RECT 281.200 149.600 282.000 149.700 ;
        RECT 295.600 150.300 296.400 150.400 ;
        RECT 337.200 150.300 338.000 150.400 ;
        RECT 295.600 149.700 338.000 150.300 ;
        RECT 295.600 149.600 296.400 149.700 ;
        RECT 337.200 149.600 338.000 149.700 ;
        RECT 343.600 150.300 344.400 150.400 ;
        RECT 350.000 150.300 350.800 150.400 ;
        RECT 353.200 150.300 354.000 150.400 ;
        RECT 356.400 150.300 357.200 150.400 ;
        RECT 343.600 149.700 357.200 150.300 ;
        RECT 343.600 149.600 344.400 149.700 ;
        RECT 350.000 149.600 350.800 149.700 ;
        RECT 353.200 149.600 354.000 149.700 ;
        RECT 356.400 149.600 357.200 149.700 ;
        RECT 367.600 150.300 368.400 150.400 ;
        RECT 378.800 150.300 379.600 150.400 ;
        RECT 367.600 149.700 379.600 150.300 ;
        RECT 367.600 149.600 368.400 149.700 ;
        RECT 378.800 149.600 379.600 149.700 ;
        RECT 383.600 150.300 384.400 150.400 ;
        RECT 386.800 150.300 387.600 150.400 ;
        RECT 383.600 149.700 387.600 150.300 ;
        RECT 383.600 149.600 384.400 149.700 ;
        RECT 386.800 149.600 387.600 149.700 ;
        RECT 393.200 150.300 394.000 150.400 ;
        RECT 401.200 150.300 402.000 150.400 ;
        RECT 407.600 150.300 408.400 150.400 ;
        RECT 393.200 149.700 408.400 150.300 ;
        RECT 393.200 149.600 394.000 149.700 ;
        RECT 401.200 149.600 402.000 149.700 ;
        RECT 407.600 149.600 408.400 149.700 ;
        RECT 417.200 150.300 418.000 150.400 ;
        RECT 425.200 150.300 426.000 150.400 ;
        RECT 417.200 149.700 426.000 150.300 ;
        RECT 417.200 149.600 418.000 149.700 ;
        RECT 425.200 149.600 426.000 149.700 ;
        RECT 452.400 150.300 453.200 150.400 ;
        RECT 455.600 150.300 456.400 150.400 ;
        RECT 452.400 149.700 456.400 150.300 ;
        RECT 452.400 149.600 453.200 149.700 ;
        RECT 455.600 149.600 456.400 149.700 ;
        RECT 468.400 150.300 469.200 150.400 ;
        RECT 487.600 150.300 488.400 150.400 ;
        RECT 468.400 149.700 488.400 150.300 ;
        RECT 468.400 149.600 469.200 149.700 ;
        RECT 487.600 149.600 488.400 149.700 ;
        RECT 500.400 150.300 501.200 150.400 ;
        RECT 503.600 150.300 504.400 150.400 ;
        RECT 516.400 150.300 517.200 150.400 ;
        RECT 500.400 149.700 517.200 150.300 ;
        RECT 500.400 149.600 501.200 149.700 ;
        RECT 503.600 149.600 504.400 149.700 ;
        RECT 516.400 149.600 517.200 149.700 ;
        RECT 39.600 148.300 40.400 148.400 ;
        RECT 41.200 148.300 42.000 148.400 ;
        RECT 39.600 147.700 42.000 148.300 ;
        RECT 39.600 147.600 40.400 147.700 ;
        RECT 41.200 147.600 42.000 147.700 ;
        RECT 58.800 148.300 59.600 148.400 ;
        RECT 62.000 148.300 62.800 148.400 ;
        RECT 58.800 147.700 62.800 148.300 ;
        RECT 58.800 147.600 59.600 147.700 ;
        RECT 62.000 147.600 62.800 147.700 ;
        RECT 65.200 148.300 66.000 148.400 ;
        RECT 90.800 148.300 91.600 148.400 ;
        RECT 65.200 147.700 91.600 148.300 ;
        RECT 65.200 147.600 66.000 147.700 ;
        RECT 90.800 147.600 91.600 147.700 ;
        RECT 161.200 148.300 162.000 148.400 ;
        RECT 193.200 148.300 194.000 148.400 ;
        RECT 161.200 147.700 194.000 148.300 ;
        RECT 161.200 147.600 162.000 147.700 ;
        RECT 193.200 147.600 194.000 147.700 ;
        RECT 196.400 148.300 197.200 148.400 ;
        RECT 206.000 148.300 206.800 148.400 ;
        RECT 215.600 148.300 216.400 148.400 ;
        RECT 196.400 147.700 216.400 148.300 ;
        RECT 196.400 147.600 197.200 147.700 ;
        RECT 206.000 147.600 206.800 147.700 ;
        RECT 215.600 147.600 216.400 147.700 ;
        RECT 234.800 148.300 235.600 148.400 ;
        RECT 262.000 148.300 262.800 148.400 ;
        RECT 234.800 147.700 262.800 148.300 ;
        RECT 234.800 147.600 235.600 147.700 ;
        RECT 262.000 147.600 262.800 147.700 ;
        RECT 266.800 148.300 267.600 148.400 ;
        RECT 287.600 148.300 288.400 148.400 ;
        RECT 266.800 147.700 288.400 148.300 ;
        RECT 266.800 147.600 267.600 147.700 ;
        RECT 287.600 147.600 288.400 147.700 ;
        RECT 314.800 148.300 315.600 148.400 ;
        RECT 329.200 148.300 330.000 148.400 ;
        RECT 314.800 147.700 330.000 148.300 ;
        RECT 314.800 147.600 315.600 147.700 ;
        RECT 329.200 147.600 330.000 147.700 ;
        RECT 386.800 148.300 387.600 148.400 ;
        RECT 401.200 148.300 402.000 148.400 ;
        RECT 418.800 148.300 419.600 148.400 ;
        RECT 386.800 147.700 419.600 148.300 ;
        RECT 386.800 147.600 387.600 147.700 ;
        RECT 401.200 147.600 402.000 147.700 ;
        RECT 418.800 147.600 419.600 147.700 ;
        RECT 452.400 148.300 453.200 148.400 ;
        RECT 510.000 148.300 510.800 148.400 ;
        RECT 452.400 147.700 510.800 148.300 ;
        RECT 452.400 147.600 453.200 147.700 ;
        RECT 510.000 147.600 510.800 147.700 ;
        RECT 511.600 148.300 512.400 148.400 ;
        RECT 518.000 148.300 518.800 148.400 ;
        RECT 511.600 147.700 518.800 148.300 ;
        RECT 511.600 147.600 512.400 147.700 ;
        RECT 518.000 147.600 518.800 147.700 ;
        RECT 20.400 145.600 21.200 146.400 ;
        RECT 31.600 146.300 32.400 146.400 ;
        RECT 39.600 146.300 40.400 146.400 ;
        RECT 50.800 146.300 51.600 146.400 ;
        RECT 31.600 145.700 51.600 146.300 ;
        RECT 31.600 145.600 32.400 145.700 ;
        RECT 39.600 145.600 40.400 145.700 ;
        RECT 50.800 145.600 51.600 145.700 ;
        RECT 66.800 146.300 67.600 146.400 ;
        RECT 73.200 146.300 74.000 146.400 ;
        RECT 87.600 146.300 88.400 146.400 ;
        RECT 66.800 145.700 88.400 146.300 ;
        RECT 66.800 145.600 67.600 145.700 ;
        RECT 73.200 145.600 74.000 145.700 ;
        RECT 87.600 145.600 88.400 145.700 ;
        RECT 116.400 146.300 117.200 146.400 ;
        RECT 118.000 146.300 118.800 146.400 ;
        RECT 116.400 145.700 118.800 146.300 ;
        RECT 116.400 145.600 117.200 145.700 ;
        RECT 118.000 145.600 118.800 145.700 ;
        RECT 172.400 146.300 173.200 146.400 ;
        RECT 194.800 146.300 195.600 146.400 ;
        RECT 172.400 145.700 195.600 146.300 ;
        RECT 172.400 145.600 173.200 145.700 ;
        RECT 194.800 145.600 195.600 145.700 ;
        RECT 202.800 146.300 203.600 146.400 ;
        RECT 207.600 146.300 208.400 146.400 ;
        RECT 210.800 146.300 211.600 146.400 ;
        RECT 202.800 145.700 211.600 146.300 ;
        RECT 202.800 145.600 203.600 145.700 ;
        RECT 207.600 145.600 208.400 145.700 ;
        RECT 210.800 145.600 211.600 145.700 ;
        RECT 262.000 146.300 262.800 146.400 ;
        RECT 263.600 146.300 264.400 146.400 ;
        RECT 266.800 146.300 267.600 146.400 ;
        RECT 330.800 146.300 331.600 146.400 ;
        RECT 262.000 145.700 331.600 146.300 ;
        RECT 262.000 145.600 262.800 145.700 ;
        RECT 263.600 145.600 264.400 145.700 ;
        RECT 266.800 145.600 267.600 145.700 ;
        RECT 330.800 145.600 331.600 145.700 ;
        RECT 375.600 146.300 376.400 146.400 ;
        RECT 383.600 146.300 384.400 146.400 ;
        RECT 375.600 145.700 384.400 146.300 ;
        RECT 375.600 145.600 376.400 145.700 ;
        RECT 383.600 145.600 384.400 145.700 ;
        RECT 393.200 146.300 394.000 146.400 ;
        RECT 412.400 146.300 413.200 146.400 ;
        RECT 454.000 146.300 454.800 146.400 ;
        RECT 462.000 146.300 462.800 146.400 ;
        RECT 393.200 145.700 462.800 146.300 ;
        RECT 393.200 145.600 394.000 145.700 ;
        RECT 412.400 145.600 413.200 145.700 ;
        RECT 454.000 145.600 454.800 145.700 ;
        RECT 462.000 145.600 462.800 145.700 ;
        RECT 486.000 146.300 486.800 146.400 ;
        RECT 489.200 146.300 490.000 146.400 ;
        RECT 486.000 145.700 490.000 146.300 ;
        RECT 486.000 145.600 486.800 145.700 ;
        RECT 489.200 145.600 490.000 145.700 ;
        RECT 490.800 146.300 491.600 146.400 ;
        RECT 497.200 146.300 498.000 146.400 ;
        RECT 490.800 145.700 498.000 146.300 ;
        RECT 490.800 145.600 491.600 145.700 ;
        RECT 497.200 145.600 498.000 145.700 ;
        RECT 514.800 146.300 515.600 146.400 ;
        RECT 524.400 146.300 525.200 146.400 ;
        RECT 514.800 145.700 525.200 146.300 ;
        RECT 514.800 145.600 515.600 145.700 ;
        RECT 524.400 145.600 525.200 145.700 ;
        RECT 97.200 144.300 98.000 144.400 ;
        RECT 116.400 144.300 117.200 144.400 ;
        RECT 97.200 143.700 117.200 144.300 ;
        RECT 97.200 143.600 98.000 143.700 ;
        RECT 116.400 143.600 117.200 143.700 ;
        RECT 143.600 144.300 144.400 144.400 ;
        RECT 146.800 144.300 147.600 144.400 ;
        RECT 143.600 143.700 147.600 144.300 ;
        RECT 143.600 143.600 144.400 143.700 ;
        RECT 146.800 143.600 147.600 143.700 ;
        RECT 161.200 144.300 162.000 144.400 ;
        RECT 180.400 144.300 181.200 144.400 ;
        RECT 161.200 143.700 181.200 144.300 ;
        RECT 161.200 143.600 162.000 143.700 ;
        RECT 180.400 143.600 181.200 143.700 ;
        RECT 321.200 144.300 322.000 144.400 ;
        RECT 343.600 144.300 344.400 144.400 ;
        RECT 321.200 143.700 344.400 144.300 ;
        RECT 321.200 143.600 322.000 143.700 ;
        RECT 343.600 143.600 344.400 143.700 ;
        RECT 396.400 144.300 397.200 144.400 ;
        RECT 401.200 144.300 402.000 144.400 ;
        RECT 415.600 144.300 416.400 144.400 ;
        RECT 396.400 143.700 416.400 144.300 ;
        RECT 396.400 143.600 397.200 143.700 ;
        RECT 401.200 143.600 402.000 143.700 ;
        RECT 415.600 143.600 416.400 143.700 ;
        RECT 417.200 144.300 418.000 144.400 ;
        RECT 420.400 144.300 421.200 144.400 ;
        RECT 417.200 143.700 421.200 144.300 ;
        RECT 417.200 143.600 418.000 143.700 ;
        RECT 420.400 143.600 421.200 143.700 ;
        RECT 450.800 144.300 451.600 144.400 ;
        RECT 530.800 144.300 531.600 144.400 ;
        RECT 450.800 143.700 531.600 144.300 ;
        RECT 450.800 143.600 451.600 143.700 ;
        RECT 530.800 143.600 531.600 143.700 ;
        RECT 12.400 142.300 13.200 142.400 ;
        RECT 28.400 142.300 29.200 142.400 ;
        RECT 71.600 142.300 72.400 142.400 ;
        RECT 12.400 141.700 72.400 142.300 ;
        RECT 12.400 141.600 13.200 141.700 ;
        RECT 28.400 141.600 29.200 141.700 ;
        RECT 71.600 141.600 72.400 141.700 ;
        RECT 89.200 142.300 90.000 142.400 ;
        RECT 98.800 142.300 99.600 142.400 ;
        RECT 105.200 142.300 106.000 142.400 ;
        RECT 89.200 141.700 106.000 142.300 ;
        RECT 89.200 141.600 90.000 141.700 ;
        RECT 98.800 141.600 99.600 141.700 ;
        RECT 105.200 141.600 106.000 141.700 ;
        RECT 233.200 142.300 234.000 142.400 ;
        RECT 249.200 142.300 250.000 142.400 ;
        RECT 233.200 141.700 250.000 142.300 ;
        RECT 233.200 141.600 234.000 141.700 ;
        RECT 249.200 141.600 250.000 141.700 ;
        RECT 310.000 142.300 310.800 142.400 ;
        RECT 332.400 142.300 333.200 142.400 ;
        RECT 338.800 142.300 339.600 142.400 ;
        RECT 310.000 141.700 339.600 142.300 ;
        RECT 310.000 141.600 310.800 141.700 ;
        RECT 332.400 141.600 333.200 141.700 ;
        RECT 338.800 141.600 339.600 141.700 ;
        RECT 370.800 142.300 371.600 142.400 ;
        RECT 454.000 142.300 454.800 142.400 ;
        RECT 370.800 141.700 454.800 142.300 ;
        RECT 370.800 141.600 371.600 141.700 ;
        RECT 454.000 141.600 454.800 141.700 ;
        RECT 463.600 142.300 464.400 142.400 ;
        RECT 474.800 142.300 475.600 142.400 ;
        RECT 463.600 141.700 475.600 142.300 ;
        RECT 463.600 141.600 464.400 141.700 ;
        RECT 474.800 141.600 475.600 141.700 ;
        RECT 478.000 142.300 478.800 142.400 ;
        RECT 482.800 142.300 483.600 142.400 ;
        RECT 478.000 141.700 483.600 142.300 ;
        RECT 478.000 141.600 478.800 141.700 ;
        RECT 482.800 141.600 483.600 141.700 ;
        RECT 503.600 142.300 504.400 142.400 ;
        RECT 535.600 142.300 536.400 142.400 ;
        RECT 503.600 141.700 536.400 142.300 ;
        RECT 503.600 141.600 504.400 141.700 ;
        RECT 535.600 141.600 536.400 141.700 ;
        RECT 20.400 140.300 21.200 140.400 ;
        RECT 23.600 140.300 24.400 140.400 ;
        RECT 20.400 139.700 24.400 140.300 ;
        RECT 20.400 139.600 21.200 139.700 ;
        RECT 23.600 139.600 24.400 139.700 ;
        RECT 100.400 140.300 101.200 140.400 ;
        RECT 102.000 140.300 102.800 140.400 ;
        RECT 100.400 139.700 102.800 140.300 ;
        RECT 100.400 139.600 101.200 139.700 ;
        RECT 102.000 139.600 102.800 139.700 ;
        RECT 228.400 140.300 229.200 140.400 ;
        RECT 250.800 140.300 251.600 140.400 ;
        RECT 228.400 139.700 251.600 140.300 ;
        RECT 228.400 139.600 229.200 139.700 ;
        RECT 250.800 139.600 251.600 139.700 ;
        RECT 318.000 140.300 318.800 140.400 ;
        RECT 345.200 140.300 346.000 140.400 ;
        RECT 318.000 139.700 346.000 140.300 ;
        RECT 318.000 139.600 318.800 139.700 ;
        RECT 345.200 139.600 346.000 139.700 ;
        RECT 374.000 140.300 374.800 140.400 ;
        RECT 442.800 140.300 443.600 140.400 ;
        RECT 374.000 139.700 443.600 140.300 ;
        RECT 374.000 139.600 374.800 139.700 ;
        RECT 442.800 139.600 443.600 139.700 ;
        RECT 481.200 140.300 482.000 140.400 ;
        RECT 489.200 140.300 490.000 140.400 ;
        RECT 481.200 139.700 490.000 140.300 ;
        RECT 481.200 139.600 482.000 139.700 ;
        RECT 489.200 139.600 490.000 139.700 ;
        RECT 532.400 140.300 533.200 140.400 ;
        RECT 534.000 140.300 534.800 140.400 ;
        RECT 532.400 139.700 534.800 140.300 ;
        RECT 532.400 139.600 533.200 139.700 ;
        RECT 534.000 139.600 534.800 139.700 ;
        RECT 2.800 138.300 3.600 138.400 ;
        RECT 7.600 138.300 8.400 138.400 ;
        RECT 33.200 138.300 34.000 138.400 ;
        RECT 441.200 138.300 442.000 138.400 ;
        RECT 2.800 137.700 34.000 138.300 ;
        RECT 2.800 137.600 3.600 137.700 ;
        RECT 7.600 137.600 8.400 137.700 ;
        RECT 33.200 137.600 34.000 137.700 ;
        RECT 314.900 137.700 442.000 138.300 ;
        RECT 314.900 136.400 315.500 137.700 ;
        RECT 441.200 137.600 442.000 137.700 ;
        RECT 7.600 136.300 8.400 136.400 ;
        RECT 15.600 136.300 16.400 136.400 ;
        RECT 36.400 136.300 37.200 136.400 ;
        RECT 7.600 135.700 37.200 136.300 ;
        RECT 7.600 135.600 8.400 135.700 ;
        RECT 15.600 135.600 16.400 135.700 ;
        RECT 36.400 135.600 37.200 135.700 ;
        RECT 78.000 136.300 78.800 136.400 ;
        RECT 84.400 136.300 85.200 136.400 ;
        RECT 92.400 136.300 93.200 136.400 ;
        RECT 111.600 136.300 112.400 136.400 ;
        RECT 78.000 135.700 112.400 136.300 ;
        RECT 78.000 135.600 78.800 135.700 ;
        RECT 84.400 135.600 85.200 135.700 ;
        RECT 92.400 135.600 93.200 135.700 ;
        RECT 111.600 135.600 112.400 135.700 ;
        RECT 114.800 136.300 115.600 136.400 ;
        RECT 134.000 136.300 134.800 136.400 ;
        RECT 114.800 135.700 134.800 136.300 ;
        RECT 114.800 135.600 115.600 135.700 ;
        RECT 134.000 135.600 134.800 135.700 ;
        RECT 142.000 136.300 142.800 136.400 ;
        RECT 145.200 136.300 146.000 136.400 ;
        RECT 142.000 135.700 146.000 136.300 ;
        RECT 142.000 135.600 142.800 135.700 ;
        RECT 145.200 135.600 146.000 135.700 ;
        RECT 241.200 136.300 242.000 136.400 ;
        RECT 242.800 136.300 243.600 136.400 ;
        RECT 241.200 135.700 243.600 136.300 ;
        RECT 241.200 135.600 242.000 135.700 ;
        RECT 242.800 135.600 243.600 135.700 ;
        RECT 246.000 136.300 246.800 136.400 ;
        RECT 252.400 136.300 253.200 136.400 ;
        RECT 246.000 135.700 253.200 136.300 ;
        RECT 246.000 135.600 246.800 135.700 ;
        RECT 252.400 135.600 253.200 135.700 ;
        RECT 257.200 136.300 258.000 136.400 ;
        RECT 273.200 136.300 274.000 136.400 ;
        RECT 314.800 136.300 315.600 136.400 ;
        RECT 257.200 135.700 315.600 136.300 ;
        RECT 257.200 135.600 258.000 135.700 ;
        RECT 273.200 135.600 274.000 135.700 ;
        RECT 314.800 135.600 315.600 135.700 ;
        RECT 356.400 136.300 357.200 136.400 ;
        RECT 361.200 136.300 362.000 136.400 ;
        RECT 356.400 135.700 362.000 136.300 ;
        RECT 356.400 135.600 357.200 135.700 ;
        RECT 361.200 135.600 362.000 135.700 ;
        RECT 362.800 136.300 363.600 136.400 ;
        RECT 370.800 136.300 371.600 136.400 ;
        RECT 362.800 135.700 371.600 136.300 ;
        RECT 362.800 135.600 363.600 135.700 ;
        RECT 370.800 135.600 371.600 135.700 ;
        RECT 372.400 136.300 373.200 136.400 ;
        RECT 385.200 136.300 386.000 136.400 ;
        RECT 372.400 135.700 386.000 136.300 ;
        RECT 372.400 135.600 373.200 135.700 ;
        RECT 385.200 135.600 386.000 135.700 ;
        RECT 412.400 136.300 413.200 136.400 ;
        RECT 426.800 136.300 427.600 136.400 ;
        RECT 481.200 136.300 482.000 136.400 ;
        RECT 412.400 135.700 482.000 136.300 ;
        RECT 412.400 135.600 413.200 135.700 ;
        RECT 426.800 135.600 427.600 135.700 ;
        RECT 481.200 135.600 482.000 135.700 ;
        RECT 6.000 134.300 6.800 134.400 ;
        RECT 18.800 134.300 19.600 134.400 ;
        RECT 33.200 134.300 34.000 134.400 ;
        RECT 6.000 133.700 34.000 134.300 ;
        RECT 6.000 133.600 6.800 133.700 ;
        RECT 18.800 133.600 19.600 133.700 ;
        RECT 33.200 133.600 34.000 133.700 ;
        RECT 41.200 134.300 42.000 134.400 ;
        RECT 70.000 134.300 70.800 134.400 ;
        RECT 41.200 133.700 70.800 134.300 ;
        RECT 41.200 133.600 42.000 133.700 ;
        RECT 70.000 133.600 70.800 133.700 ;
        RECT 122.800 134.300 123.600 134.400 ;
        RECT 151.600 134.300 152.400 134.400 ;
        RECT 122.800 133.700 152.400 134.300 ;
        RECT 122.800 133.600 123.600 133.700 ;
        RECT 151.600 133.600 152.400 133.700 ;
        RECT 161.200 134.300 162.000 134.400 ;
        RECT 166.000 134.300 166.800 134.400 ;
        RECT 161.200 133.700 166.800 134.300 ;
        RECT 161.200 133.600 162.000 133.700 ;
        RECT 166.000 133.600 166.800 133.700 ;
        RECT 167.600 134.300 168.400 134.400 ;
        RECT 172.400 134.300 173.200 134.400 ;
        RECT 167.600 133.700 173.200 134.300 ;
        RECT 167.600 133.600 168.400 133.700 ;
        RECT 172.400 133.600 173.200 133.700 ;
        RECT 202.800 134.300 203.600 134.400 ;
        RECT 218.800 134.300 219.600 134.400 ;
        RECT 202.800 133.700 219.600 134.300 ;
        RECT 202.800 133.600 203.600 133.700 ;
        RECT 218.800 133.600 219.600 133.700 ;
        RECT 226.800 134.300 227.600 134.400 ;
        RECT 231.600 134.300 232.400 134.400 ;
        RECT 226.800 133.700 232.400 134.300 ;
        RECT 226.800 133.600 227.600 133.700 ;
        RECT 231.600 133.600 232.400 133.700 ;
        RECT 238.000 134.300 238.800 134.400 ;
        RECT 249.200 134.300 250.000 134.400 ;
        RECT 252.400 134.300 253.200 134.400 ;
        RECT 260.400 134.300 261.200 134.400 ;
        RECT 238.000 133.700 261.200 134.300 ;
        RECT 238.000 133.600 238.800 133.700 ;
        RECT 249.200 133.600 250.000 133.700 ;
        RECT 252.400 133.600 253.200 133.700 ;
        RECT 260.400 133.600 261.200 133.700 ;
        RECT 292.400 134.300 293.200 134.400 ;
        RECT 306.800 134.300 307.600 134.400 ;
        RECT 292.400 133.700 307.600 134.300 ;
        RECT 292.400 133.600 293.200 133.700 ;
        RECT 306.800 133.600 307.600 133.700 ;
        RECT 361.200 134.300 362.000 134.400 ;
        RECT 364.400 134.300 365.200 134.400 ;
        RECT 361.200 133.700 365.200 134.300 ;
        RECT 361.200 133.600 362.000 133.700 ;
        RECT 364.400 133.600 365.200 133.700 ;
        RECT 366.000 134.300 366.800 134.400 ;
        RECT 375.600 134.300 376.400 134.400 ;
        RECT 394.800 134.300 395.600 134.400 ;
        RECT 366.000 133.700 395.600 134.300 ;
        RECT 366.000 133.600 366.800 133.700 ;
        RECT 375.600 133.600 376.400 133.700 ;
        RECT 394.800 133.600 395.600 133.700 ;
        RECT 412.400 134.300 413.200 134.400 ;
        RECT 422.000 134.300 422.800 134.400 ;
        RECT 412.400 133.700 422.800 134.300 ;
        RECT 412.400 133.600 413.200 133.700 ;
        RECT 422.000 133.600 422.800 133.700 ;
        RECT 442.800 134.300 443.600 134.400 ;
        RECT 470.000 134.300 470.800 134.400 ;
        RECT 442.800 133.700 470.800 134.300 ;
        RECT 442.800 133.600 443.600 133.700 ;
        RECT 470.000 133.600 470.800 133.700 ;
        RECT 4.400 132.300 5.200 132.400 ;
        RECT 9.200 132.300 10.000 132.400 ;
        RECT 4.400 131.700 10.000 132.300 ;
        RECT 4.400 131.600 5.200 131.700 ;
        RECT 9.200 131.600 10.000 131.700 ;
        RECT 17.200 132.300 18.000 132.400 ;
        RECT 26.800 132.300 27.600 132.400 ;
        RECT 17.200 131.700 27.600 132.300 ;
        RECT 17.200 131.600 18.000 131.700 ;
        RECT 26.800 131.600 27.600 131.700 ;
        RECT 28.400 132.300 29.200 132.400 ;
        RECT 34.800 132.300 35.600 132.400 ;
        RECT 97.200 132.300 98.000 132.400 ;
        RECT 111.600 132.300 112.400 132.400 ;
        RECT 28.400 131.700 48.300 132.300 ;
        RECT 28.400 131.600 29.200 131.700 ;
        RECT 34.800 131.600 35.600 131.700 ;
        RECT 47.700 130.400 48.300 131.700 ;
        RECT 97.200 131.700 112.400 132.300 ;
        RECT 97.200 131.600 98.000 131.700 ;
        RECT 111.600 131.600 112.400 131.700 ;
        RECT 159.600 132.300 160.400 132.400 ;
        RECT 162.800 132.300 163.600 132.400 ;
        RECT 183.600 132.300 184.400 132.400 ;
        RECT 217.200 132.300 218.000 132.400 ;
        RECT 159.600 131.700 218.000 132.300 ;
        RECT 159.600 131.600 160.400 131.700 ;
        RECT 162.800 131.600 163.600 131.700 ;
        RECT 183.600 131.600 184.400 131.700 ;
        RECT 217.200 131.600 218.000 131.700 ;
        RECT 230.000 132.300 230.800 132.400 ;
        RECT 233.200 132.300 234.000 132.400 ;
        RECT 230.000 131.700 234.000 132.300 ;
        RECT 230.000 131.600 230.800 131.700 ;
        RECT 233.200 131.600 234.000 131.700 ;
        RECT 254.000 132.300 254.800 132.400 ;
        RECT 263.600 132.300 264.400 132.400 ;
        RECT 254.000 131.700 264.400 132.300 ;
        RECT 254.000 131.600 254.800 131.700 ;
        RECT 263.600 131.600 264.400 131.700 ;
        RECT 310.000 132.300 310.800 132.400 ;
        RECT 314.800 132.300 315.600 132.400 ;
        RECT 310.000 131.700 315.600 132.300 ;
        RECT 310.000 131.600 310.800 131.700 ;
        RECT 314.800 131.600 315.600 131.700 ;
        RECT 335.600 132.300 336.400 132.400 ;
        RECT 367.600 132.300 368.400 132.400 ;
        RECT 335.600 131.700 368.400 132.300 ;
        RECT 335.600 131.600 336.400 131.700 ;
        RECT 367.600 131.600 368.400 131.700 ;
        RECT 382.000 132.300 382.800 132.400 ;
        RECT 439.600 132.300 440.400 132.400 ;
        RECT 455.600 132.300 456.400 132.400 ;
        RECT 382.000 131.700 456.400 132.300 ;
        RECT 382.000 131.600 382.800 131.700 ;
        RECT 439.600 131.600 440.400 131.700 ;
        RECT 455.600 131.600 456.400 131.700 ;
        RECT 500.400 132.300 501.200 132.400 ;
        RECT 506.800 132.300 507.600 132.400 ;
        RECT 500.400 131.700 507.600 132.300 ;
        RECT 500.400 131.600 501.200 131.700 ;
        RECT 506.800 131.600 507.600 131.700 ;
        RECT 38.000 130.300 38.800 130.400 ;
        RECT 44.400 130.300 45.200 130.400 ;
        RECT 38.000 129.700 45.200 130.300 ;
        RECT 38.000 129.600 38.800 129.700 ;
        RECT 44.400 129.600 45.200 129.700 ;
        RECT 47.600 130.300 48.400 130.400 ;
        RECT 58.800 130.300 59.600 130.400 ;
        RECT 86.000 130.300 86.800 130.400 ;
        RECT 47.600 129.700 86.800 130.300 ;
        RECT 47.600 129.600 48.400 129.700 ;
        RECT 58.800 129.600 59.600 129.700 ;
        RECT 86.000 129.600 86.800 129.700 ;
        RECT 156.400 130.300 157.200 130.400 ;
        RECT 169.200 130.300 170.000 130.400 ;
        RECT 156.400 129.700 170.000 130.300 ;
        RECT 156.400 129.600 157.200 129.700 ;
        RECT 169.200 129.600 170.000 129.700 ;
        RECT 172.400 130.300 173.200 130.400 ;
        RECT 178.800 130.300 179.600 130.400 ;
        RECT 193.200 130.300 194.000 130.400 ;
        RECT 220.400 130.300 221.200 130.400 ;
        RECT 222.000 130.300 222.800 130.400 ;
        RECT 233.200 130.300 234.000 130.400 ;
        RECT 172.400 129.700 234.000 130.300 ;
        RECT 172.400 129.600 173.200 129.700 ;
        RECT 178.800 129.600 179.600 129.700 ;
        RECT 193.200 129.600 194.000 129.700 ;
        RECT 220.400 129.600 221.200 129.700 ;
        RECT 222.000 129.600 222.800 129.700 ;
        RECT 233.200 129.600 234.000 129.700 ;
        RECT 249.200 130.300 250.000 130.400 ;
        RECT 260.400 130.300 261.200 130.400 ;
        RECT 249.200 129.700 261.200 130.300 ;
        RECT 249.200 129.600 250.000 129.700 ;
        RECT 260.400 129.600 261.200 129.700 ;
        RECT 306.800 130.300 307.600 130.400 ;
        RECT 316.400 130.300 317.200 130.400 ;
        RECT 306.800 129.700 317.200 130.300 ;
        RECT 306.800 129.600 307.600 129.700 ;
        RECT 316.400 129.600 317.200 129.700 ;
        RECT 410.800 130.300 411.600 130.400 ;
        RECT 436.400 130.300 437.200 130.400 ;
        RECT 410.800 129.700 437.200 130.300 ;
        RECT 410.800 129.600 411.600 129.700 ;
        RECT 436.400 129.600 437.200 129.700 ;
        RECT 449.200 130.300 450.000 130.400 ;
        RECT 481.200 130.300 482.000 130.400 ;
        RECT 449.200 129.700 482.000 130.300 ;
        RECT 449.200 129.600 450.000 129.700 ;
        RECT 481.200 129.600 482.000 129.700 ;
        RECT 497.200 130.300 498.000 130.400 ;
        RECT 513.200 130.300 514.000 130.400 ;
        RECT 519.600 130.300 520.400 130.400 ;
        RECT 497.200 129.700 520.400 130.300 ;
        RECT 497.200 129.600 498.000 129.700 ;
        RECT 513.200 129.600 514.000 129.700 ;
        RECT 519.600 129.600 520.400 129.700 ;
        RECT 22.000 128.300 22.800 128.400 ;
        RECT 25.200 128.300 26.000 128.400 ;
        RECT 31.600 128.300 32.400 128.400 ;
        RECT 22.000 127.700 32.400 128.300 ;
        RECT 22.000 127.600 22.800 127.700 ;
        RECT 25.200 127.600 26.000 127.700 ;
        RECT 31.600 127.600 32.400 127.700 ;
        RECT 33.200 128.300 34.000 128.400 ;
        RECT 41.200 128.300 42.000 128.400 ;
        RECT 33.200 127.700 42.000 128.300 ;
        RECT 33.200 127.600 34.000 127.700 ;
        RECT 41.200 127.600 42.000 127.700 ;
        RECT 159.600 128.300 160.400 128.400 ;
        RECT 164.400 128.300 165.200 128.400 ;
        RECT 159.600 127.700 165.200 128.300 ;
        RECT 159.600 127.600 160.400 127.700 ;
        RECT 164.400 127.600 165.200 127.700 ;
        RECT 185.200 128.300 186.000 128.400 ;
        RECT 190.000 128.300 190.800 128.400 ;
        RECT 185.200 127.700 190.800 128.300 ;
        RECT 185.200 127.600 186.000 127.700 ;
        RECT 190.000 127.600 190.800 127.700 ;
        RECT 231.600 128.300 232.400 128.400 ;
        RECT 274.800 128.300 275.600 128.400 ;
        RECT 231.600 127.700 275.600 128.300 ;
        RECT 231.600 127.600 232.400 127.700 ;
        RECT 274.800 127.600 275.600 127.700 ;
        RECT 388.400 128.300 389.200 128.400 ;
        RECT 447.600 128.300 448.400 128.400 ;
        RECT 388.400 127.700 448.400 128.300 ;
        RECT 388.400 127.600 389.200 127.700 ;
        RECT 447.600 127.600 448.400 127.700 ;
        RECT 454.000 128.300 454.800 128.400 ;
        RECT 470.000 128.300 470.800 128.400 ;
        RECT 454.000 127.700 470.800 128.300 ;
        RECT 454.000 127.600 454.800 127.700 ;
        RECT 470.000 127.600 470.800 127.700 ;
        RECT 22.000 126.300 22.800 126.400 ;
        RECT 26.800 126.300 27.600 126.400 ;
        RECT 295.600 126.300 296.400 126.400 ;
        RECT 22.000 125.700 27.600 126.300 ;
        RECT 22.000 125.600 22.800 125.700 ;
        RECT 26.800 125.600 27.600 125.700 ;
        RECT 116.500 125.700 296.400 126.300 ;
        RECT 116.500 124.400 117.100 125.700 ;
        RECT 295.600 125.600 296.400 125.700 ;
        RECT 425.200 126.300 426.000 126.400 ;
        RECT 454.000 126.300 454.800 126.400 ;
        RECT 425.200 125.700 454.800 126.300 ;
        RECT 425.200 125.600 426.000 125.700 ;
        RECT 454.000 125.600 454.800 125.700 ;
        RECT 505.200 126.300 506.000 126.400 ;
        RECT 506.800 126.300 507.600 126.400 ;
        RECT 505.200 125.700 507.600 126.300 ;
        RECT 505.200 125.600 506.000 125.700 ;
        RECT 506.800 125.600 507.600 125.700 ;
        RECT 116.400 123.600 117.200 124.400 ;
        RECT 402.800 124.300 403.600 124.400 ;
        RECT 462.000 124.300 462.800 124.400 ;
        RECT 402.800 123.700 462.800 124.300 ;
        RECT 402.800 123.600 403.600 123.700 ;
        RECT 462.000 123.600 462.800 123.700 ;
        RECT 4.400 122.300 5.200 122.400 ;
        RECT 20.400 122.300 21.200 122.400 ;
        RECT 4.400 121.700 21.200 122.300 ;
        RECT 4.400 121.600 5.200 121.700 ;
        RECT 20.400 121.600 21.200 121.700 ;
        RECT 30.000 121.600 30.800 122.400 ;
        RECT 86.000 122.300 86.800 122.400 ;
        RECT 94.000 122.300 94.800 122.400 ;
        RECT 119.600 122.300 120.400 122.400 ;
        RECT 86.000 121.700 120.400 122.300 ;
        RECT 86.000 121.600 86.800 121.700 ;
        RECT 94.000 121.600 94.800 121.700 ;
        RECT 119.600 121.600 120.400 121.700 ;
        RECT 164.400 122.300 165.200 122.400 ;
        RECT 196.400 122.300 197.200 122.400 ;
        RECT 199.600 122.300 200.400 122.400 ;
        RECT 164.400 121.700 200.400 122.300 ;
        RECT 164.400 121.600 165.200 121.700 ;
        RECT 196.400 121.600 197.200 121.700 ;
        RECT 199.600 121.600 200.400 121.700 ;
        RECT 378.800 122.300 379.600 122.400 ;
        RECT 382.000 122.300 382.800 122.400 ;
        RECT 378.800 121.700 382.800 122.300 ;
        RECT 378.800 121.600 379.600 121.700 ;
        RECT 382.000 121.600 382.800 121.700 ;
        RECT 394.800 122.300 395.600 122.400 ;
        RECT 407.600 122.300 408.400 122.400 ;
        RECT 394.800 121.700 408.400 122.300 ;
        RECT 394.800 121.600 395.600 121.700 ;
        RECT 407.600 121.600 408.400 121.700 ;
        RECT 46.000 120.300 46.800 120.400 ;
        RECT 57.200 120.300 58.000 120.400 ;
        RECT 46.000 119.700 58.000 120.300 ;
        RECT 46.000 119.600 46.800 119.700 ;
        RECT 57.200 119.600 58.000 119.700 ;
        RECT 60.400 120.300 61.200 120.400 ;
        RECT 66.800 120.300 67.600 120.400 ;
        RECT 60.400 119.700 67.600 120.300 ;
        RECT 60.400 119.600 61.200 119.700 ;
        RECT 66.800 119.600 67.600 119.700 ;
        RECT 214.000 120.300 214.800 120.400 ;
        RECT 266.800 120.300 267.600 120.400 ;
        RECT 214.000 119.700 267.600 120.300 ;
        RECT 214.000 119.600 214.800 119.700 ;
        RECT 266.800 119.600 267.600 119.700 ;
        RECT 390.000 120.300 390.800 120.400 ;
        RECT 420.400 120.300 421.200 120.400 ;
        RECT 390.000 119.700 421.200 120.300 ;
        RECT 390.000 119.600 390.800 119.700 ;
        RECT 420.400 119.600 421.200 119.700 ;
        RECT 431.600 120.300 432.400 120.400 ;
        RECT 455.600 120.300 456.400 120.400 ;
        RECT 431.600 119.700 456.400 120.300 ;
        RECT 431.600 119.600 432.400 119.700 ;
        RECT 455.600 119.600 456.400 119.700 ;
        RECT 514.800 120.300 515.600 120.400 ;
        RECT 542.000 120.300 542.800 120.400 ;
        RECT 514.800 119.700 542.800 120.300 ;
        RECT 514.800 119.600 515.600 119.700 ;
        RECT 542.000 119.600 542.800 119.700 ;
        RECT 100.400 118.300 101.200 118.400 ;
        RECT 102.000 118.300 102.800 118.400 ;
        RECT 100.400 117.700 102.800 118.300 ;
        RECT 100.400 117.600 101.200 117.700 ;
        RECT 102.000 117.600 102.800 117.700 ;
        RECT 222.000 118.300 222.800 118.400 ;
        RECT 250.800 118.300 251.600 118.400 ;
        RECT 222.000 117.700 251.600 118.300 ;
        RECT 222.000 117.600 222.800 117.700 ;
        RECT 250.800 117.600 251.600 117.700 ;
        RECT 377.200 118.300 378.000 118.400 ;
        RECT 442.800 118.300 443.600 118.400 ;
        RECT 377.200 117.700 443.600 118.300 ;
        RECT 377.200 117.600 378.000 117.700 ;
        RECT 442.800 117.600 443.600 117.700 ;
        RECT 15.600 116.300 16.400 116.400 ;
        RECT 20.400 116.300 21.200 116.400 ;
        RECT 68.400 116.300 69.200 116.400 ;
        RECT 15.600 115.700 69.200 116.300 ;
        RECT 15.600 115.600 16.400 115.700 ;
        RECT 20.400 115.600 21.200 115.700 ;
        RECT 68.400 115.600 69.200 115.700 ;
        RECT 159.600 116.300 160.400 116.400 ;
        RECT 180.400 116.300 181.200 116.400 ;
        RECT 214.000 116.300 214.800 116.400 ;
        RECT 159.600 115.700 214.800 116.300 ;
        RECT 159.600 115.600 160.400 115.700 ;
        RECT 180.400 115.600 181.200 115.700 ;
        RECT 214.000 115.600 214.800 115.700 ;
        RECT 364.400 116.300 365.200 116.400 ;
        RECT 393.200 116.300 394.000 116.400 ;
        RECT 364.400 115.700 394.000 116.300 ;
        RECT 364.400 115.600 365.200 115.700 ;
        RECT 393.200 115.600 394.000 115.700 ;
        RECT 415.600 116.300 416.400 116.400 ;
        RECT 492.400 116.300 493.200 116.400 ;
        RECT 415.600 115.700 493.200 116.300 ;
        RECT 415.600 115.600 416.400 115.700 ;
        RECT 492.400 115.600 493.200 115.700 ;
        RECT 14.000 114.300 14.800 114.400 ;
        RECT 18.800 114.300 19.600 114.400 ;
        RECT 28.400 114.300 29.200 114.400 ;
        RECT 14.000 113.700 29.200 114.300 ;
        RECT 14.000 113.600 14.800 113.700 ;
        RECT 18.800 113.600 19.600 113.700 ;
        RECT 28.400 113.600 29.200 113.700 ;
        RECT 164.400 114.300 165.200 114.400 ;
        RECT 178.800 114.300 179.600 114.400 ;
        RECT 196.400 114.300 197.200 114.400 ;
        RECT 164.400 113.700 197.200 114.300 ;
        RECT 164.400 113.600 165.200 113.700 ;
        RECT 178.800 113.600 179.600 113.700 ;
        RECT 196.400 113.600 197.200 113.700 ;
        RECT 246.000 114.300 246.800 114.400 ;
        RECT 252.400 114.300 253.200 114.400 ;
        RECT 246.000 113.700 253.200 114.300 ;
        RECT 246.000 113.600 246.800 113.700 ;
        RECT 252.400 113.600 253.200 113.700 ;
        RECT 372.400 114.300 373.200 114.400 ;
        RECT 460.400 114.300 461.200 114.400 ;
        RECT 372.400 113.700 461.200 114.300 ;
        RECT 372.400 113.600 373.200 113.700 ;
        RECT 460.400 113.600 461.200 113.700 ;
        RECT 484.400 114.300 485.200 114.400 ;
        RECT 487.600 114.300 488.400 114.400 ;
        RECT 500.400 114.300 501.200 114.400 ;
        RECT 484.400 113.700 501.200 114.300 ;
        RECT 484.400 113.600 485.200 113.700 ;
        RECT 487.600 113.600 488.400 113.700 ;
        RECT 500.400 113.600 501.200 113.700 ;
        RECT 505.200 114.300 506.000 114.400 ;
        RECT 513.200 114.300 514.000 114.400 ;
        RECT 505.200 113.700 514.000 114.300 ;
        RECT 505.200 113.600 506.000 113.700 ;
        RECT 513.200 113.600 514.000 113.700 ;
        RECT 4.400 111.600 5.200 112.400 ;
        RECT 6.000 112.300 6.800 112.400 ;
        RECT 10.800 112.300 11.600 112.400 ;
        RECT 6.000 111.700 11.600 112.300 ;
        RECT 6.000 111.600 6.800 111.700 ;
        RECT 10.800 111.600 11.600 111.700 ;
        RECT 17.200 112.300 18.000 112.400 ;
        RECT 25.200 112.300 26.000 112.400 ;
        RECT 17.200 111.700 26.000 112.300 ;
        RECT 17.200 111.600 18.000 111.700 ;
        RECT 25.200 111.600 26.000 111.700 ;
        RECT 26.800 112.300 27.600 112.400 ;
        RECT 31.600 112.300 32.400 112.400 ;
        RECT 26.800 111.700 32.400 112.300 ;
        RECT 26.800 111.600 27.600 111.700 ;
        RECT 31.600 111.600 32.400 111.700 ;
        RECT 82.800 112.300 83.600 112.400 ;
        RECT 90.800 112.300 91.600 112.400 ;
        RECT 130.800 112.300 131.600 112.400 ;
        RECT 82.800 111.700 131.600 112.300 ;
        RECT 82.800 111.600 83.600 111.700 ;
        RECT 90.800 111.600 91.600 111.700 ;
        RECT 130.800 111.600 131.600 111.700 ;
        RECT 134.000 112.300 134.800 112.400 ;
        RECT 167.600 112.300 168.400 112.400 ;
        RECT 134.000 111.700 168.400 112.300 ;
        RECT 134.000 111.600 134.800 111.700 ;
        RECT 167.600 111.600 168.400 111.700 ;
        RECT 212.400 112.300 213.200 112.400 ;
        RECT 239.600 112.300 240.400 112.400 ;
        RECT 212.400 111.700 240.400 112.300 ;
        RECT 212.400 111.600 213.200 111.700 ;
        RECT 239.600 111.600 240.400 111.700 ;
        RECT 247.600 111.600 248.400 112.400 ;
        RECT 313.200 112.300 314.000 112.400 ;
        RECT 318.000 112.300 318.800 112.400 ;
        RECT 385.200 112.300 386.000 112.400 ;
        RECT 313.200 111.700 318.800 112.300 ;
        RECT 313.200 111.600 314.000 111.700 ;
        RECT 318.000 111.600 318.800 111.700 ;
        RECT 321.300 111.700 386.000 112.300 ;
        RECT 321.300 110.400 321.900 111.700 ;
        RECT 385.200 111.600 386.000 111.700 ;
        RECT 404.400 112.300 405.200 112.400 ;
        RECT 414.000 112.300 414.800 112.400 ;
        RECT 404.400 111.700 414.800 112.300 ;
        RECT 404.400 111.600 405.200 111.700 ;
        RECT 414.000 111.600 414.800 111.700 ;
        RECT 420.400 112.300 421.200 112.400 ;
        RECT 439.600 112.300 440.400 112.400 ;
        RECT 420.400 111.700 440.400 112.300 ;
        RECT 420.400 111.600 421.200 111.700 ;
        RECT 439.600 111.600 440.400 111.700 ;
        RECT 455.600 112.300 456.400 112.400 ;
        RECT 471.600 112.300 472.400 112.400 ;
        RECT 455.600 111.700 472.400 112.300 ;
        RECT 455.600 111.600 456.400 111.700 ;
        RECT 471.600 111.600 472.400 111.700 ;
        RECT 473.200 112.300 474.000 112.400 ;
        RECT 495.600 112.300 496.400 112.400 ;
        RECT 473.200 111.700 496.400 112.300 ;
        RECT 473.200 111.600 474.000 111.700 ;
        RECT 495.600 111.600 496.400 111.700 ;
        RECT 497.200 112.300 498.000 112.400 ;
        RECT 503.600 112.300 504.400 112.400 ;
        RECT 505.200 112.300 506.000 112.400 ;
        RECT 497.200 111.700 506.000 112.300 ;
        RECT 497.200 111.600 498.000 111.700 ;
        RECT 503.600 111.600 504.400 111.700 ;
        RECT 505.200 111.600 506.000 111.700 ;
        RECT 14.000 110.300 14.800 110.400 ;
        RECT 22.000 110.300 22.800 110.400 ;
        RECT 14.000 109.700 22.800 110.300 ;
        RECT 14.000 109.600 14.800 109.700 ;
        RECT 22.000 109.600 22.800 109.700 ;
        RECT 70.000 110.300 70.800 110.400 ;
        RECT 87.600 110.300 88.400 110.400 ;
        RECT 70.000 109.700 88.400 110.300 ;
        RECT 70.000 109.600 70.800 109.700 ;
        RECT 87.600 109.600 88.400 109.700 ;
        RECT 116.400 110.300 117.200 110.400 ;
        RECT 127.600 110.300 128.400 110.400 ;
        RECT 116.400 109.700 128.400 110.300 ;
        RECT 116.400 109.600 117.200 109.700 ;
        RECT 127.600 109.600 128.400 109.700 ;
        RECT 148.400 110.300 149.200 110.400 ;
        RECT 154.800 110.300 155.600 110.400 ;
        RECT 148.400 109.700 155.600 110.300 ;
        RECT 148.400 109.600 149.200 109.700 ;
        RECT 154.800 109.600 155.600 109.700 ;
        RECT 167.600 110.300 168.400 110.400 ;
        RECT 170.800 110.300 171.600 110.400 ;
        RECT 167.600 109.700 171.600 110.300 ;
        RECT 167.600 109.600 168.400 109.700 ;
        RECT 170.800 109.600 171.600 109.700 ;
        RECT 220.400 110.300 221.200 110.400 ;
        RECT 225.200 110.300 226.000 110.400 ;
        RECT 220.400 109.700 226.000 110.300 ;
        RECT 220.400 109.600 221.200 109.700 ;
        RECT 225.200 109.600 226.000 109.700 ;
        RECT 236.400 110.300 237.200 110.400 ;
        RECT 255.600 110.300 256.400 110.400 ;
        RECT 258.800 110.300 259.600 110.400 ;
        RECT 236.400 109.700 259.600 110.300 ;
        RECT 236.400 109.600 237.200 109.700 ;
        RECT 255.600 109.600 256.400 109.700 ;
        RECT 258.800 109.600 259.600 109.700 ;
        RECT 274.800 110.300 275.600 110.400 ;
        RECT 321.200 110.300 322.000 110.400 ;
        RECT 274.800 109.700 322.000 110.300 ;
        RECT 274.800 109.600 275.600 109.700 ;
        RECT 321.200 109.600 322.000 109.700 ;
        RECT 369.200 110.300 370.000 110.400 ;
        RECT 378.800 110.300 379.600 110.400 ;
        RECT 412.400 110.300 413.200 110.400 ;
        RECT 369.200 109.700 413.200 110.300 ;
        RECT 369.200 109.600 370.000 109.700 ;
        RECT 378.800 109.600 379.600 109.700 ;
        RECT 412.400 109.600 413.200 109.700 ;
        RECT 417.200 110.300 418.000 110.400 ;
        RECT 431.600 110.300 432.400 110.400 ;
        RECT 417.200 109.700 432.400 110.300 ;
        RECT 417.200 109.600 418.000 109.700 ;
        RECT 431.600 109.600 432.400 109.700 ;
        RECT 436.400 110.300 437.200 110.400 ;
        RECT 447.600 110.300 448.400 110.400 ;
        RECT 436.400 109.700 448.400 110.300 ;
        RECT 436.400 109.600 437.200 109.700 ;
        RECT 447.600 109.600 448.400 109.700 ;
        RECT 457.200 110.300 458.000 110.400 ;
        RECT 462.000 110.300 462.800 110.400 ;
        RECT 457.200 109.700 462.800 110.300 ;
        RECT 457.200 109.600 458.000 109.700 ;
        RECT 462.000 109.600 462.800 109.700 ;
        RECT 463.600 110.300 464.400 110.400 ;
        RECT 466.800 110.300 467.600 110.400 ;
        RECT 463.600 109.700 467.600 110.300 ;
        RECT 463.600 109.600 464.400 109.700 ;
        RECT 466.800 109.600 467.600 109.700 ;
        RECT 476.400 110.300 477.200 110.400 ;
        RECT 478.000 110.300 478.800 110.400 ;
        RECT 479.600 110.300 480.400 110.400 ;
        RECT 476.400 109.700 480.400 110.300 ;
        RECT 476.400 109.600 477.200 109.700 ;
        RECT 478.000 109.600 478.800 109.700 ;
        RECT 479.600 109.600 480.400 109.700 ;
        RECT 482.800 110.300 483.600 110.400 ;
        RECT 490.800 110.300 491.600 110.400 ;
        RECT 482.800 109.700 491.600 110.300 ;
        RECT 482.800 109.600 483.600 109.700 ;
        RECT 490.800 109.600 491.600 109.700 ;
        RECT 4.400 108.300 5.200 108.400 ;
        RECT 7.600 108.300 8.400 108.400 ;
        RECT 4.400 107.700 8.400 108.300 ;
        RECT 4.400 107.600 5.200 107.700 ;
        RECT 7.600 107.600 8.400 107.700 ;
        RECT 41.200 108.300 42.000 108.400 ;
        RECT 52.400 108.300 53.200 108.400 ;
        RECT 58.800 108.300 59.600 108.400 ;
        RECT 41.200 107.700 59.600 108.300 ;
        RECT 41.200 107.600 42.000 107.700 ;
        RECT 52.400 107.600 53.200 107.700 ;
        RECT 58.800 107.600 59.600 107.700 ;
        RECT 79.600 108.300 80.400 108.400 ;
        RECT 84.400 108.300 85.200 108.400 ;
        RECT 79.600 107.700 85.200 108.300 ;
        RECT 79.600 107.600 80.400 107.700 ;
        RECT 84.400 107.600 85.200 107.700 ;
        RECT 145.200 108.300 146.000 108.400 ;
        RECT 148.400 108.300 149.200 108.400 ;
        RECT 154.800 108.300 155.600 108.400 ;
        RECT 145.200 107.700 155.600 108.300 ;
        RECT 145.200 107.600 146.000 107.700 ;
        RECT 148.400 107.600 149.200 107.700 ;
        RECT 154.800 107.600 155.600 107.700 ;
        RECT 174.000 108.300 174.800 108.400 ;
        RECT 183.600 108.300 184.400 108.400 ;
        RECT 174.000 107.700 184.400 108.300 ;
        RECT 174.000 107.600 174.800 107.700 ;
        RECT 183.600 107.600 184.400 107.700 ;
        RECT 193.200 108.300 194.000 108.400 ;
        RECT 215.600 108.300 216.400 108.400 ;
        RECT 193.200 107.700 216.400 108.300 ;
        RECT 193.200 107.600 194.000 107.700 ;
        RECT 215.600 107.600 216.400 107.700 ;
        RECT 246.000 108.300 246.800 108.400 ;
        RECT 249.200 108.300 250.000 108.400 ;
        RECT 250.800 108.300 251.600 108.400 ;
        RECT 246.000 107.700 251.600 108.300 ;
        RECT 246.000 107.600 246.800 107.700 ;
        RECT 249.200 107.600 250.000 107.700 ;
        RECT 250.800 107.600 251.600 107.700 ;
        RECT 294.000 108.300 294.800 108.400 ;
        RECT 316.400 108.300 317.200 108.400 ;
        RECT 294.000 107.700 317.200 108.300 ;
        RECT 294.000 107.600 294.800 107.700 ;
        RECT 316.400 107.600 317.200 107.700 ;
        RECT 351.600 108.300 352.400 108.400 ;
        RECT 377.200 108.300 378.000 108.400 ;
        RECT 351.600 107.700 378.000 108.300 ;
        RECT 351.600 107.600 352.400 107.700 ;
        RECT 377.200 107.600 378.000 107.700 ;
        RECT 399.600 108.300 400.400 108.400 ;
        RECT 406.000 108.300 406.800 108.400 ;
        RECT 399.600 107.700 406.800 108.300 ;
        RECT 399.600 107.600 400.400 107.700 ;
        RECT 406.000 107.600 406.800 107.700 ;
        RECT 423.600 108.300 424.400 108.400 ;
        RECT 433.200 108.300 434.000 108.400 ;
        RECT 423.600 107.700 434.000 108.300 ;
        RECT 423.600 107.600 424.400 107.700 ;
        RECT 433.200 107.600 434.000 107.700 ;
        RECT 446.000 108.300 446.800 108.400 ;
        RECT 449.200 108.300 450.000 108.400 ;
        RECT 446.000 107.700 450.000 108.300 ;
        RECT 446.000 107.600 446.800 107.700 ;
        RECT 449.200 107.600 450.000 107.700 ;
        RECT 455.600 107.600 456.400 108.400 ;
        RECT 458.800 108.300 459.600 108.400 ;
        RECT 473.200 108.300 474.000 108.400 ;
        RECT 458.800 107.700 474.000 108.300 ;
        RECT 458.800 107.600 459.600 107.700 ;
        RECT 473.200 107.600 474.000 107.700 ;
        RECT 482.800 108.300 483.600 108.400 ;
        RECT 486.000 108.300 486.800 108.400 ;
        RECT 492.400 108.300 493.200 108.400 ;
        RECT 482.800 107.700 493.200 108.300 ;
        RECT 482.800 107.600 483.600 107.700 ;
        RECT 486.000 107.600 486.800 107.700 ;
        RECT 492.400 107.600 493.200 107.700 ;
        RECT 498.800 108.300 499.600 108.400 ;
        RECT 514.800 108.300 515.600 108.400 ;
        RECT 498.800 107.700 515.600 108.300 ;
        RECT 498.800 107.600 499.600 107.700 ;
        RECT 514.800 107.600 515.600 107.700 ;
        RECT 33.200 106.300 34.000 106.400 ;
        RECT 63.600 106.300 64.400 106.400 ;
        RECT 33.200 105.700 64.400 106.300 ;
        RECT 33.200 105.600 34.000 105.700 ;
        RECT 63.600 105.600 64.400 105.700 ;
        RECT 100.400 106.300 101.200 106.400 ;
        RECT 114.800 106.300 115.600 106.400 ;
        RECT 100.400 105.700 115.600 106.300 ;
        RECT 100.400 105.600 101.200 105.700 ;
        RECT 114.800 105.600 115.600 105.700 ;
        RECT 140.400 106.300 141.200 106.400 ;
        RECT 146.800 106.300 147.600 106.400 ;
        RECT 148.400 106.300 149.200 106.400 ;
        RECT 140.400 105.700 149.200 106.300 ;
        RECT 140.400 105.600 141.200 105.700 ;
        RECT 146.800 105.600 147.600 105.700 ;
        RECT 148.400 105.600 149.200 105.700 ;
        RECT 174.000 106.300 174.800 106.400 ;
        RECT 177.200 106.300 178.000 106.400 ;
        RECT 207.600 106.300 208.400 106.400 ;
        RECT 174.000 105.700 208.400 106.300 ;
        RECT 174.000 105.600 174.800 105.700 ;
        RECT 177.200 105.600 178.000 105.700 ;
        RECT 207.600 105.600 208.400 105.700 ;
        RECT 212.400 106.300 213.200 106.400 ;
        RECT 225.200 106.300 226.000 106.400 ;
        RECT 212.400 105.700 226.000 106.300 ;
        RECT 212.400 105.600 213.200 105.700 ;
        RECT 225.200 105.600 226.000 105.700 ;
        RECT 233.200 106.300 234.000 106.400 ;
        RECT 236.400 106.300 237.200 106.400 ;
        RECT 233.200 105.700 237.200 106.300 ;
        RECT 233.200 105.600 234.000 105.700 ;
        RECT 236.400 105.600 237.200 105.700 ;
        RECT 239.600 106.300 240.400 106.400 ;
        RECT 244.400 106.300 245.200 106.400 ;
        RECT 257.200 106.300 258.000 106.400 ;
        RECT 239.600 105.700 258.000 106.300 ;
        RECT 239.600 105.600 240.400 105.700 ;
        RECT 244.400 105.600 245.200 105.700 ;
        RECT 257.200 105.600 258.000 105.700 ;
        RECT 290.800 106.300 291.600 106.400 ;
        RECT 311.600 106.300 312.400 106.400 ;
        RECT 324.400 106.300 325.200 106.400 ;
        RECT 338.800 106.300 339.600 106.400 ;
        RECT 354.800 106.300 355.600 106.400 ;
        RECT 290.800 105.700 355.600 106.300 ;
        RECT 290.800 105.600 291.600 105.700 ;
        RECT 311.600 105.600 312.400 105.700 ;
        RECT 324.400 105.600 325.200 105.700 ;
        RECT 338.800 105.600 339.600 105.700 ;
        RECT 354.800 105.600 355.600 105.700 ;
        RECT 362.800 106.300 363.600 106.400 ;
        RECT 391.600 106.300 392.400 106.400 ;
        RECT 362.800 105.700 392.400 106.300 ;
        RECT 362.800 105.600 363.600 105.700 ;
        RECT 391.600 105.600 392.400 105.700 ;
        RECT 396.400 106.300 397.200 106.400 ;
        RECT 404.400 106.300 405.200 106.400 ;
        RECT 396.400 105.700 405.200 106.300 ;
        RECT 396.400 105.600 397.200 105.700 ;
        RECT 404.400 105.600 405.200 105.700 ;
        RECT 471.600 106.300 472.400 106.400 ;
        RECT 481.200 106.300 482.000 106.400 ;
        RECT 489.200 106.300 490.000 106.400 ;
        RECT 471.600 105.700 490.000 106.300 ;
        RECT 471.600 105.600 472.400 105.700 ;
        RECT 481.200 105.600 482.000 105.700 ;
        RECT 489.200 105.600 490.000 105.700 ;
        RECT 490.800 106.300 491.600 106.400 ;
        RECT 500.400 106.300 501.200 106.400 ;
        RECT 490.800 105.700 501.200 106.300 ;
        RECT 490.800 105.600 491.600 105.700 ;
        RECT 500.400 105.600 501.200 105.700 ;
        RECT 511.600 106.300 512.400 106.400 ;
        RECT 537.200 106.300 538.000 106.400 ;
        RECT 511.600 105.700 538.000 106.300 ;
        RECT 511.600 105.600 512.400 105.700 ;
        RECT 537.200 105.600 538.000 105.700 ;
        RECT 81.200 104.300 82.000 104.400 ;
        RECT 97.200 104.300 98.000 104.400 ;
        RECT 81.200 103.700 98.000 104.300 ;
        RECT 81.200 103.600 82.000 103.700 ;
        RECT 97.200 103.600 98.000 103.700 ;
        RECT 140.400 104.300 141.200 104.400 ;
        RECT 161.200 104.300 162.000 104.400 ;
        RECT 175.600 104.300 176.400 104.400 ;
        RECT 140.400 103.700 176.400 104.300 ;
        RECT 140.400 103.600 141.200 103.700 ;
        RECT 161.200 103.600 162.000 103.700 ;
        RECT 175.600 103.600 176.400 103.700 ;
        RECT 225.200 104.300 226.000 104.400 ;
        RECT 254.000 104.300 254.800 104.400 ;
        RECT 303.600 104.300 304.400 104.400 ;
        RECT 225.200 103.700 304.400 104.300 ;
        RECT 225.200 103.600 226.000 103.700 ;
        RECT 254.000 103.600 254.800 103.700 ;
        RECT 303.600 103.600 304.400 103.700 ;
        RECT 313.200 104.300 314.000 104.400 ;
        RECT 372.400 104.300 373.200 104.400 ;
        RECT 313.200 103.700 373.200 104.300 ;
        RECT 313.200 103.600 314.000 103.700 ;
        RECT 372.400 103.600 373.200 103.700 ;
        RECT 385.200 104.300 386.000 104.400 ;
        RECT 394.800 104.300 395.600 104.400 ;
        RECT 385.200 103.700 395.600 104.300 ;
        RECT 385.200 103.600 386.000 103.700 ;
        RECT 394.800 103.600 395.600 103.700 ;
        RECT 431.600 104.300 432.400 104.400 ;
        RECT 446.000 104.300 446.800 104.400 ;
        RECT 431.600 103.700 446.800 104.300 ;
        RECT 431.600 103.600 432.400 103.700 ;
        RECT 446.000 103.600 446.800 103.700 ;
        RECT 31.600 102.300 32.400 102.400 ;
        RECT 44.400 102.300 45.200 102.400 ;
        RECT 31.600 101.700 45.200 102.300 ;
        RECT 31.600 101.600 32.400 101.700 ;
        RECT 44.400 101.600 45.200 101.700 ;
        RECT 143.600 102.300 144.400 102.400 ;
        RECT 145.200 102.300 146.000 102.400 ;
        RECT 150.000 102.300 150.800 102.400 ;
        RECT 143.600 101.700 150.800 102.300 ;
        RECT 143.600 101.600 144.400 101.700 ;
        RECT 145.200 101.600 146.000 101.700 ;
        RECT 150.000 101.600 150.800 101.700 ;
        RECT 234.800 102.300 235.600 102.400 ;
        RECT 250.800 102.300 251.600 102.400 ;
        RECT 234.800 101.700 251.600 102.300 ;
        RECT 234.800 101.600 235.600 101.700 ;
        RECT 250.800 101.600 251.600 101.700 ;
        RECT 369.200 102.300 370.000 102.400 ;
        RECT 374.000 102.300 374.800 102.400 ;
        RECT 369.200 101.700 374.800 102.300 ;
        RECT 369.200 101.600 370.000 101.700 ;
        RECT 374.000 101.600 374.800 101.700 ;
        RECT 394.800 102.300 395.600 102.400 ;
        RECT 422.000 102.300 422.800 102.400 ;
        RECT 394.800 101.700 422.800 102.300 ;
        RECT 394.800 101.600 395.600 101.700 ;
        RECT 422.000 101.600 422.800 101.700 ;
        RECT 441.200 102.300 442.000 102.400 ;
        RECT 468.400 102.300 469.200 102.400 ;
        RECT 441.200 101.700 469.200 102.300 ;
        RECT 441.200 101.600 442.000 101.700 ;
        RECT 468.400 101.600 469.200 101.700 ;
        RECT 103.600 100.300 104.400 100.400 ;
        RECT 108.400 100.300 109.200 100.400 ;
        RECT 103.600 99.700 109.200 100.300 ;
        RECT 103.600 99.600 104.400 99.700 ;
        RECT 108.400 99.600 109.200 99.700 ;
        RECT 138.800 100.300 139.600 100.400 ;
        RECT 188.400 100.300 189.200 100.400 ;
        RECT 222.000 100.300 222.800 100.400 ;
        RECT 138.800 99.700 222.800 100.300 ;
        RECT 138.800 99.600 139.600 99.700 ;
        RECT 188.400 99.600 189.200 99.700 ;
        RECT 222.000 99.600 222.800 99.700 ;
        RECT 246.000 100.300 246.800 100.400 ;
        RECT 262.000 100.300 262.800 100.400 ;
        RECT 246.000 99.700 262.800 100.300 ;
        RECT 246.000 99.600 246.800 99.700 ;
        RECT 262.000 99.600 262.800 99.700 ;
        RECT 286.000 100.300 286.800 100.400 ;
        RECT 290.800 100.300 291.600 100.400 ;
        RECT 286.000 99.700 291.600 100.300 ;
        RECT 286.000 99.600 286.800 99.700 ;
        RECT 290.800 99.600 291.600 99.700 ;
        RECT 337.200 100.300 338.000 100.400 ;
        RECT 342.000 100.300 342.800 100.400 ;
        RECT 337.200 99.700 342.800 100.300 ;
        RECT 337.200 99.600 338.000 99.700 ;
        RECT 342.000 99.600 342.800 99.700 ;
        RECT 370.800 100.300 371.600 100.400 ;
        RECT 383.600 100.300 384.400 100.400 ;
        RECT 370.800 99.700 384.400 100.300 ;
        RECT 370.800 99.600 371.600 99.700 ;
        RECT 383.600 99.600 384.400 99.700 ;
        RECT 393.200 100.300 394.000 100.400 ;
        RECT 446.000 100.300 446.800 100.400 ;
        RECT 393.200 99.700 446.800 100.300 ;
        RECT 393.200 99.600 394.000 99.700 ;
        RECT 446.000 99.600 446.800 99.700 ;
        RECT 497.200 99.600 498.000 100.400 ;
        RECT 503.600 100.300 504.400 100.400 ;
        RECT 537.200 100.300 538.000 100.400 ;
        RECT 503.600 99.700 538.000 100.300 ;
        RECT 503.600 99.600 504.400 99.700 ;
        RECT 537.200 99.600 538.000 99.700 ;
        RECT 28.400 98.300 29.200 98.400 ;
        RECT 33.200 98.300 34.000 98.400 ;
        RECT 42.800 98.300 43.600 98.400 ;
        RECT 44.400 98.300 45.200 98.400 ;
        RECT 28.400 97.700 45.200 98.300 ;
        RECT 28.400 97.600 29.200 97.700 ;
        RECT 33.200 97.600 34.000 97.700 ;
        RECT 42.800 97.600 43.600 97.700 ;
        RECT 44.400 97.600 45.200 97.700 ;
        RECT 46.000 98.300 46.800 98.400 ;
        RECT 49.200 98.300 50.000 98.400 ;
        RECT 46.000 97.700 50.000 98.300 ;
        RECT 46.000 97.600 46.800 97.700 ;
        RECT 49.200 97.600 50.000 97.700 ;
        RECT 153.200 98.300 154.000 98.400 ;
        RECT 174.000 98.300 174.800 98.400 ;
        RECT 183.600 98.300 184.400 98.400 ;
        RECT 153.200 97.700 184.400 98.300 ;
        RECT 153.200 97.600 154.000 97.700 ;
        RECT 174.000 97.600 174.800 97.700 ;
        RECT 183.600 97.600 184.400 97.700 ;
        RECT 209.200 98.300 210.000 98.400 ;
        RECT 218.800 98.300 219.600 98.400 ;
        RECT 209.200 97.700 219.600 98.300 ;
        RECT 209.200 97.600 210.000 97.700 ;
        RECT 218.800 97.600 219.600 97.700 ;
        RECT 225.200 98.300 226.000 98.400 ;
        RECT 228.400 98.300 229.200 98.400 ;
        RECT 225.200 97.700 229.200 98.300 ;
        RECT 225.200 97.600 226.000 97.700 ;
        RECT 228.400 97.600 229.200 97.700 ;
        RECT 262.000 98.300 262.800 98.400 ;
        RECT 308.400 98.300 309.200 98.400 ;
        RECT 262.000 97.700 309.200 98.300 ;
        RECT 262.000 97.600 262.800 97.700 ;
        RECT 308.400 97.600 309.200 97.700 ;
        RECT 367.600 98.300 368.400 98.400 ;
        RECT 409.200 98.300 410.000 98.400 ;
        RECT 367.600 97.700 410.000 98.300 ;
        RECT 367.600 97.600 368.400 97.700 ;
        RECT 409.200 97.600 410.000 97.700 ;
        RECT 415.600 98.300 416.400 98.400 ;
        RECT 455.600 98.300 456.400 98.400 ;
        RECT 415.600 97.700 456.400 98.300 ;
        RECT 415.600 97.600 416.400 97.700 ;
        RECT 455.600 97.600 456.400 97.700 ;
        RECT 458.800 98.300 459.600 98.400 ;
        RECT 474.800 98.300 475.600 98.400 ;
        RECT 458.800 97.700 475.600 98.300 ;
        RECT 458.800 97.600 459.600 97.700 ;
        RECT 474.800 97.600 475.600 97.700 ;
        RECT 478.000 98.300 478.800 98.400 ;
        RECT 502.000 98.300 502.800 98.400 ;
        RECT 508.400 98.300 509.200 98.400 ;
        RECT 518.000 98.300 518.800 98.400 ;
        RECT 478.000 97.700 518.800 98.300 ;
        RECT 478.000 97.600 478.800 97.700 ;
        RECT 502.000 97.600 502.800 97.700 ;
        RECT 508.400 97.600 509.200 97.700 ;
        RECT 518.000 97.600 518.800 97.700 ;
        RECT 14.000 96.300 14.800 96.400 ;
        RECT 23.600 96.300 24.400 96.400 ;
        RECT 14.000 95.700 24.400 96.300 ;
        RECT 14.000 95.600 14.800 95.700 ;
        RECT 23.600 95.600 24.400 95.700 ;
        RECT 39.600 96.300 40.400 96.400 ;
        RECT 46.000 96.300 46.800 96.400 ;
        RECT 39.600 95.700 46.800 96.300 ;
        RECT 39.600 95.600 40.400 95.700 ;
        RECT 46.000 95.600 46.800 95.700 ;
        RECT 79.600 96.300 80.400 96.400 ;
        RECT 87.600 96.300 88.400 96.400 ;
        RECT 79.600 95.700 88.400 96.300 ;
        RECT 79.600 95.600 80.400 95.700 ;
        RECT 87.600 95.600 88.400 95.700 ;
        RECT 137.200 96.300 138.000 96.400 ;
        RECT 142.000 96.300 142.800 96.400 ;
        RECT 137.200 95.700 142.800 96.300 ;
        RECT 137.200 95.600 138.000 95.700 ;
        RECT 142.000 95.600 142.800 95.700 ;
        RECT 207.600 96.300 208.400 96.400 ;
        RECT 222.000 96.300 222.800 96.400 ;
        RECT 207.600 95.700 222.800 96.300 ;
        RECT 207.600 95.600 208.400 95.700 ;
        RECT 222.000 95.600 222.800 95.700 ;
        RECT 226.800 96.300 227.600 96.400 ;
        RECT 234.800 96.300 235.600 96.400 ;
        RECT 226.800 95.700 235.600 96.300 ;
        RECT 226.800 95.600 227.600 95.700 ;
        RECT 234.800 95.600 235.600 95.700 ;
        RECT 242.800 96.300 243.600 96.400 ;
        RECT 249.200 96.300 250.000 96.400 ;
        RECT 260.400 96.300 261.200 96.400 ;
        RECT 242.800 95.700 261.200 96.300 ;
        RECT 242.800 95.600 243.600 95.700 ;
        RECT 249.200 95.600 250.000 95.700 ;
        RECT 260.400 95.600 261.200 95.700 ;
        RECT 303.600 96.300 304.400 96.400 ;
        RECT 306.800 96.300 307.600 96.400 ;
        RECT 303.600 95.700 307.600 96.300 ;
        RECT 303.600 95.600 304.400 95.700 ;
        RECT 306.800 95.600 307.600 95.700 ;
        RECT 354.800 96.300 355.600 96.400 ;
        RECT 370.800 96.300 371.600 96.400 ;
        RECT 354.800 95.700 371.600 96.300 ;
        RECT 354.800 95.600 355.600 95.700 ;
        RECT 370.800 95.600 371.600 95.700 ;
        RECT 390.000 96.300 390.800 96.400 ;
        RECT 410.800 96.300 411.600 96.400 ;
        RECT 438.000 96.300 438.800 96.400 ;
        RECT 452.400 96.300 453.200 96.400 ;
        RECT 390.000 95.700 409.900 96.300 ;
        RECT 390.000 95.600 390.800 95.700 ;
        RECT 15.600 94.300 16.400 94.400 ;
        RECT 30.000 94.300 30.800 94.400 ;
        RECT 15.600 93.700 30.800 94.300 ;
        RECT 15.600 93.600 16.400 93.700 ;
        RECT 30.000 93.600 30.800 93.700 ;
        RECT 50.800 94.300 51.600 94.400 ;
        RECT 52.400 94.300 53.200 94.400 ;
        RECT 50.800 93.700 53.200 94.300 ;
        RECT 50.800 93.600 51.600 93.700 ;
        RECT 52.400 93.600 53.200 93.700 ;
        RECT 58.800 94.300 59.600 94.400 ;
        RECT 90.800 94.300 91.600 94.400 ;
        RECT 58.800 93.700 91.600 94.300 ;
        RECT 58.800 93.600 59.600 93.700 ;
        RECT 90.800 93.600 91.600 93.700 ;
        RECT 111.600 94.300 112.400 94.400 ;
        RECT 135.600 94.300 136.400 94.400 ;
        RECT 111.600 93.700 136.400 94.300 ;
        RECT 111.600 93.600 112.400 93.700 ;
        RECT 135.600 93.600 136.400 93.700 ;
        RECT 193.200 93.600 194.000 94.400 ;
        RECT 204.400 94.300 205.200 94.400 ;
        RECT 212.400 94.300 213.200 94.400 ;
        RECT 204.400 93.700 213.200 94.300 ;
        RECT 204.400 93.600 205.200 93.700 ;
        RECT 212.400 93.600 213.200 93.700 ;
        RECT 218.800 94.300 219.600 94.400 ;
        RECT 223.600 94.300 224.400 94.400 ;
        RECT 218.800 93.700 224.400 94.300 ;
        RECT 218.800 93.600 219.600 93.700 ;
        RECT 223.600 93.600 224.400 93.700 ;
        RECT 225.200 94.300 226.000 94.400 ;
        RECT 228.400 94.300 229.200 94.400 ;
        RECT 225.200 93.700 229.200 94.300 ;
        RECT 225.200 93.600 226.000 93.700 ;
        RECT 228.400 93.600 229.200 93.700 ;
        RECT 231.600 94.300 232.400 94.400 ;
        RECT 236.400 94.300 237.200 94.400 ;
        RECT 231.600 93.700 237.200 94.300 ;
        RECT 231.600 93.600 232.400 93.700 ;
        RECT 236.400 93.600 237.200 93.700 ;
        RECT 263.600 94.300 264.400 94.400 ;
        RECT 289.200 94.300 290.000 94.400 ;
        RECT 263.600 93.700 290.000 94.300 ;
        RECT 263.600 93.600 264.400 93.700 ;
        RECT 289.200 93.600 290.000 93.700 ;
        RECT 327.600 94.300 328.400 94.400 ;
        RECT 345.200 94.300 346.000 94.400 ;
        RECT 327.600 93.700 346.000 94.300 ;
        RECT 327.600 93.600 328.400 93.700 ;
        RECT 345.200 93.600 346.000 93.700 ;
        RECT 353.200 94.300 354.000 94.400 ;
        RECT 396.400 94.300 397.200 94.400 ;
        RECT 353.200 93.700 397.200 94.300 ;
        RECT 353.200 93.600 354.000 93.700 ;
        RECT 396.400 93.600 397.200 93.700 ;
        RECT 398.000 94.300 398.800 94.400 ;
        RECT 402.800 94.300 403.600 94.400 ;
        RECT 404.400 94.300 405.200 94.400 ;
        RECT 398.000 93.700 405.200 94.300 ;
        RECT 398.000 93.600 398.800 93.700 ;
        RECT 402.800 93.600 403.600 93.700 ;
        RECT 404.400 93.600 405.200 93.700 ;
        RECT 407.600 93.600 408.400 94.400 ;
        RECT 409.300 94.300 409.900 95.700 ;
        RECT 410.800 95.700 453.200 96.300 ;
        RECT 410.800 95.600 411.600 95.700 ;
        RECT 438.000 95.600 438.800 95.700 ;
        RECT 452.400 95.600 453.200 95.700 ;
        RECT 465.200 96.300 466.000 96.400 ;
        RECT 468.400 96.300 469.200 96.400 ;
        RECT 465.200 95.700 469.200 96.300 ;
        RECT 465.200 95.600 466.000 95.700 ;
        RECT 468.400 95.600 469.200 95.700 ;
        RECT 498.800 96.300 499.600 96.400 ;
        RECT 534.000 96.300 534.800 96.400 ;
        RECT 498.800 95.700 534.800 96.300 ;
        RECT 498.800 95.600 499.600 95.700 ;
        RECT 534.000 95.600 534.800 95.700 ;
        RECT 438.000 94.300 438.800 94.400 ;
        RECT 409.300 93.700 438.800 94.300 ;
        RECT 438.000 93.600 438.800 93.700 ;
        RECT 441.200 94.300 442.000 94.400 ;
        RECT 458.800 94.300 459.600 94.400 ;
        RECT 441.200 93.700 459.600 94.300 ;
        RECT 441.200 93.600 442.000 93.700 ;
        RECT 458.800 93.600 459.600 93.700 ;
        RECT 465.200 94.300 466.000 94.400 ;
        RECT 479.600 94.300 480.400 94.400 ;
        RECT 465.200 93.700 480.400 94.300 ;
        RECT 465.200 93.600 466.000 93.700 ;
        RECT 479.600 93.600 480.400 93.700 ;
        RECT 20.400 92.300 21.200 92.400 ;
        RECT 23.600 92.300 24.400 92.400 ;
        RECT 20.400 91.700 24.400 92.300 ;
        RECT 20.400 91.600 21.200 91.700 ;
        RECT 23.600 91.600 24.400 91.700 ;
        RECT 26.800 92.300 27.600 92.400 ;
        RECT 39.600 92.300 40.400 92.400 ;
        RECT 26.800 91.700 40.400 92.300 ;
        RECT 26.800 91.600 27.600 91.700 ;
        RECT 39.600 91.600 40.400 91.700 ;
        RECT 82.800 92.300 83.600 92.400 ;
        RECT 87.600 92.300 88.400 92.400 ;
        RECT 90.800 92.300 91.600 92.400 ;
        RECT 95.600 92.300 96.400 92.400 ;
        RECT 82.800 91.700 96.400 92.300 ;
        RECT 82.800 91.600 83.600 91.700 ;
        RECT 87.600 91.600 88.400 91.700 ;
        RECT 90.800 91.600 91.600 91.700 ;
        RECT 95.600 91.600 96.400 91.700 ;
        RECT 97.200 92.300 98.000 92.400 ;
        RECT 100.400 92.300 101.200 92.400 ;
        RECT 97.200 91.700 101.200 92.300 ;
        RECT 97.200 91.600 98.000 91.700 ;
        RECT 100.400 91.600 101.200 91.700 ;
        RECT 150.000 92.300 150.800 92.400 ;
        RECT 153.200 92.300 154.000 92.400 ;
        RECT 241.200 92.300 242.000 92.400 ;
        RECT 247.600 92.300 248.400 92.400 ;
        RECT 257.200 92.300 258.000 92.400 ;
        RECT 150.000 91.700 154.000 92.300 ;
        RECT 150.000 91.600 150.800 91.700 ;
        RECT 153.200 91.600 154.000 91.700 ;
        RECT 212.500 91.700 258.000 92.300 ;
        RECT 212.500 90.400 213.100 91.700 ;
        RECT 241.200 91.600 242.000 91.700 ;
        RECT 247.600 91.600 248.400 91.700 ;
        RECT 257.200 91.600 258.000 91.700 ;
        RECT 314.800 92.300 315.600 92.400 ;
        RECT 343.600 92.300 344.400 92.400 ;
        RECT 348.400 92.300 349.200 92.400 ;
        RECT 314.800 91.700 349.200 92.300 ;
        RECT 314.800 91.600 315.600 91.700 ;
        RECT 343.600 91.600 344.400 91.700 ;
        RECT 348.400 91.600 349.200 91.700 ;
        RECT 390.000 92.300 390.800 92.400 ;
        RECT 415.600 92.300 416.400 92.400 ;
        RECT 390.000 91.700 416.400 92.300 ;
        RECT 390.000 91.600 390.800 91.700 ;
        RECT 415.600 91.600 416.400 91.700 ;
        RECT 463.600 92.300 464.400 92.400 ;
        RECT 487.600 92.300 488.400 92.400 ;
        RECT 463.600 91.700 488.400 92.300 ;
        RECT 463.600 91.600 464.400 91.700 ;
        RECT 487.600 91.600 488.400 91.700 ;
        RECT 511.600 92.300 512.400 92.400 ;
        RECT 526.000 92.300 526.800 92.400 ;
        RECT 511.600 91.700 526.800 92.300 ;
        RECT 511.600 91.600 512.400 91.700 ;
        RECT 526.000 91.600 526.800 91.700 ;
        RECT 1.200 90.300 2.000 90.400 ;
        RECT 15.600 90.300 16.400 90.400 ;
        RECT 17.200 90.300 18.000 90.400 ;
        RECT 22.000 90.300 22.800 90.400 ;
        RECT 1.200 89.700 22.800 90.300 ;
        RECT 1.200 89.600 2.000 89.700 ;
        RECT 15.600 89.600 16.400 89.700 ;
        RECT 17.200 89.600 18.000 89.700 ;
        RECT 22.000 89.600 22.800 89.700 ;
        RECT 23.600 90.300 24.400 90.400 ;
        RECT 41.200 90.300 42.000 90.400 ;
        RECT 23.600 89.700 42.000 90.300 ;
        RECT 23.600 89.600 24.400 89.700 ;
        RECT 41.200 89.600 42.000 89.700 ;
        RECT 153.200 90.300 154.000 90.400 ;
        RECT 161.200 90.300 162.000 90.400 ;
        RECT 153.200 89.700 162.000 90.300 ;
        RECT 153.200 89.600 154.000 89.700 ;
        RECT 161.200 89.600 162.000 89.700 ;
        RECT 199.600 90.300 200.400 90.400 ;
        RECT 212.400 90.300 213.200 90.400 ;
        RECT 199.600 89.700 213.200 90.300 ;
        RECT 199.600 89.600 200.400 89.700 ;
        RECT 212.400 89.600 213.200 89.700 ;
        RECT 222.000 90.300 222.800 90.400 ;
        RECT 226.800 90.300 227.600 90.400 ;
        RECT 222.000 89.700 227.600 90.300 ;
        RECT 222.000 89.600 222.800 89.700 ;
        RECT 226.800 89.600 227.600 89.700 ;
        RECT 386.800 90.300 387.600 90.400 ;
        RECT 390.000 90.300 390.800 90.400 ;
        RECT 393.200 90.300 394.000 90.400 ;
        RECT 386.800 89.700 394.000 90.300 ;
        RECT 386.800 89.600 387.600 89.700 ;
        RECT 390.000 89.600 390.800 89.700 ;
        RECT 393.200 89.600 394.000 89.700 ;
        RECT 396.400 90.300 397.200 90.400 ;
        RECT 404.400 90.300 405.200 90.400 ;
        RECT 396.400 89.700 405.200 90.300 ;
        RECT 396.400 89.600 397.200 89.700 ;
        RECT 404.400 89.600 405.200 89.700 ;
        RECT 407.600 90.300 408.400 90.400 ;
        RECT 412.400 90.300 413.200 90.400 ;
        RECT 449.200 90.300 450.000 90.400 ;
        RECT 455.600 90.300 456.400 90.400 ;
        RECT 468.400 90.300 469.200 90.400 ;
        RECT 407.600 89.700 469.200 90.300 ;
        RECT 407.600 89.600 408.400 89.700 ;
        RECT 412.400 89.600 413.200 89.700 ;
        RECT 449.200 89.600 450.000 89.700 ;
        RECT 455.600 89.600 456.400 89.700 ;
        RECT 468.400 89.600 469.200 89.700 ;
        RECT 473.200 90.300 474.000 90.400 ;
        RECT 478.000 90.300 478.800 90.400 ;
        RECT 473.200 89.700 478.800 90.300 ;
        RECT 473.200 89.600 474.000 89.700 ;
        RECT 478.000 89.600 478.800 89.700 ;
        RECT 4.400 88.300 5.200 88.400 ;
        RECT 12.400 88.300 13.200 88.400 ;
        RECT 18.800 88.300 19.600 88.400 ;
        RECT 4.400 87.700 19.600 88.300 ;
        RECT 4.400 87.600 5.200 87.700 ;
        RECT 12.400 87.600 13.200 87.700 ;
        RECT 18.800 87.600 19.600 87.700 ;
        RECT 20.400 88.300 21.200 88.400 ;
        RECT 25.200 88.300 26.000 88.400 ;
        RECT 20.400 87.700 26.000 88.300 ;
        RECT 20.400 87.600 21.200 87.700 ;
        RECT 25.200 87.600 26.000 87.700 ;
        RECT 30.000 88.300 30.800 88.400 ;
        RECT 38.000 88.300 38.800 88.400 ;
        RECT 30.000 87.700 38.800 88.300 ;
        RECT 30.000 87.600 30.800 87.700 ;
        RECT 38.000 87.600 38.800 87.700 ;
        RECT 154.800 88.300 155.600 88.400 ;
        RECT 161.200 88.300 162.000 88.400 ;
        RECT 154.800 87.700 162.000 88.300 ;
        RECT 154.800 87.600 155.600 87.700 ;
        RECT 161.200 87.600 162.000 87.700 ;
        RECT 204.400 88.300 205.200 88.400 ;
        RECT 238.000 88.300 238.800 88.400 ;
        RECT 204.400 87.700 238.800 88.300 ;
        RECT 204.400 87.600 205.200 87.700 ;
        RECT 238.000 87.600 238.800 87.700 ;
        RECT 385.200 88.300 386.000 88.400 ;
        RECT 439.600 88.300 440.400 88.400 ;
        RECT 385.200 87.700 440.400 88.300 ;
        RECT 385.200 87.600 386.000 87.700 ;
        RECT 439.600 87.600 440.400 87.700 ;
        RECT 185.200 86.300 186.000 86.400 ;
        RECT 263.600 86.300 264.400 86.400 ;
        RECT 185.200 85.700 264.400 86.300 ;
        RECT 185.200 85.600 186.000 85.700 ;
        RECT 263.600 85.600 264.400 85.700 ;
        RECT 402.800 86.300 403.600 86.400 ;
        RECT 417.200 86.300 418.000 86.400 ;
        RECT 430.000 86.300 430.800 86.400 ;
        RECT 402.800 85.700 430.800 86.300 ;
        RECT 402.800 85.600 403.600 85.700 ;
        RECT 417.200 85.600 418.000 85.700 ;
        RECT 430.000 85.600 430.800 85.700 ;
        RECT 436.400 86.300 437.200 86.400 ;
        RECT 442.800 86.300 443.600 86.400 ;
        RECT 436.400 85.700 443.600 86.300 ;
        RECT 436.400 85.600 437.200 85.700 ;
        RECT 442.800 85.600 443.600 85.700 ;
        RECT 326.000 84.300 326.800 84.400 ;
        RECT 342.000 84.300 342.800 84.400 ;
        RECT 326.000 83.700 342.800 84.300 ;
        RECT 326.000 83.600 326.800 83.700 ;
        RECT 342.000 83.600 342.800 83.700 ;
        RECT 378.800 84.300 379.600 84.400 ;
        RECT 418.800 84.300 419.600 84.400 ;
        RECT 378.800 83.700 419.600 84.300 ;
        RECT 378.800 83.600 379.600 83.700 ;
        RECT 418.800 83.600 419.600 83.700 ;
        RECT 433.200 84.300 434.000 84.400 ;
        RECT 441.200 84.300 442.000 84.400 ;
        RECT 433.200 83.700 442.000 84.300 ;
        RECT 433.200 83.600 434.000 83.700 ;
        RECT 441.200 83.600 442.000 83.700 ;
        RECT 442.800 84.300 443.600 84.400 ;
        RECT 444.400 84.300 445.200 84.400 ;
        RECT 442.800 83.700 445.200 84.300 ;
        RECT 442.800 83.600 443.600 83.700 ;
        RECT 444.400 83.600 445.200 83.700 ;
        RECT 15.600 82.300 16.400 82.400 ;
        RECT 30.000 82.300 30.800 82.400 ;
        RECT 15.600 81.700 30.800 82.300 ;
        RECT 15.600 81.600 16.400 81.700 ;
        RECT 30.000 81.600 30.800 81.700 ;
        RECT 62.000 82.300 62.800 82.400 ;
        RECT 65.200 82.300 66.000 82.400 ;
        RECT 62.000 81.700 66.000 82.300 ;
        RECT 62.000 81.600 62.800 81.700 ;
        RECT 65.200 81.600 66.000 81.700 ;
        RECT 353.200 81.600 354.000 82.400 ;
        RECT 436.400 82.300 437.200 82.400 ;
        RECT 446.000 82.300 446.800 82.400 ;
        RECT 436.400 81.700 446.800 82.300 ;
        RECT 436.400 81.600 437.200 81.700 ;
        RECT 446.000 81.600 446.800 81.700 ;
        RECT 542.000 82.300 542.800 82.400 ;
        RECT 545.200 82.300 546.000 82.400 ;
        RECT 542.000 81.700 546.000 82.300 ;
        RECT 542.000 81.600 542.800 81.700 ;
        RECT 545.200 81.600 546.000 81.700 ;
        RECT 134.000 80.300 134.800 80.400 ;
        RECT 145.200 80.300 146.000 80.400 ;
        RECT 134.000 79.700 146.000 80.300 ;
        RECT 134.000 79.600 134.800 79.700 ;
        RECT 145.200 79.600 146.000 79.700 ;
        RECT 185.200 80.300 186.000 80.400 ;
        RECT 193.200 80.300 194.000 80.400 ;
        RECT 185.200 79.700 194.000 80.300 ;
        RECT 185.200 79.600 186.000 79.700 ;
        RECT 193.200 79.600 194.000 79.700 ;
        RECT 228.400 80.300 229.200 80.400 ;
        RECT 231.600 80.300 232.400 80.400 ;
        RECT 228.400 79.700 232.400 80.300 ;
        RECT 228.400 79.600 229.200 79.700 ;
        RECT 231.600 79.600 232.400 79.700 ;
        RECT 286.000 80.300 286.800 80.400 ;
        RECT 290.800 80.300 291.600 80.400 ;
        RECT 286.000 79.700 291.600 80.300 ;
        RECT 286.000 79.600 286.800 79.700 ;
        RECT 290.800 79.600 291.600 79.700 ;
        RECT 308.400 80.300 309.200 80.400 ;
        RECT 378.800 80.300 379.600 80.400 ;
        RECT 308.400 79.700 379.600 80.300 ;
        RECT 308.400 79.600 309.200 79.700 ;
        RECT 378.800 79.600 379.600 79.700 ;
        RECT 466.800 78.300 467.600 78.400 ;
        RECT 484.400 78.300 485.200 78.400 ;
        RECT 466.800 77.700 485.200 78.300 ;
        RECT 466.800 77.600 467.600 77.700 ;
        RECT 484.400 77.600 485.200 77.700 ;
        RECT 305.200 76.300 306.000 76.400 ;
        RECT 326.000 76.300 326.800 76.400 ;
        RECT 305.200 75.700 326.800 76.300 ;
        RECT 305.200 75.600 306.000 75.700 ;
        RECT 326.000 75.600 326.800 75.700 ;
        RECT 334.000 76.300 334.800 76.400 ;
        RECT 372.400 76.300 373.200 76.400 ;
        RECT 334.000 75.700 373.200 76.300 ;
        RECT 334.000 75.600 334.800 75.700 ;
        RECT 372.400 75.600 373.200 75.700 ;
        RECT 497.200 76.300 498.000 76.400 ;
        RECT 498.800 76.300 499.600 76.400 ;
        RECT 497.200 75.700 499.600 76.300 ;
        RECT 497.200 75.600 498.000 75.700 ;
        RECT 498.800 75.600 499.600 75.700 ;
        RECT 503.600 76.300 504.400 76.400 ;
        RECT 506.800 76.300 507.600 76.400 ;
        RECT 514.800 76.300 515.600 76.400 ;
        RECT 503.600 75.700 515.600 76.300 ;
        RECT 503.600 75.600 504.400 75.700 ;
        RECT 506.800 75.600 507.600 75.700 ;
        RECT 514.800 75.600 515.600 75.700 ;
        RECT 7.600 74.300 8.400 74.400 ;
        RECT 52.400 74.300 53.200 74.400 ;
        RECT 84.400 74.300 85.200 74.400 ;
        RECT 7.600 73.700 85.200 74.300 ;
        RECT 7.600 73.600 8.400 73.700 ;
        RECT 52.400 73.600 53.200 73.700 ;
        RECT 84.400 73.600 85.200 73.700 ;
        RECT 228.400 74.300 229.200 74.400 ;
        RECT 247.600 74.300 248.400 74.400 ;
        RECT 313.200 74.300 314.000 74.400 ;
        RECT 228.400 73.700 314.000 74.300 ;
        RECT 228.400 73.600 229.200 73.700 ;
        RECT 247.600 73.600 248.400 73.700 ;
        RECT 313.200 73.600 314.000 73.700 ;
        RECT 358.000 74.300 358.800 74.400 ;
        RECT 375.600 74.300 376.400 74.400 ;
        RECT 358.000 73.700 376.400 74.300 ;
        RECT 358.000 73.600 358.800 73.700 ;
        RECT 375.600 73.600 376.400 73.700 ;
        RECT 377.200 74.300 378.000 74.400 ;
        RECT 391.600 74.300 392.400 74.400 ;
        RECT 377.200 73.700 392.400 74.300 ;
        RECT 377.200 73.600 378.000 73.700 ;
        RECT 391.600 73.600 392.400 73.700 ;
        RECT 447.600 74.300 448.400 74.400 ;
        RECT 450.800 74.300 451.600 74.400 ;
        RECT 447.600 73.700 451.600 74.300 ;
        RECT 447.600 73.600 448.400 73.700 ;
        RECT 450.800 73.600 451.600 73.700 ;
        RECT 471.600 73.600 472.400 74.400 ;
        RECT 484.400 74.300 485.200 74.400 ;
        RECT 510.000 74.300 510.800 74.400 ;
        RECT 484.400 73.700 510.800 74.300 ;
        RECT 484.400 73.600 485.200 73.700 ;
        RECT 510.000 73.600 510.800 73.700 ;
        RECT 36.400 72.300 37.200 72.400 ;
        RECT 39.600 72.300 40.400 72.400 ;
        RECT 36.400 71.700 40.400 72.300 ;
        RECT 36.400 71.600 37.200 71.700 ;
        RECT 39.600 71.600 40.400 71.700 ;
        RECT 58.800 71.600 59.600 72.400 ;
        RECT 162.800 72.300 163.600 72.400 ;
        RECT 167.600 72.300 168.400 72.400 ;
        RECT 177.200 72.300 178.000 72.400 ;
        RECT 162.800 71.700 178.000 72.300 ;
        RECT 162.800 71.600 163.600 71.700 ;
        RECT 167.600 71.600 168.400 71.700 ;
        RECT 177.200 71.600 178.000 71.700 ;
        RECT 252.400 72.300 253.200 72.400 ;
        RECT 257.200 72.300 258.000 72.400 ;
        RECT 330.800 72.300 331.600 72.400 ;
        RECT 385.200 72.300 386.000 72.400 ;
        RECT 252.400 71.700 310.700 72.300 ;
        RECT 252.400 71.600 253.200 71.700 ;
        RECT 257.200 71.600 258.000 71.700 ;
        RECT 310.100 70.400 310.700 71.700 ;
        RECT 330.800 71.700 386.000 72.300 ;
        RECT 330.800 71.600 331.600 71.700 ;
        RECT 385.200 71.600 386.000 71.700 ;
        RECT 391.600 72.300 392.400 72.400 ;
        RECT 396.400 72.300 397.200 72.400 ;
        RECT 391.600 71.700 397.200 72.300 ;
        RECT 391.600 71.600 392.400 71.700 ;
        RECT 396.400 71.600 397.200 71.700 ;
        RECT 425.200 72.300 426.000 72.400 ;
        RECT 470.000 72.300 470.800 72.400 ;
        RECT 425.200 71.700 470.800 72.300 ;
        RECT 425.200 71.600 426.000 71.700 ;
        RECT 470.000 71.600 470.800 71.700 ;
        RECT 490.800 72.300 491.600 72.400 ;
        RECT 503.600 72.300 504.400 72.400 ;
        RECT 505.200 72.300 506.000 72.400 ;
        RECT 508.400 72.300 509.200 72.400 ;
        RECT 490.800 71.700 509.200 72.300 ;
        RECT 490.800 71.600 491.600 71.700 ;
        RECT 503.600 71.600 504.400 71.700 ;
        RECT 505.200 71.600 506.000 71.700 ;
        RECT 508.400 71.600 509.200 71.700 ;
        RECT 9.200 70.300 10.000 70.400 ;
        RECT 12.400 70.300 13.200 70.400 ;
        RECT 9.200 69.700 13.200 70.300 ;
        RECT 9.200 69.600 10.000 69.700 ;
        RECT 12.400 69.600 13.200 69.700 ;
        RECT 22.000 70.300 22.800 70.400 ;
        RECT 26.800 70.300 27.600 70.400 ;
        RECT 22.000 69.700 27.600 70.300 ;
        RECT 22.000 69.600 22.800 69.700 ;
        RECT 26.800 69.600 27.600 69.700 ;
        RECT 28.400 70.300 29.200 70.400 ;
        RECT 46.000 70.300 46.800 70.400 ;
        RECT 28.400 69.700 46.800 70.300 ;
        RECT 28.400 69.600 29.200 69.700 ;
        RECT 46.000 69.600 46.800 69.700 ;
        RECT 49.200 70.300 50.000 70.400 ;
        RECT 54.000 70.300 54.800 70.400 ;
        RECT 49.200 69.700 54.800 70.300 ;
        RECT 49.200 69.600 50.000 69.700 ;
        RECT 54.000 69.600 54.800 69.700 ;
        RECT 78.000 70.300 78.800 70.400 ;
        RECT 87.600 70.300 88.400 70.400 ;
        RECT 116.400 70.300 117.200 70.400 ;
        RECT 130.800 70.300 131.600 70.400 ;
        RECT 78.000 69.700 131.600 70.300 ;
        RECT 78.000 69.600 78.800 69.700 ;
        RECT 87.600 69.600 88.400 69.700 ;
        RECT 116.400 69.600 117.200 69.700 ;
        RECT 130.800 69.600 131.600 69.700 ;
        RECT 196.400 70.300 197.200 70.400 ;
        RECT 210.800 70.300 211.600 70.400 ;
        RECT 217.200 70.300 218.000 70.400 ;
        RECT 196.400 69.700 218.000 70.300 ;
        RECT 196.400 69.600 197.200 69.700 ;
        RECT 210.800 69.600 211.600 69.700 ;
        RECT 217.200 69.600 218.000 69.700 ;
        RECT 273.200 70.300 274.000 70.400 ;
        RECT 308.400 70.300 309.200 70.400 ;
        RECT 273.200 69.700 309.200 70.300 ;
        RECT 273.200 69.600 274.000 69.700 ;
        RECT 308.400 69.600 309.200 69.700 ;
        RECT 310.000 70.300 310.800 70.400 ;
        RECT 314.800 70.300 315.600 70.400 ;
        RECT 310.000 69.700 315.600 70.300 ;
        RECT 310.000 69.600 310.800 69.700 ;
        RECT 314.800 69.600 315.600 69.700 ;
        RECT 369.200 70.300 370.000 70.400 ;
        RECT 374.000 70.300 374.800 70.400 ;
        RECT 388.400 70.300 389.200 70.400 ;
        RECT 369.200 69.700 389.200 70.300 ;
        RECT 369.200 69.600 370.000 69.700 ;
        RECT 374.000 69.600 374.800 69.700 ;
        RECT 388.400 69.600 389.200 69.700 ;
        RECT 446.000 70.300 446.800 70.400 ;
        RECT 454.000 70.300 454.800 70.400 ;
        RECT 446.000 69.700 454.800 70.300 ;
        RECT 446.000 69.600 446.800 69.700 ;
        RECT 454.000 69.600 454.800 69.700 ;
        RECT 460.400 70.300 461.200 70.400 ;
        RECT 490.800 70.300 491.600 70.400 ;
        RECT 460.400 69.700 491.600 70.300 ;
        RECT 460.400 69.600 461.200 69.700 ;
        RECT 490.800 69.600 491.600 69.700 ;
        RECT 492.400 70.300 493.200 70.400 ;
        RECT 497.200 70.300 498.000 70.400 ;
        RECT 492.400 69.700 498.000 70.300 ;
        RECT 492.400 69.600 493.200 69.700 ;
        RECT 497.200 69.600 498.000 69.700 ;
        RECT 500.400 70.300 501.200 70.400 ;
        RECT 510.000 70.300 510.800 70.400 ;
        RECT 500.400 69.700 510.800 70.300 ;
        RECT 500.400 69.600 501.200 69.700 ;
        RECT 510.000 69.600 510.800 69.700 ;
        RECT 6.000 68.300 6.800 68.400 ;
        RECT 30.000 68.300 30.800 68.400 ;
        RECT 6.000 67.700 30.800 68.300 ;
        RECT 6.000 67.600 6.800 67.700 ;
        RECT 30.000 67.600 30.800 67.700 ;
        RECT 31.600 68.300 32.400 68.400 ;
        RECT 42.800 68.300 43.600 68.400 ;
        RECT 31.600 67.700 43.600 68.300 ;
        RECT 31.600 67.600 32.400 67.700 ;
        RECT 42.800 67.600 43.600 67.700 ;
        RECT 62.000 68.300 62.800 68.400 ;
        RECT 74.800 68.300 75.600 68.400 ;
        RECT 62.000 67.700 75.600 68.300 ;
        RECT 62.000 67.600 62.800 67.700 ;
        RECT 74.800 67.600 75.600 67.700 ;
        RECT 111.600 68.300 112.400 68.400 ;
        RECT 134.000 68.300 134.800 68.400 ;
        RECT 111.600 67.700 134.800 68.300 ;
        RECT 111.600 67.600 112.400 67.700 ;
        RECT 134.000 67.600 134.800 67.700 ;
        RECT 153.200 68.300 154.000 68.400 ;
        RECT 159.600 68.300 160.400 68.400 ;
        RECT 153.200 67.700 160.400 68.300 ;
        RECT 153.200 67.600 154.000 67.700 ;
        RECT 159.600 67.600 160.400 67.700 ;
        RECT 327.600 68.300 328.400 68.400 ;
        RECT 380.400 68.300 381.200 68.400 ;
        RECT 327.600 67.700 381.200 68.300 ;
        RECT 327.600 67.600 328.400 67.700 ;
        RECT 380.400 67.600 381.200 67.700 ;
        RECT 386.800 68.300 387.600 68.400 ;
        RECT 393.200 68.300 394.000 68.400 ;
        RECT 386.800 67.700 394.000 68.300 ;
        RECT 386.800 67.600 387.600 67.700 ;
        RECT 393.200 67.600 394.000 67.700 ;
        RECT 399.600 68.300 400.400 68.400 ;
        RECT 458.800 68.300 459.600 68.400 ;
        RECT 399.600 67.700 459.600 68.300 ;
        RECT 399.600 67.600 400.400 67.700 ;
        RECT 458.800 67.600 459.600 67.700 ;
        RECT 465.200 68.300 466.000 68.400 ;
        RECT 474.800 68.300 475.600 68.400 ;
        RECT 465.200 67.700 475.600 68.300 ;
        RECT 465.200 67.600 466.000 67.700 ;
        RECT 474.800 67.600 475.600 67.700 ;
        RECT 482.800 68.300 483.600 68.400 ;
        RECT 502.000 68.300 502.800 68.400 ;
        RECT 482.800 67.700 502.800 68.300 ;
        RECT 482.800 67.600 483.600 67.700 ;
        RECT 502.000 67.600 502.800 67.700 ;
        RECT 510.000 68.300 510.800 68.400 ;
        RECT 516.400 68.300 517.200 68.400 ;
        RECT 510.000 67.700 517.200 68.300 ;
        RECT 510.000 67.600 510.800 67.700 ;
        RECT 516.400 67.600 517.200 67.700 ;
        RECT 2.800 66.300 3.600 66.400 ;
        RECT 18.800 66.300 19.600 66.400 ;
        RECT 2.800 65.700 19.600 66.300 ;
        RECT 2.800 65.600 3.600 65.700 ;
        RECT 18.800 65.600 19.600 65.700 ;
        RECT 34.800 66.300 35.600 66.400 ;
        RECT 39.600 66.300 40.400 66.400 ;
        RECT 34.800 65.700 40.400 66.300 ;
        RECT 34.800 65.600 35.600 65.700 ;
        RECT 39.600 65.600 40.400 65.700 ;
        RECT 87.600 66.300 88.400 66.400 ;
        RECT 108.400 66.300 109.200 66.400 ;
        RECT 150.000 66.300 150.800 66.400 ;
        RECT 164.400 66.300 165.200 66.400 ;
        RECT 188.400 66.300 189.200 66.400 ;
        RECT 198.000 66.300 198.800 66.400 ;
        RECT 225.200 66.300 226.000 66.400 ;
        RECT 87.600 65.700 226.000 66.300 ;
        RECT 87.600 65.600 88.400 65.700 ;
        RECT 108.400 65.600 109.200 65.700 ;
        RECT 150.000 65.600 150.800 65.700 ;
        RECT 164.400 65.600 165.200 65.700 ;
        RECT 188.400 65.600 189.200 65.700 ;
        RECT 198.000 65.600 198.800 65.700 ;
        RECT 225.200 65.600 226.000 65.700 ;
        RECT 242.800 66.300 243.600 66.400 ;
        RECT 262.000 66.300 262.800 66.400 ;
        RECT 242.800 65.700 262.800 66.300 ;
        RECT 242.800 65.600 243.600 65.700 ;
        RECT 262.000 65.600 262.800 65.700 ;
        RECT 263.600 66.300 264.400 66.400 ;
        RECT 266.800 66.300 267.600 66.400 ;
        RECT 263.600 65.700 267.600 66.300 ;
        RECT 263.600 65.600 264.400 65.700 ;
        RECT 266.800 65.600 267.600 65.700 ;
        RECT 294.000 66.300 294.800 66.400 ;
        RECT 311.600 66.300 312.400 66.400 ;
        RECT 294.000 65.700 312.400 66.300 ;
        RECT 294.000 65.600 294.800 65.700 ;
        RECT 311.600 65.600 312.400 65.700 ;
        RECT 319.600 66.300 320.400 66.400 ;
        RECT 324.400 66.300 325.200 66.400 ;
        RECT 319.600 65.700 325.200 66.300 ;
        RECT 319.600 65.600 320.400 65.700 ;
        RECT 324.400 65.600 325.200 65.700 ;
        RECT 449.200 66.300 450.000 66.400 ;
        RECT 458.800 66.300 459.600 66.400 ;
        RECT 449.200 65.700 459.600 66.300 ;
        RECT 449.200 65.600 450.000 65.700 ;
        RECT 458.800 65.600 459.600 65.700 ;
        RECT 503.600 66.300 504.400 66.400 ;
        RECT 535.600 66.300 536.400 66.400 ;
        RECT 503.600 65.700 536.400 66.300 ;
        RECT 503.600 65.600 504.400 65.700 ;
        RECT 535.600 65.600 536.400 65.700 ;
        RECT 25.200 64.300 26.000 64.400 ;
        RECT 36.400 64.300 37.200 64.400 ;
        RECT 25.200 63.700 37.200 64.300 ;
        RECT 25.200 63.600 26.000 63.700 ;
        RECT 36.400 63.600 37.200 63.700 ;
        RECT 38.000 64.300 38.800 64.400 ;
        RECT 44.400 64.300 45.200 64.400 ;
        RECT 38.000 63.700 45.200 64.300 ;
        RECT 38.000 63.600 38.800 63.700 ;
        RECT 44.400 63.600 45.200 63.700 ;
        RECT 255.600 64.300 256.400 64.400 ;
        RECT 294.000 64.300 294.800 64.400 ;
        RECT 255.600 63.700 294.800 64.300 ;
        RECT 255.600 63.600 256.400 63.700 ;
        RECT 294.000 63.600 294.800 63.700 ;
        RECT 303.600 64.300 304.400 64.400 ;
        RECT 321.200 64.300 322.000 64.400 ;
        RECT 303.600 63.700 322.000 64.300 ;
        RECT 303.600 63.600 304.400 63.700 ;
        RECT 321.200 63.600 322.000 63.700 ;
        RECT 335.600 64.300 336.400 64.400 ;
        RECT 354.800 64.300 355.600 64.400 ;
        RECT 335.600 63.700 355.600 64.300 ;
        RECT 335.600 63.600 336.400 63.700 ;
        RECT 354.800 63.600 355.600 63.700 ;
        RECT 394.800 64.300 395.600 64.400 ;
        RECT 404.400 64.300 405.200 64.400 ;
        RECT 394.800 63.700 405.200 64.300 ;
        RECT 394.800 63.600 395.600 63.700 ;
        RECT 404.400 63.600 405.200 63.700 ;
        RECT 447.600 64.300 448.400 64.400 ;
        RECT 450.800 64.300 451.600 64.400 ;
        RECT 447.600 63.700 451.600 64.300 ;
        RECT 447.600 63.600 448.400 63.700 ;
        RECT 450.800 63.600 451.600 63.700 ;
        RECT 455.600 64.300 456.400 64.400 ;
        RECT 479.600 64.300 480.400 64.400 ;
        RECT 455.600 63.700 480.400 64.300 ;
        RECT 455.600 63.600 456.400 63.700 ;
        RECT 479.600 63.600 480.400 63.700 ;
        RECT 30.000 62.300 30.800 62.400 ;
        RECT 34.800 62.300 35.600 62.400 ;
        RECT 30.000 61.700 35.600 62.300 ;
        RECT 30.000 61.600 30.800 61.700 ;
        RECT 34.800 61.600 35.600 61.700 ;
        RECT 148.400 61.600 149.200 62.400 ;
        RECT 337.200 62.300 338.000 62.400 ;
        RECT 343.600 62.300 344.400 62.400 ;
        RECT 367.600 62.300 368.400 62.400 ;
        RECT 377.200 62.300 378.000 62.400 ;
        RECT 337.200 61.700 378.000 62.300 ;
        RECT 337.200 61.600 338.000 61.700 ;
        RECT 343.600 61.600 344.400 61.700 ;
        RECT 367.600 61.600 368.400 61.700 ;
        RECT 377.200 61.600 378.000 61.700 ;
        RECT 380.400 62.300 381.200 62.400 ;
        RECT 450.800 62.300 451.600 62.400 ;
        RECT 454.000 62.300 454.800 62.400 ;
        RECT 380.400 61.700 449.900 62.300 ;
        RECT 380.400 61.600 381.200 61.700 ;
        RECT 49.200 60.300 50.000 60.400 ;
        RECT 55.600 60.300 56.400 60.400 ;
        RECT 49.200 59.700 56.400 60.300 ;
        RECT 49.200 59.600 50.000 59.700 ;
        RECT 55.600 59.600 56.400 59.700 ;
        RECT 132.400 60.300 133.200 60.400 ;
        RECT 214.000 60.300 214.800 60.400 ;
        RECT 218.800 60.300 219.600 60.400 ;
        RECT 230.000 60.300 230.800 60.400 ;
        RECT 249.200 60.300 250.000 60.400 ;
        RECT 132.400 59.700 171.500 60.300 ;
        RECT 132.400 59.600 133.200 59.700 ;
        RECT 170.900 58.400 171.500 59.700 ;
        RECT 214.000 59.700 250.000 60.300 ;
        RECT 214.000 59.600 214.800 59.700 ;
        RECT 218.800 59.600 219.600 59.700 ;
        RECT 230.000 59.600 230.800 59.700 ;
        RECT 249.200 59.600 250.000 59.700 ;
        RECT 290.800 60.300 291.600 60.400 ;
        RECT 297.200 60.300 298.000 60.400 ;
        RECT 290.800 59.700 298.000 60.300 ;
        RECT 290.800 59.600 291.600 59.700 ;
        RECT 297.200 59.600 298.000 59.700 ;
        RECT 327.600 60.300 328.400 60.400 ;
        RECT 385.200 60.300 386.000 60.400 ;
        RECT 391.600 60.300 392.400 60.400 ;
        RECT 327.600 59.700 384.300 60.300 ;
        RECT 327.600 59.600 328.400 59.700 ;
        RECT 10.800 58.300 11.600 58.400 ;
        RECT 22.000 58.300 22.800 58.400 ;
        RECT 10.800 57.700 22.800 58.300 ;
        RECT 10.800 57.600 11.600 57.700 ;
        RECT 22.000 57.600 22.800 57.700 ;
        RECT 81.200 58.300 82.000 58.400 ;
        RECT 138.800 58.300 139.600 58.400 ;
        RECT 169.200 58.300 170.000 58.400 ;
        RECT 81.200 57.700 170.000 58.300 ;
        RECT 81.200 57.600 82.000 57.700 ;
        RECT 138.800 57.600 139.600 57.700 ;
        RECT 169.200 57.600 170.000 57.700 ;
        RECT 170.800 58.300 171.600 58.400 ;
        RECT 242.800 58.300 243.600 58.400 ;
        RECT 170.800 57.700 243.600 58.300 ;
        RECT 170.800 57.600 171.600 57.700 ;
        RECT 242.800 57.600 243.600 57.700 ;
        RECT 332.400 58.300 333.200 58.400 ;
        RECT 367.600 58.300 368.400 58.400 ;
        RECT 332.400 57.700 368.400 58.300 ;
        RECT 383.700 58.300 384.300 59.700 ;
        RECT 385.200 59.700 392.400 60.300 ;
        RECT 449.300 60.300 449.900 61.700 ;
        RECT 450.800 61.700 454.800 62.300 ;
        RECT 450.800 61.600 451.600 61.700 ;
        RECT 454.000 61.600 454.800 61.700 ;
        RECT 468.400 61.600 469.200 62.400 ;
        RECT 460.400 60.300 461.200 60.400 ;
        RECT 449.300 59.700 461.200 60.300 ;
        RECT 385.200 59.600 386.000 59.700 ;
        RECT 391.600 59.600 392.400 59.700 ;
        RECT 460.400 59.600 461.200 59.700 ;
        RECT 466.800 60.300 467.600 60.400 ;
        RECT 487.600 60.300 488.400 60.400 ;
        RECT 466.800 59.700 488.400 60.300 ;
        RECT 466.800 59.600 467.600 59.700 ;
        RECT 487.600 59.600 488.400 59.700 ;
        RECT 471.600 58.300 472.400 58.400 ;
        RECT 383.700 57.700 472.400 58.300 ;
        RECT 332.400 57.600 333.200 57.700 ;
        RECT 367.600 57.600 368.400 57.700 ;
        RECT 471.600 57.600 472.400 57.700 ;
        RECT 494.000 58.300 494.800 58.400 ;
        RECT 500.400 58.300 501.200 58.400 ;
        RECT 506.800 58.300 507.600 58.400 ;
        RECT 494.000 57.700 507.600 58.300 ;
        RECT 494.000 57.600 494.800 57.700 ;
        RECT 500.400 57.600 501.200 57.700 ;
        RECT 506.800 57.600 507.600 57.700 ;
        RECT 4.400 56.300 5.200 56.400 ;
        RECT 9.200 56.300 10.000 56.400 ;
        RECT 12.400 56.300 13.200 56.400 ;
        RECT 4.400 55.700 13.200 56.300 ;
        RECT 4.400 55.600 5.200 55.700 ;
        RECT 9.200 55.600 10.000 55.700 ;
        RECT 12.400 55.600 13.200 55.700 ;
        RECT 20.400 56.300 21.200 56.400 ;
        RECT 30.000 56.300 30.800 56.400 ;
        RECT 20.400 55.700 30.800 56.300 ;
        RECT 20.400 55.600 21.200 55.700 ;
        RECT 30.000 55.600 30.800 55.700 ;
        RECT 103.600 56.300 104.400 56.400 ;
        RECT 135.600 56.300 136.400 56.400 ;
        RECT 103.600 55.700 136.400 56.300 ;
        RECT 103.600 55.600 104.400 55.700 ;
        RECT 135.600 55.600 136.400 55.700 ;
        RECT 137.200 56.300 138.000 56.400 ;
        RECT 143.600 56.300 144.400 56.400 ;
        RECT 137.200 55.700 144.400 56.300 ;
        RECT 137.200 55.600 138.000 55.700 ;
        RECT 143.600 55.600 144.400 55.700 ;
        RECT 145.200 56.300 146.000 56.400 ;
        RECT 159.600 56.300 160.400 56.400 ;
        RECT 145.200 55.700 160.400 56.300 ;
        RECT 145.200 55.600 146.000 55.700 ;
        RECT 159.600 55.600 160.400 55.700 ;
        RECT 234.800 56.300 235.600 56.400 ;
        RECT 255.600 56.300 256.400 56.400 ;
        RECT 234.800 55.700 256.400 56.300 ;
        RECT 234.800 55.600 235.600 55.700 ;
        RECT 255.600 55.600 256.400 55.700 ;
        RECT 324.400 56.300 325.200 56.400 ;
        RECT 353.200 56.300 354.000 56.400 ;
        RECT 354.800 56.300 355.600 56.400 ;
        RECT 324.400 55.700 355.600 56.300 ;
        RECT 324.400 55.600 325.200 55.700 ;
        RECT 353.200 55.600 354.000 55.700 ;
        RECT 354.800 55.600 355.600 55.700 ;
        RECT 358.000 56.300 358.800 56.400 ;
        RECT 372.400 56.300 373.200 56.400 ;
        RECT 418.800 56.300 419.600 56.400 ;
        RECT 358.000 55.700 419.600 56.300 ;
        RECT 358.000 55.600 358.800 55.700 ;
        RECT 372.400 55.600 373.200 55.700 ;
        RECT 418.800 55.600 419.600 55.700 ;
        RECT 420.400 56.300 421.200 56.400 ;
        RECT 433.200 56.300 434.000 56.400 ;
        RECT 462.000 56.300 462.800 56.400 ;
        RECT 420.400 55.700 434.000 56.300 ;
        RECT 420.400 55.600 421.200 55.700 ;
        RECT 433.200 55.600 434.000 55.700 ;
        RECT 434.900 55.700 462.800 56.300 ;
        RECT 1.200 54.300 2.000 54.400 ;
        RECT 2.800 54.300 3.600 54.400 ;
        RECT 4.400 54.300 5.200 54.400 ;
        RECT 1.200 53.700 5.200 54.300 ;
        RECT 1.200 53.600 2.000 53.700 ;
        RECT 2.800 53.600 3.600 53.700 ;
        RECT 4.400 53.600 5.200 53.700 ;
        RECT 10.800 54.300 11.600 54.400 ;
        RECT 17.200 54.300 18.000 54.400 ;
        RECT 10.800 53.700 18.000 54.300 ;
        RECT 10.800 53.600 11.600 53.700 ;
        RECT 17.200 53.600 18.000 53.700 ;
        RECT 23.600 54.300 24.400 54.400 ;
        RECT 31.600 54.300 32.400 54.400 ;
        RECT 46.000 54.300 46.800 54.400 ;
        RECT 23.600 53.700 46.800 54.300 ;
        RECT 23.600 53.600 24.400 53.700 ;
        RECT 31.600 53.600 32.400 53.700 ;
        RECT 46.000 53.600 46.800 53.700 ;
        RECT 130.800 54.300 131.600 54.400 ;
        RECT 162.800 54.300 163.600 54.400 ;
        RECT 174.000 54.300 174.800 54.400 ;
        RECT 202.800 54.300 203.600 54.400 ;
        RECT 247.600 54.300 248.400 54.400 ;
        RECT 308.400 54.300 309.200 54.400 ;
        RECT 130.800 53.700 309.200 54.300 ;
        RECT 130.800 53.600 131.600 53.700 ;
        RECT 162.800 53.600 163.600 53.700 ;
        RECT 174.000 53.600 174.800 53.700 ;
        RECT 202.800 53.600 203.600 53.700 ;
        RECT 247.600 53.600 248.400 53.700 ;
        RECT 308.400 53.600 309.200 53.700 ;
        RECT 318.000 54.300 318.800 54.400 ;
        RECT 358.000 54.300 358.800 54.400 ;
        RECT 369.200 54.300 370.000 54.400 ;
        RECT 318.000 53.700 370.000 54.300 ;
        RECT 318.000 53.600 318.800 53.700 ;
        RECT 358.000 53.600 358.800 53.700 ;
        RECT 369.200 53.600 370.000 53.700 ;
        RECT 386.800 54.300 387.600 54.400 ;
        RECT 407.600 54.300 408.400 54.400 ;
        RECT 386.800 53.700 408.400 54.300 ;
        RECT 386.800 53.600 387.600 53.700 ;
        RECT 407.600 53.600 408.400 53.700 ;
        RECT 410.800 54.300 411.600 54.400 ;
        RECT 425.200 54.300 426.000 54.400 ;
        RECT 410.800 53.700 426.000 54.300 ;
        RECT 410.800 53.600 411.600 53.700 ;
        RECT 425.200 53.600 426.000 53.700 ;
        RECT 430.000 54.300 430.800 54.400 ;
        RECT 434.900 54.300 435.500 55.700 ;
        RECT 462.000 55.600 462.800 55.700 ;
        RECT 476.400 56.300 477.200 56.400 ;
        RECT 492.400 56.300 493.200 56.400 ;
        RECT 514.800 56.300 515.600 56.400 ;
        RECT 476.400 55.700 515.600 56.300 ;
        RECT 476.400 55.600 477.200 55.700 ;
        RECT 492.400 55.600 493.200 55.700 ;
        RECT 514.800 55.600 515.600 55.700 ;
        RECT 476.400 54.300 477.200 54.400 ;
        RECT 430.000 53.700 435.500 54.300 ;
        RECT 441.300 53.700 477.200 54.300 ;
        RECT 430.000 53.600 430.800 53.700 ;
        RECT 18.800 52.300 19.600 52.400 ;
        RECT 26.800 52.300 27.600 52.400 ;
        RECT 18.800 51.700 27.600 52.300 ;
        RECT 18.800 51.600 19.600 51.700 ;
        RECT 26.800 51.600 27.600 51.700 ;
        RECT 122.800 52.300 123.600 52.400 ;
        RECT 145.200 52.300 146.000 52.400 ;
        RECT 154.800 52.300 155.600 52.400 ;
        RECT 122.800 51.700 155.600 52.300 ;
        RECT 122.800 51.600 123.600 51.700 ;
        RECT 145.200 51.600 146.000 51.700 ;
        RECT 154.800 51.600 155.600 51.700 ;
        RECT 158.000 52.300 158.800 52.400 ;
        RECT 161.200 52.300 162.000 52.400 ;
        RECT 162.800 52.300 163.600 52.400 ;
        RECT 158.000 51.700 163.600 52.300 ;
        RECT 158.000 51.600 158.800 51.700 ;
        RECT 161.200 51.600 162.000 51.700 ;
        RECT 162.800 51.600 163.600 51.700 ;
        RECT 190.000 52.300 190.800 52.400 ;
        RECT 215.600 52.300 216.400 52.400 ;
        RECT 190.000 51.700 216.400 52.300 ;
        RECT 190.000 51.600 190.800 51.700 ;
        RECT 215.600 51.600 216.400 51.700 ;
        RECT 222.000 52.300 222.800 52.400 ;
        RECT 226.800 52.300 227.600 52.400 ;
        RECT 236.400 52.300 237.200 52.400 ;
        RECT 222.000 51.700 237.200 52.300 ;
        RECT 222.000 51.600 222.800 51.700 ;
        RECT 226.800 51.600 227.600 51.700 ;
        RECT 236.400 51.600 237.200 51.700 ;
        RECT 354.800 52.300 355.600 52.400 ;
        RECT 359.600 52.300 360.400 52.400 ;
        RECT 362.800 52.300 363.600 52.400 ;
        RECT 354.800 51.700 363.600 52.300 ;
        RECT 354.800 51.600 355.600 51.700 ;
        RECT 359.600 51.600 360.400 51.700 ;
        RECT 362.800 51.600 363.600 51.700 ;
        RECT 364.400 52.300 365.200 52.400 ;
        RECT 369.200 52.300 370.000 52.400 ;
        RECT 364.400 51.700 370.000 52.300 ;
        RECT 364.400 51.600 365.200 51.700 ;
        RECT 369.200 51.600 370.000 51.700 ;
        RECT 412.400 52.300 413.200 52.400 ;
        RECT 417.200 52.300 418.000 52.400 ;
        RECT 412.400 51.700 418.000 52.300 ;
        RECT 412.400 51.600 413.200 51.700 ;
        RECT 417.200 51.600 418.000 51.700 ;
        RECT 418.800 52.300 419.600 52.400 ;
        RECT 441.300 52.300 441.900 53.700 ;
        RECT 476.400 53.600 477.200 53.700 ;
        RECT 497.200 54.300 498.000 54.400 ;
        RECT 502.000 54.300 502.800 54.400 ;
        RECT 497.200 53.700 502.800 54.300 ;
        RECT 497.200 53.600 498.000 53.700 ;
        RECT 502.000 53.600 502.800 53.700 ;
        RECT 511.600 54.300 512.400 54.400 ;
        RECT 534.000 54.300 534.800 54.400 ;
        RECT 511.600 53.700 534.800 54.300 ;
        RECT 511.600 53.600 512.400 53.700 ;
        RECT 534.000 53.600 534.800 53.700 ;
        RECT 418.800 51.700 441.900 52.300 ;
        RECT 418.800 51.600 419.600 51.700 ;
        RECT 442.800 51.600 443.600 52.400 ;
        RECT 449.200 52.300 450.000 52.400 ;
        RECT 482.800 52.300 483.600 52.400 ;
        RECT 449.200 51.700 483.600 52.300 ;
        RECT 449.200 51.600 450.000 51.700 ;
        RECT 482.800 51.600 483.600 51.700 ;
        RECT 484.400 52.300 485.200 52.400 ;
        RECT 508.400 52.300 509.200 52.400 ;
        RECT 484.400 51.700 509.200 52.300 ;
        RECT 484.400 51.600 485.200 51.700 ;
        RECT 508.400 51.600 509.200 51.700 ;
        RECT 510.000 52.300 510.800 52.400 ;
        RECT 534.000 52.300 534.800 52.400 ;
        RECT 510.000 51.700 534.800 52.300 ;
        RECT 510.000 51.600 510.800 51.700 ;
        RECT 534.000 51.600 534.800 51.700 ;
        RECT 4.400 50.300 5.200 50.400 ;
        RECT 15.600 50.300 16.400 50.400 ;
        RECT 25.200 50.300 26.000 50.400 ;
        RECT 4.400 49.700 26.000 50.300 ;
        RECT 4.400 49.600 5.200 49.700 ;
        RECT 15.600 49.600 16.400 49.700 ;
        RECT 25.200 49.600 26.000 49.700 ;
        RECT 134.000 50.300 134.800 50.400 ;
        RECT 148.400 50.300 149.200 50.400 ;
        RECT 134.000 49.700 149.200 50.300 ;
        RECT 134.000 49.600 134.800 49.700 ;
        RECT 148.400 49.600 149.200 49.700 ;
        RECT 177.200 50.300 178.000 50.400 ;
        RECT 180.400 50.300 181.200 50.400 ;
        RECT 177.200 49.700 181.200 50.300 ;
        RECT 177.200 49.600 178.000 49.700 ;
        RECT 180.400 49.600 181.200 49.700 ;
        RECT 225.200 50.300 226.000 50.400 ;
        RECT 233.200 50.300 234.000 50.400 ;
        RECT 225.200 49.700 234.000 50.300 ;
        RECT 225.200 49.600 226.000 49.700 ;
        RECT 233.200 49.600 234.000 49.700 ;
        RECT 239.600 50.300 240.400 50.400 ;
        RECT 262.000 50.300 262.800 50.400 ;
        RECT 279.600 50.300 280.400 50.400 ;
        RECT 284.400 50.300 285.200 50.400 ;
        RECT 314.800 50.300 315.600 50.400 ;
        RECT 239.600 49.700 315.600 50.300 ;
        RECT 239.600 49.600 240.400 49.700 ;
        RECT 262.000 49.600 262.800 49.700 ;
        RECT 279.600 49.600 280.400 49.700 ;
        RECT 284.400 49.600 285.200 49.700 ;
        RECT 314.800 49.600 315.600 49.700 ;
        RECT 369.200 50.300 370.000 50.400 ;
        RECT 436.400 50.300 437.200 50.400 ;
        RECT 369.200 49.700 437.200 50.300 ;
        RECT 369.200 49.600 370.000 49.700 ;
        RECT 436.400 49.600 437.200 49.700 ;
        RECT 521.200 50.300 522.000 50.400 ;
        RECT 530.800 50.300 531.600 50.400 ;
        RECT 546.800 50.300 547.600 50.400 ;
        RECT 521.200 49.700 547.600 50.300 ;
        RECT 521.200 49.600 522.000 49.700 ;
        RECT 530.800 49.600 531.600 49.700 ;
        RECT 546.800 49.600 547.600 49.700 ;
        RECT 415.600 48.300 416.400 48.400 ;
        RECT 418.800 48.300 419.600 48.400 ;
        RECT 415.600 47.700 419.600 48.300 ;
        RECT 415.600 47.600 416.400 47.700 ;
        RECT 418.800 47.600 419.600 47.700 ;
        RECT 430.000 48.300 430.800 48.400 ;
        RECT 447.600 48.300 448.400 48.400 ;
        RECT 430.000 47.700 448.400 48.300 ;
        RECT 430.000 47.600 430.800 47.700 ;
        RECT 447.600 47.600 448.400 47.700 ;
        RECT 433.200 46.300 434.000 46.400 ;
        RECT 478.000 46.300 478.800 46.400 ;
        RECT 433.200 45.700 478.800 46.300 ;
        RECT 433.200 45.600 434.000 45.700 ;
        RECT 478.000 45.600 478.800 45.700 ;
        RECT 503.600 46.300 504.400 46.400 ;
        RECT 506.800 46.300 507.600 46.400 ;
        RECT 503.600 45.700 507.600 46.300 ;
        RECT 503.600 45.600 504.400 45.700 ;
        RECT 506.800 45.600 507.600 45.700 ;
        RECT 54.000 44.300 54.800 44.400 ;
        RECT 57.200 44.300 58.000 44.400 ;
        RECT 54.000 43.700 58.000 44.300 ;
        RECT 54.000 43.600 54.800 43.700 ;
        RECT 57.200 43.600 58.000 43.700 ;
        RECT 497.200 43.600 498.000 44.400 ;
        RECT 166.000 42.300 166.800 42.400 ;
        RECT 169.200 42.300 170.000 42.400 ;
        RECT 166.000 41.700 170.000 42.300 ;
        RECT 166.000 41.600 166.800 41.700 ;
        RECT 169.200 41.600 170.000 41.700 ;
        RECT 185.200 42.300 186.000 42.400 ;
        RECT 193.200 42.300 194.000 42.400 ;
        RECT 185.200 41.700 194.000 42.300 ;
        RECT 185.200 41.600 186.000 41.700 ;
        RECT 193.200 41.600 194.000 41.700 ;
        RECT 247.600 42.300 248.400 42.400 ;
        RECT 252.400 42.300 253.200 42.400 ;
        RECT 247.600 41.700 253.200 42.300 ;
        RECT 247.600 41.600 248.400 41.700 ;
        RECT 252.400 41.600 253.200 41.700 ;
        RECT 465.200 42.300 466.000 42.400 ;
        RECT 468.400 42.300 469.200 42.400 ;
        RECT 465.200 41.700 469.200 42.300 ;
        RECT 465.200 41.600 466.000 41.700 ;
        RECT 468.400 41.600 469.200 41.700 ;
        RECT 22.000 40.300 22.800 40.400 ;
        RECT 26.800 40.300 27.600 40.400 ;
        RECT 22.000 39.700 27.600 40.300 ;
        RECT 22.000 39.600 22.800 39.700 ;
        RECT 26.800 39.600 27.600 39.700 ;
        RECT 162.800 40.300 163.600 40.400 ;
        RECT 166.000 40.300 166.800 40.400 ;
        RECT 178.800 40.300 179.600 40.400 ;
        RECT 162.800 39.700 179.600 40.300 ;
        RECT 162.800 39.600 163.600 39.700 ;
        RECT 166.000 39.600 166.800 39.700 ;
        RECT 178.800 39.600 179.600 39.700 ;
        RECT 180.400 40.300 181.200 40.400 ;
        RECT 194.800 40.300 195.600 40.400 ;
        RECT 180.400 39.700 195.600 40.300 ;
        RECT 180.400 39.600 181.200 39.700 ;
        RECT 194.800 39.600 195.600 39.700 ;
        RECT 20.400 37.600 21.200 38.400 ;
        RECT 482.800 38.300 483.600 38.400 ;
        RECT 487.600 38.300 488.400 38.400 ;
        RECT 482.800 37.700 488.400 38.300 ;
        RECT 482.800 37.600 483.600 37.700 ;
        RECT 487.600 37.600 488.400 37.700 ;
        RECT 519.600 37.600 520.400 38.400 ;
        RECT 530.800 38.300 531.600 38.400 ;
        RECT 532.400 38.300 533.200 38.400 ;
        RECT 530.800 37.700 533.200 38.300 ;
        RECT 530.800 37.600 531.600 37.700 ;
        RECT 532.400 37.600 533.200 37.700 ;
        RECT 135.600 34.300 136.400 34.400 ;
        RECT 407.600 34.300 408.400 34.400 ;
        RECT 135.600 33.700 408.400 34.300 ;
        RECT 135.600 33.600 136.400 33.700 ;
        RECT 407.600 33.600 408.400 33.700 ;
        RECT 476.400 34.300 477.200 34.400 ;
        RECT 479.600 34.300 480.400 34.400 ;
        RECT 476.400 33.700 480.400 34.300 ;
        RECT 476.400 33.600 477.200 33.700 ;
        RECT 479.600 33.600 480.400 33.700 ;
        RECT 527.600 34.300 528.400 34.400 ;
        RECT 542.000 34.300 542.800 34.400 ;
        RECT 527.600 33.700 542.800 34.300 ;
        RECT 527.600 33.600 528.400 33.700 ;
        RECT 542.000 33.600 542.800 33.700 ;
        RECT 207.600 32.300 208.400 32.400 ;
        RECT 218.800 32.300 219.600 32.400 ;
        RECT 207.600 31.700 219.600 32.300 ;
        RECT 207.600 31.600 208.400 31.700 ;
        RECT 218.800 31.600 219.600 31.700 ;
        RECT 222.000 32.300 222.800 32.400 ;
        RECT 226.800 32.300 227.600 32.400 ;
        RECT 222.000 31.700 227.600 32.300 ;
        RECT 222.000 31.600 222.800 31.700 ;
        RECT 226.800 31.600 227.600 31.700 ;
        RECT 487.600 32.300 488.400 32.400 ;
        RECT 518.000 32.300 518.800 32.400 ;
        RECT 487.600 31.700 518.800 32.300 ;
        RECT 487.600 31.600 488.400 31.700 ;
        RECT 518.000 31.600 518.800 31.700 ;
        RECT 522.800 32.300 523.600 32.400 ;
        RECT 532.400 32.300 533.200 32.400 ;
        RECT 522.800 31.700 533.200 32.300 ;
        RECT 522.800 31.600 523.600 31.700 ;
        RECT 532.400 31.600 533.200 31.700 ;
        RECT 31.600 30.300 32.400 30.400 ;
        RECT 46.000 30.300 46.800 30.400 ;
        RECT 31.600 29.700 46.800 30.300 ;
        RECT 31.600 29.600 32.400 29.700 ;
        RECT 46.000 29.600 46.800 29.700 ;
        RECT 74.800 30.300 75.600 30.400 ;
        RECT 79.600 30.300 80.400 30.400 ;
        RECT 74.800 29.700 80.400 30.300 ;
        RECT 74.800 29.600 75.600 29.700 ;
        RECT 79.600 29.600 80.400 29.700 ;
        RECT 114.800 30.300 115.600 30.400 ;
        RECT 119.600 30.300 120.400 30.400 ;
        RECT 162.800 30.300 163.600 30.400 ;
        RECT 114.800 29.700 163.600 30.300 ;
        RECT 114.800 29.600 115.600 29.700 ;
        RECT 119.600 29.600 120.400 29.700 ;
        RECT 162.800 29.600 163.600 29.700 ;
        RECT 212.400 30.300 213.200 30.400 ;
        RECT 222.000 30.300 222.800 30.400 ;
        RECT 212.400 29.700 222.800 30.300 ;
        RECT 212.400 29.600 213.200 29.700 ;
        RECT 222.000 29.600 222.800 29.700 ;
        RECT 270.000 30.300 270.800 30.400 ;
        RECT 281.200 30.300 282.000 30.400 ;
        RECT 270.000 29.700 282.000 30.300 ;
        RECT 270.000 29.600 270.800 29.700 ;
        RECT 281.200 29.600 282.000 29.700 ;
        RECT 287.600 30.300 288.400 30.400 ;
        RECT 324.400 30.300 325.200 30.400 ;
        RECT 287.600 29.700 325.200 30.300 ;
        RECT 287.600 29.600 288.400 29.700 ;
        RECT 324.400 29.600 325.200 29.700 ;
        RECT 476.400 30.300 477.200 30.400 ;
        RECT 524.400 30.300 525.200 30.400 ;
        RECT 476.400 29.700 525.200 30.300 ;
        RECT 476.400 29.600 477.200 29.700 ;
        RECT 524.400 29.600 525.200 29.700 ;
        RECT 55.600 28.300 56.400 28.400 ;
        RECT 57.200 28.300 58.000 28.400 ;
        RECT 55.600 27.700 58.000 28.300 ;
        RECT 55.600 27.600 56.400 27.700 ;
        RECT 57.200 27.600 58.000 27.700 ;
        RECT 188.400 28.300 189.200 28.400 ;
        RECT 204.400 28.300 205.200 28.400 ;
        RECT 188.400 27.700 205.200 28.300 ;
        RECT 188.400 27.600 189.200 27.700 ;
        RECT 204.400 27.600 205.200 27.700 ;
        RECT 270.000 28.300 270.800 28.400 ;
        RECT 279.600 28.300 280.400 28.400 ;
        RECT 286.000 28.300 286.800 28.400 ;
        RECT 270.000 27.700 286.800 28.300 ;
        RECT 270.000 27.600 270.800 27.700 ;
        RECT 279.600 27.600 280.400 27.700 ;
        RECT 286.000 27.600 286.800 27.700 ;
        RECT 287.600 28.300 288.400 28.400 ;
        RECT 308.400 28.300 309.200 28.400 ;
        RECT 287.600 27.700 309.200 28.300 ;
        RECT 287.600 27.600 288.400 27.700 ;
        RECT 308.400 27.600 309.200 27.700 ;
        RECT 385.200 27.600 386.000 28.400 ;
        RECT 402.800 28.300 403.600 28.400 ;
        RECT 518.000 28.300 518.800 28.400 ;
        RECT 402.800 27.700 518.800 28.300 ;
        RECT 402.800 27.600 403.600 27.700 ;
        RECT 518.000 27.600 518.800 27.700 ;
        RECT 223.600 26.300 224.400 26.400 ;
        RECT 226.800 26.300 227.600 26.400 ;
        RECT 223.600 25.700 227.600 26.300 ;
        RECT 223.600 25.600 224.400 25.700 ;
        RECT 226.800 25.600 227.600 25.700 ;
        RECT 247.600 26.300 248.400 26.400 ;
        RECT 305.200 26.300 306.000 26.400 ;
        RECT 247.600 25.700 306.000 26.300 ;
        RECT 247.600 25.600 248.400 25.700 ;
        RECT 305.200 25.600 306.000 25.700 ;
        RECT 449.200 26.300 450.000 26.400 ;
        RECT 468.400 26.300 469.200 26.400 ;
        RECT 482.800 26.300 483.600 26.400 ;
        RECT 498.800 26.300 499.600 26.400 ;
        RECT 521.200 26.300 522.000 26.400 ;
        RECT 449.200 25.700 522.000 26.300 ;
        RECT 449.200 25.600 450.000 25.700 ;
        RECT 468.400 25.600 469.200 25.700 ;
        RECT 482.800 25.600 483.600 25.700 ;
        RECT 498.800 25.600 499.600 25.700 ;
        RECT 521.200 25.600 522.000 25.700 ;
        RECT 92.400 24.300 93.200 24.400 ;
        RECT 119.600 24.300 120.400 24.400 ;
        RECT 92.400 23.700 120.400 24.300 ;
        RECT 92.400 23.600 93.200 23.700 ;
        RECT 119.600 23.600 120.400 23.700 ;
        RECT 122.800 24.300 123.600 24.400 ;
        RECT 135.600 24.300 136.400 24.400 ;
        RECT 122.800 23.700 136.400 24.300 ;
        RECT 122.800 23.600 123.600 23.700 ;
        RECT 135.600 23.600 136.400 23.700 ;
        RECT 153.200 24.300 154.000 24.400 ;
        RECT 234.800 24.300 235.600 24.400 ;
        RECT 153.200 23.700 235.600 24.300 ;
        RECT 153.200 23.600 154.000 23.700 ;
        RECT 234.800 23.600 235.600 23.700 ;
        RECT 250.800 24.300 251.600 24.400 ;
        RECT 271.600 24.300 272.400 24.400 ;
        RECT 250.800 23.700 272.400 24.300 ;
        RECT 250.800 23.600 251.600 23.700 ;
        RECT 271.600 23.600 272.400 23.700 ;
        RECT 471.600 24.300 472.400 24.400 ;
        RECT 497.200 24.300 498.000 24.400 ;
        RECT 498.800 24.300 499.600 24.400 ;
        RECT 471.600 23.700 499.600 24.300 ;
        RECT 471.600 23.600 472.400 23.700 ;
        RECT 497.200 23.600 498.000 23.700 ;
        RECT 498.800 23.600 499.600 23.700 ;
        RECT 500.400 24.300 501.200 24.400 ;
        RECT 502.000 24.300 502.800 24.400 ;
        RECT 500.400 23.700 502.800 24.300 ;
        RECT 500.400 23.600 501.200 23.700 ;
        RECT 502.000 23.600 502.800 23.700 ;
        RECT 60.400 22.300 61.200 22.400 ;
        RECT 66.800 22.300 67.600 22.400 ;
        RECT 90.800 22.300 91.600 22.400 ;
        RECT 94.000 22.300 94.800 22.400 ;
        RECT 60.400 21.700 94.800 22.300 ;
        RECT 60.400 21.600 61.200 21.700 ;
        RECT 66.800 21.600 67.600 21.700 ;
        RECT 90.800 21.600 91.600 21.700 ;
        RECT 94.000 21.600 94.800 21.700 ;
        RECT 100.400 22.300 101.200 22.400 ;
        RECT 106.800 22.300 107.600 22.400 ;
        RECT 150.000 22.300 150.800 22.400 ;
        RECT 154.800 22.300 155.600 22.400 ;
        RECT 185.200 22.300 186.000 22.400 ;
        RECT 198.000 22.300 198.800 22.400 ;
        RECT 100.400 21.700 198.800 22.300 ;
        RECT 100.400 21.600 101.200 21.700 ;
        RECT 106.800 21.600 107.600 21.700 ;
        RECT 150.000 21.600 150.800 21.700 ;
        RECT 154.800 21.600 155.600 21.700 ;
        RECT 185.200 21.600 186.000 21.700 ;
        RECT 198.000 21.600 198.800 21.700 ;
        RECT 202.800 22.300 203.600 22.400 ;
        RECT 233.200 22.300 234.000 22.400 ;
        RECT 202.800 21.700 234.000 22.300 ;
        RECT 202.800 21.600 203.600 21.700 ;
        RECT 233.200 21.600 234.000 21.700 ;
        RECT 244.400 22.300 245.200 22.400 ;
        RECT 270.000 22.300 270.800 22.400 ;
        RECT 244.400 21.700 270.800 22.300 ;
        RECT 244.400 21.600 245.200 21.700 ;
        RECT 270.000 21.600 270.800 21.700 ;
        RECT 335.600 22.300 336.400 22.400 ;
        RECT 343.600 22.300 344.400 22.400 ;
        RECT 335.600 21.700 344.400 22.300 ;
        RECT 335.600 21.600 336.400 21.700 ;
        RECT 343.600 21.600 344.400 21.700 ;
        RECT 367.600 22.300 368.400 22.400 ;
        RECT 377.200 22.300 378.000 22.400 ;
        RECT 367.600 21.700 378.000 22.300 ;
        RECT 367.600 21.600 368.400 21.700 ;
        RECT 377.200 21.600 378.000 21.700 ;
        RECT 390.000 22.300 390.800 22.400 ;
        RECT 398.000 22.300 398.800 22.400 ;
        RECT 390.000 21.700 398.800 22.300 ;
        RECT 390.000 21.600 390.800 21.700 ;
        RECT 398.000 21.600 398.800 21.700 ;
        RECT 428.400 22.300 429.200 22.400 ;
        RECT 433.200 22.300 434.000 22.400 ;
        RECT 428.400 21.700 434.000 22.300 ;
        RECT 428.400 21.600 429.200 21.700 ;
        RECT 433.200 21.600 434.000 21.700 ;
        RECT 503.600 21.600 504.400 22.400 ;
        RECT 2.800 20.300 3.600 20.400 ;
        RECT 9.200 20.300 10.000 20.400 ;
        RECT 2.800 19.700 10.000 20.300 ;
        RECT 2.800 19.600 3.600 19.700 ;
        RECT 9.200 19.600 10.000 19.700 ;
        RECT 103.600 20.300 104.400 20.400 ;
        RECT 121.200 20.300 122.000 20.400 ;
        RECT 103.600 19.700 122.000 20.300 ;
        RECT 103.600 19.600 104.400 19.700 ;
        RECT 121.200 19.600 122.000 19.700 ;
        RECT 262.000 20.300 262.800 20.400 ;
        RECT 266.800 20.300 267.600 20.400 ;
        RECT 262.000 19.700 267.600 20.300 ;
        RECT 262.000 19.600 262.800 19.700 ;
        RECT 266.800 19.600 267.600 19.700 ;
        RECT 306.800 20.300 307.600 20.400 ;
        RECT 340.400 20.300 341.200 20.400 ;
        RECT 354.800 20.300 355.600 20.400 ;
        RECT 359.600 20.300 360.400 20.400 ;
        RECT 386.800 20.300 387.600 20.400 ;
        RECT 306.800 19.700 387.600 20.300 ;
        RECT 306.800 19.600 307.600 19.700 ;
        RECT 340.400 19.600 341.200 19.700 ;
        RECT 354.800 19.600 355.600 19.700 ;
        RECT 359.600 19.600 360.400 19.700 ;
        RECT 386.800 19.600 387.600 19.700 ;
        RECT 231.600 18.300 232.400 18.400 ;
        RECT 238.000 18.300 238.800 18.400 ;
        RECT 246.000 18.300 246.800 18.400 ;
        RECT 265.200 18.300 266.000 18.400 ;
        RECT 231.600 17.700 266.000 18.300 ;
        RECT 231.600 17.600 232.400 17.700 ;
        RECT 238.000 17.600 238.800 17.700 ;
        RECT 246.000 17.600 246.800 17.700 ;
        RECT 265.200 17.600 266.000 17.700 ;
        RECT 266.800 18.300 267.600 18.400 ;
        RECT 289.200 18.300 290.000 18.400 ;
        RECT 266.800 17.700 290.000 18.300 ;
        RECT 266.800 17.600 267.600 17.700 ;
        RECT 289.200 17.600 290.000 17.700 ;
        RECT 18.800 16.300 19.600 16.400 ;
        RECT 52.400 16.300 53.200 16.400 ;
        RECT 87.600 16.300 88.400 16.400 ;
        RECT 100.400 16.300 101.200 16.400 ;
        RECT 18.800 15.700 101.200 16.300 ;
        RECT 18.800 15.600 19.600 15.700 ;
        RECT 52.400 15.600 53.200 15.700 ;
        RECT 87.600 15.600 88.400 15.700 ;
        RECT 100.400 15.600 101.200 15.700 ;
        RECT 239.600 16.300 240.400 16.400 ;
        RECT 266.800 16.300 267.600 16.400 ;
        RECT 239.600 15.700 267.600 16.300 ;
        RECT 239.600 15.600 240.400 15.700 ;
        RECT 266.800 15.600 267.600 15.700 ;
        RECT 386.800 16.300 387.600 16.400 ;
        RECT 412.400 16.300 413.200 16.400 ;
        RECT 433.200 16.300 434.000 16.400 ;
        RECT 386.800 15.700 434.000 16.300 ;
        RECT 386.800 15.600 387.600 15.700 ;
        RECT 412.400 15.600 413.200 15.700 ;
        RECT 433.200 15.600 434.000 15.700 ;
        RECT 20.400 14.300 21.200 14.400 ;
        RECT 22.000 14.300 22.800 14.400 ;
        RECT 20.400 13.700 22.800 14.300 ;
        RECT 20.400 13.600 21.200 13.700 ;
        RECT 22.000 13.600 22.800 13.700 ;
        RECT 49.200 14.300 50.000 14.400 ;
        RECT 70.000 14.300 70.800 14.400 ;
        RECT 49.200 13.700 70.800 14.300 ;
        RECT 49.200 13.600 50.000 13.700 ;
        RECT 70.000 13.600 70.800 13.700 ;
        RECT 82.800 14.300 83.600 14.400 ;
        RECT 97.200 14.300 98.000 14.400 ;
        RECT 82.800 13.700 98.000 14.300 ;
        RECT 82.800 13.600 83.600 13.700 ;
        RECT 97.200 13.600 98.000 13.700 ;
        RECT 142.000 14.300 142.800 14.400 ;
        RECT 158.000 14.300 158.800 14.400 ;
        RECT 142.000 13.700 158.800 14.300 ;
        RECT 142.000 13.600 142.800 13.700 ;
        RECT 158.000 13.600 158.800 13.700 ;
        RECT 194.800 14.300 195.600 14.400 ;
        RECT 223.600 14.300 224.400 14.400 ;
        RECT 194.800 13.700 224.400 14.300 ;
        RECT 194.800 13.600 195.600 13.700 ;
        RECT 223.600 13.600 224.400 13.700 ;
        RECT 226.800 14.300 227.600 14.400 ;
        RECT 244.400 14.300 245.200 14.400 ;
        RECT 226.800 13.700 245.200 14.300 ;
        RECT 226.800 13.600 227.600 13.700 ;
        RECT 244.400 13.600 245.200 13.700 ;
        RECT 255.600 14.300 256.400 14.400 ;
        RECT 257.200 14.300 258.000 14.400 ;
        RECT 263.600 14.300 264.400 14.400 ;
        RECT 255.600 13.700 264.400 14.300 ;
        RECT 255.600 13.600 256.400 13.700 ;
        RECT 257.200 13.600 258.000 13.700 ;
        RECT 263.600 13.600 264.400 13.700 ;
        RECT 268.400 14.300 269.200 14.400 ;
        RECT 279.600 14.300 280.400 14.400 ;
        RECT 268.400 13.700 280.400 14.300 ;
        RECT 268.400 13.600 269.200 13.700 ;
        RECT 279.600 13.600 280.400 13.700 ;
        RECT 308.400 14.300 309.200 14.400 ;
        RECT 324.400 14.300 325.200 14.400 ;
        RECT 330.800 14.300 331.600 14.400 ;
        RECT 308.400 13.700 331.600 14.300 ;
        RECT 308.400 13.600 309.200 13.700 ;
        RECT 324.400 13.600 325.200 13.700 ;
        RECT 330.800 13.600 331.600 13.700 ;
        RECT 68.400 12.300 69.200 12.400 ;
        RECT 79.600 12.300 80.400 12.400 ;
        RECT 68.400 11.700 80.400 12.300 ;
        RECT 68.400 11.600 69.200 11.700 ;
        RECT 79.600 11.600 80.400 11.700 ;
        RECT 116.400 12.300 117.200 12.400 ;
        RECT 225.200 12.300 226.000 12.400 ;
        RECT 116.400 11.700 226.000 12.300 ;
        RECT 116.400 11.600 117.200 11.700 ;
        RECT 225.200 11.600 226.000 11.700 ;
        RECT 242.800 12.300 243.600 12.400 ;
        RECT 255.600 12.300 256.400 12.400 ;
        RECT 242.800 11.700 256.400 12.300 ;
        RECT 242.800 11.600 243.600 11.700 ;
        RECT 255.600 11.600 256.400 11.700 ;
        RECT 265.200 12.300 266.000 12.400 ;
        RECT 271.600 12.300 272.400 12.400 ;
        RECT 290.800 12.300 291.600 12.400 ;
        RECT 265.200 11.700 291.600 12.300 ;
        RECT 265.200 11.600 266.000 11.700 ;
        RECT 271.600 11.600 272.400 11.700 ;
        RECT 290.800 11.600 291.600 11.700 ;
        RECT 329.200 12.300 330.000 12.400 ;
        RECT 358.000 12.300 358.800 12.400 ;
        RECT 329.200 11.700 358.800 12.300 ;
        RECT 329.200 11.600 330.000 11.700 ;
        RECT 358.000 11.600 358.800 11.700 ;
        RECT 396.400 12.300 397.200 12.400 ;
        RECT 399.600 12.300 400.400 12.400 ;
        RECT 396.400 11.700 400.400 12.300 ;
        RECT 396.400 11.600 397.200 11.700 ;
        RECT 399.600 11.600 400.400 11.700 ;
        RECT 458.800 12.300 459.600 12.400 ;
        RECT 462.000 12.300 462.800 12.400 ;
        RECT 458.800 11.700 462.800 12.300 ;
        RECT 458.800 11.600 459.600 11.700 ;
        RECT 462.000 11.600 462.800 11.700 ;
        RECT 545.200 11.600 546.000 12.400 ;
        RECT 166.000 10.300 166.800 10.400 ;
        RECT 185.200 10.300 186.000 10.400 ;
        RECT 166.000 9.700 186.000 10.300 ;
        RECT 166.000 9.600 166.800 9.700 ;
        RECT 185.200 9.600 186.000 9.700 ;
        RECT 222.000 10.300 222.800 10.400 ;
        RECT 230.000 10.300 230.800 10.400 ;
        RECT 249.200 10.300 250.000 10.400 ;
        RECT 254.000 10.300 254.800 10.400 ;
        RECT 274.800 10.300 275.600 10.400 ;
        RECT 222.000 9.700 275.600 10.300 ;
        RECT 222.000 9.600 222.800 9.700 ;
        RECT 230.000 9.600 230.800 9.700 ;
        RECT 249.200 9.600 250.000 9.700 ;
        RECT 254.000 9.600 254.800 9.700 ;
        RECT 274.800 9.600 275.600 9.700 ;
        RECT 278.000 10.300 278.800 10.400 ;
        RECT 287.600 10.300 288.400 10.400 ;
        RECT 278.000 9.700 288.400 10.300 ;
        RECT 278.000 9.600 278.800 9.700 ;
        RECT 287.600 9.600 288.400 9.700 ;
        RECT 332.400 10.300 333.200 10.400 ;
        RECT 338.800 10.300 339.600 10.400 ;
        RECT 332.400 9.700 339.600 10.300 ;
        RECT 332.400 9.600 333.200 9.700 ;
        RECT 338.800 9.600 339.600 9.700 ;
        RECT 225.200 8.300 226.000 8.400 ;
        RECT 228.400 8.300 229.200 8.400 ;
        RECT 225.200 7.700 229.200 8.300 ;
        RECT 225.200 7.600 226.000 7.700 ;
        RECT 228.400 7.600 229.200 7.700 ;
        RECT 236.400 8.300 237.200 8.400 ;
        RECT 239.600 8.300 240.400 8.400 ;
        RECT 236.400 7.700 240.400 8.300 ;
        RECT 236.400 7.600 237.200 7.700 ;
        RECT 239.600 7.600 240.400 7.700 ;
        RECT 254.000 8.300 254.800 8.400 ;
        RECT 310.000 8.300 310.800 8.400 ;
        RECT 254.000 7.700 310.800 8.300 ;
        RECT 254.000 7.600 254.800 7.700 ;
        RECT 310.000 7.600 310.800 7.700 ;
      LAYER metal4 ;
        RECT 26.600 321.400 27.800 374.600 ;
        RECT 13.800 251.400 15.000 296.600 ;
        RECT 23.400 257.400 24.600 278.600 ;
        RECT 29.800 267.400 31.000 272.600 ;
        RECT 33.000 255.400 34.200 306.600 ;
        RECT 20.200 225.400 21.400 246.600 ;
        RECT 4.200 111.400 5.400 152.600 ;
        RECT 20.200 121.400 21.400 146.600 ;
        RECT 23.400 139.400 24.600 206.600 ;
        RECT 29.800 185.400 31.000 246.600 ;
        RECT 33.000 193.400 34.200 226.600 ;
        RECT 39.400 211.400 40.600 286.600 ;
        RECT 45.800 265.400 47.000 304.600 ;
        RECT 26.600 125.400 27.800 182.600 ;
        RECT 42.600 167.400 43.800 208.600 ;
        RECT 45.800 193.400 47.000 256.600 ;
        RECT 52.200 249.400 53.400 300.600 ;
        RECT 55.400 265.400 56.600 316.600 ;
        RECT 61.800 227.400 63.000 250.600 ;
        RECT 68.200 249.400 69.400 304.600 ;
        RECT 71.400 265.400 72.600 364.600 ;
        RECT 74.600 295.400 75.800 344.600 ;
        RECT 74.600 265.400 75.800 284.600 ;
        RECT 29.800 121.400 31.000 166.600 ;
        RECT 49.000 159.400 50.200 198.600 ;
        RECT 29.800 81.400 31.000 94.600 ;
        RECT 39.400 91.400 40.600 148.600 ;
        RECT 42.600 97.400 43.800 154.600 ;
        RECT 45.800 53.400 47.000 120.600 ;
        RECT 52.200 93.400 53.400 184.600 ;
        RECT 68.200 115.400 69.400 208.600 ;
        RECT 81.000 153.400 82.200 340.600 ;
        RECT 93.800 173.400 95.000 200.600 ;
        RECT 58.600 71.400 59.800 108.600 ;
        RECT 87.400 91.400 88.600 168.600 ;
        RECT 100.200 139.400 101.400 200.600 ;
        RECT 109.800 197.400 111.000 286.600 ;
        RECT 132.200 267.400 133.400 300.600 ;
        RECT 132.200 187.400 133.400 228.600 ;
        RECT 135.400 217.400 136.600 270.600 ;
        RECT 141.800 264.600 143.000 270.600 ;
        RECT 140.200 263.400 143.000 264.600 ;
        RECT 100.200 91.400 101.400 118.600 ;
        RECT 116.200 69.400 117.400 146.600 ;
        RECT 145.000 135.400 146.200 262.600 ;
        RECT 154.600 241.400 155.800 268.600 ;
        RECT 157.800 253.400 159.000 278.600 ;
        RECT 167.400 231.400 168.600 260.600 ;
        RECT 173.800 259.400 175.000 276.600 ;
        RECT 177.000 231.400 178.200 306.600 ;
        RECT 180.200 299.400 181.400 330.600 ;
        RECT 237.800 321.400 239.000 344.600 ;
        RECT 285.800 323.400 287.000 346.600 ;
        RECT 324.200 337.400 325.400 364.600 ;
        RECT 164.200 127.400 165.400 224.600 ;
        RECT 20.200 13.400 21.400 38.600 ;
        RECT 55.400 27.400 56.600 60.600 ;
        RECT 145.000 55.400 146.200 102.600 ;
        RECT 148.200 49.400 149.400 106.600 ;
        RECT 183.400 97.400 184.600 236.600 ;
        RECT 189.800 127.400 191.000 290.600 ;
        RECT 205.800 237.400 207.000 284.600 ;
        RECT 193.000 93.400 194.200 130.600 ;
        RECT 196.200 113.400 197.400 148.600 ;
        RECT 212.200 105.400 213.400 182.600 ;
        RECT 215.400 151.400 216.600 276.600 ;
        RECT 225.000 205.400 226.200 280.600 ;
        RECT 225.000 103.400 226.200 194.600 ;
        RECT 228.200 175.400 229.400 194.600 ;
        RECT 231.400 127.400 232.600 206.600 ;
        RECT 234.600 205.400 235.800 290.600 ;
        RECT 241.000 257.400 242.200 292.600 ;
        RECT 247.400 175.400 248.600 274.600 ;
        RECT 282.600 249.400 283.800 280.600 ;
        RECT 289.000 255.400 290.200 268.600 ;
        RECT 241.000 135.400 242.200 158.600 ;
        RECT 250.600 139.400 251.800 204.600 ;
        RECT 260.200 201.400 261.400 228.600 ;
        RECT 282.600 173.400 283.800 192.600 ;
        RECT 295.400 125.400 296.600 276.600 ;
        RECT 301.800 173.400 303.000 266.600 ;
        RECT 161.000 51.400 162.200 88.600 ;
        RECT 228.200 73.400 229.400 98.600 ;
        RECT 247.400 53.400 248.600 112.600 ;
        RECT 308.200 13.400 309.400 170.600 ;
        RECT 333.800 165.400 335.000 298.600 ;
        RECT 337.000 291.400 338.200 332.600 ;
        RECT 359.400 327.400 360.600 374.600 ;
        RECT 365.800 303.400 367.000 368.600 ;
        RECT 372.200 329.400 373.400 350.600 ;
        RECT 346.600 247.400 347.800 298.600 ;
        RECT 375.400 289.400 376.600 322.600 ;
        RECT 391.400 321.400 392.600 372.600 ;
        RECT 397.800 327.400 399.000 358.600 ;
        RECT 442.600 353.400 443.800 358.600 ;
        RECT 410.600 343.400 411.800 350.600 ;
        RECT 385.000 291.400 386.200 296.600 ;
        RECT 401.000 289.400 402.200 334.600 ;
        RECT 404.200 307.400 405.400 328.600 ;
        RECT 407.400 289.400 408.600 330.600 ;
        RECT 436.200 329.400 437.400 334.600 ;
        RECT 449.000 331.400 450.200 350.600 ;
        RECT 337.000 215.400 338.200 220.600 ;
        RECT 349.800 177.400 351.000 210.600 ;
        RECT 353.000 193.400 354.200 274.600 ;
        RECT 359.400 177.400 360.600 240.600 ;
        RECT 375.400 209.400 376.600 218.600 ;
        RECT 381.800 207.400 383.000 258.600 ;
        RECT 407.400 215.400 408.600 272.600 ;
        RECT 372.200 113.400 373.400 158.600 ;
        RECT 375.400 145.400 376.600 190.600 ;
        RECT 353.000 55.400 354.200 82.600 ;
        RECT 362.600 51.400 363.800 106.600 ;
        RECT 369.000 53.400 370.200 102.600 ;
        RECT 385.000 87.400 386.200 136.600 ;
        RECT 394.600 121.400 395.800 200.600 ;
        RECT 397.800 157.400 399.000 212.600 ;
        RECT 401.000 147.400 402.200 174.600 ;
        RECT 410.600 129.400 411.800 216.600 ;
        RECT 445.800 215.400 447.000 260.600 ;
        RECT 455.400 213.400 456.600 258.600 ;
        RECT 458.600 227.400 459.800 338.600 ;
        RECT 413.800 201.400 415.000 208.600 ;
        RECT 417.000 149.400 418.200 180.600 ;
        RECT 436.200 109.400 437.400 194.600 ;
        RECT 385.000 27.400 386.200 60.600 ;
        RECT 407.400 53.400 408.600 94.600 ;
        RECT 433.000 21.400 434.200 56.600 ;
        RECT 442.600 51.400 443.800 84.600 ;
        RECT 445.800 81.400 447.000 108.600 ;
        RECT 455.400 107.400 456.600 206.600 ;
        RECT 458.600 203.400 459.800 222.600 ;
        RECT 465.000 211.400 466.200 346.600 ;
        RECT 468.200 261.400 469.400 340.600 ;
        RECT 474.600 317.400 475.800 336.600 ;
        RECT 461.800 145.400 463.000 202.600 ;
        RECT 465.000 159.400 466.200 190.600 ;
        RECT 468.200 89.400 469.400 180.600 ;
        RECT 471.400 173.400 472.600 228.600 ;
        RECT 474.600 141.400 475.800 228.600 ;
        RECT 477.800 179.400 479.000 294.600 ;
        RECT 481.000 189.400 482.200 258.600 ;
        RECT 500.200 217.400 501.400 292.600 ;
        RECT 477.800 109.400 479.000 174.600 ;
        RECT 481.000 139.400 482.200 180.600 ;
        RECT 468.200 41.400 469.400 62.600 ;
        RECT 471.400 23.400 472.600 74.600 ;
        RECT 487.400 31.400 488.600 212.600 ;
        RECT 497.000 165.400 498.200 176.600 ;
        RECT 500.200 131.400 501.400 200.600 ;
        RECT 503.400 149.400 504.600 304.600 ;
        RECT 497.000 75.400 498.200 100.600 ;
        RECT 503.400 71.400 504.600 112.600 ;
        RECT 497.000 23.400 498.200 44.600 ;
        RECT 500.200 23.400 501.400 70.600 ;
        RECT 503.400 21.400 504.600 46.600 ;
        RECT 506.600 45.400 507.800 126.600 ;
        RECT 509.800 69.400 511.000 252.600 ;
        RECT 522.600 221.400 523.800 344.600 ;
        RECT 525.800 279.400 527.000 368.600 ;
        RECT 519.400 37.400 520.600 154.600 ;
        RECT 522.600 31.400 523.800 204.600 ;
        RECT 525.800 171.400 527.000 226.600 ;
        RECT 532.200 191.400 533.400 300.600 ;
        RECT 535.400 211.400 536.600 296.600 ;
        RECT 538.600 187.400 539.800 344.600 ;
        RECT 532.200 37.400 533.400 140.600 ;
        RECT 541.800 33.400 543.000 258.600 ;
        RECT 545.000 11.400 546.200 180.600 ;
  END
END i2c_master_top
END LIBRARY

