magic
tech scmos
magscale 1 2
timestamp 1618241807
<< metal1 >>
rect 1866 1814 1878 1816
rect 1851 1806 1853 1814
rect 1861 1806 1863 1814
rect 1871 1806 1873 1814
rect 1881 1806 1883 1814
rect 1891 1806 1893 1814
rect 1866 1804 1878 1806
rect 429 1757 467 1763
rect 2436 1737 2467 1743
rect 45 1717 82 1723
rect 958 1717 995 1723
rect 1069 1717 1106 1723
rect 1854 1717 1948 1723
rect 2318 1717 2355 1723
rect 2429 1717 2444 1723
rect 2525 1677 2540 1683
rect 2420 1636 2422 1644
rect 666 1614 678 1616
rect 651 1606 653 1614
rect 661 1606 663 1614
rect 671 1606 673 1614
rect 681 1606 683 1614
rect 691 1606 693 1614
rect 666 1604 678 1606
rect 1844 1576 1846 1584
rect 45 1497 82 1503
rect 957 1483 963 1503
rect 788 1477 883 1483
rect 909 1477 947 1483
rect 957 1477 988 1483
rect 909 1457 915 1477
rect 1085 1483 1091 1503
rect 1124 1497 1139 1503
rect 1284 1497 1299 1503
rect 1869 1503 1875 1523
rect 1869 1497 1971 1503
rect 2141 1503 2147 1523
rect 2404 1516 2412 1524
rect 2141 1497 2179 1503
rect 2372 1497 2403 1503
rect 1076 1477 1091 1483
rect 1988 1477 2003 1483
rect 1092 1457 1107 1463
rect 1197 1457 1235 1463
rect 1997 1457 2003 1477
rect 2461 1477 2499 1483
rect 2013 1457 2028 1463
rect 2461 1457 2467 1477
rect 1396 1436 1398 1444
rect 2058 1436 2060 1444
rect 2244 1436 2248 1444
rect 1866 1414 1878 1416
rect 1851 1406 1853 1414
rect 1861 1406 1863 1414
rect 1871 1406 1873 1414
rect 1881 1406 1883 1414
rect 1891 1406 1893 1414
rect 1866 1404 1878 1406
rect 621 1357 684 1363
rect 429 1337 451 1343
rect 516 1337 531 1343
rect 605 1337 700 1343
rect 1565 1337 1596 1343
rect 2004 1337 2019 1343
rect 2253 1337 2268 1343
rect 45 1317 82 1323
rect 628 1317 723 1323
rect 1693 1317 1747 1323
rect 1780 1317 1795 1323
rect 1828 1317 1900 1323
rect 2020 1317 2035 1323
rect 2068 1317 2083 1323
rect 1821 1297 1868 1303
rect 2077 1297 2083 1317
rect 2276 1317 2291 1323
rect 2301 1317 2332 1323
rect 2301 1297 2307 1317
rect 2388 1317 2403 1323
rect 2036 1236 2038 1244
rect 666 1214 678 1216
rect 651 1206 653 1214
rect 661 1206 663 1214
rect 671 1206 673 1214
rect 681 1206 683 1214
rect 691 1206 693 1214
rect 666 1204 678 1206
rect 660 1137 723 1143
rect 1741 1137 1756 1143
rect 2492 1137 2540 1143
rect 804 1116 808 1124
rect 1364 1117 1379 1123
rect 45 1097 82 1103
rect 749 1097 771 1103
rect 765 1084 771 1097
rect 1469 1097 1484 1103
rect 1773 1097 1795 1103
rect 2436 1097 2467 1103
rect 461 1077 499 1083
rect 461 1057 467 1077
rect 1773 1077 1788 1083
rect 1844 1077 1923 1083
rect 1949 1077 2003 1083
rect 1946 1036 1948 1044
rect 1866 1014 1878 1016
rect 1851 1006 1853 1014
rect 1861 1006 1863 1014
rect 1871 1006 1873 1014
rect 1881 1006 1883 1014
rect 1891 1006 1893 1014
rect 1866 1004 1878 1006
rect 605 943 611 963
rect 804 957 835 963
rect 2148 956 2156 964
rect 596 937 611 943
rect 628 937 707 943
rect 765 937 787 943
rect 1565 937 1603 943
rect 45 917 82 923
rect 468 917 524 923
rect 1524 917 1539 923
rect 1597 917 1619 923
rect 1741 917 1779 923
rect 1508 897 1523 903
rect 1821 897 1907 903
rect 2356 897 2371 903
rect 2106 876 2108 884
rect 2180 877 2195 883
rect 1732 836 1734 844
rect 2036 836 2038 844
rect 666 814 678 816
rect 651 806 653 814
rect 661 806 663 814
rect 671 806 673 814
rect 681 806 683 814
rect 691 806 693 814
rect 666 804 678 806
rect 1773 777 1788 783
rect 509 697 524 703
rect 1188 697 1203 703
rect 1373 697 1452 703
rect 1556 697 1587 703
rect 1725 697 1740 703
rect 460 692 468 696
rect 1428 677 1443 683
rect 1636 677 1651 683
rect 1709 677 1724 683
rect 1421 663 1427 676
rect 1405 657 1427 663
rect 2500 657 2515 663
rect 2356 636 2360 644
rect 1866 614 1878 616
rect 1851 606 1853 614
rect 1861 606 1863 614
rect 1871 606 1873 614
rect 1881 606 1883 614
rect 1891 606 1893 614
rect 1866 604 1878 606
rect 2506 576 2508 584
rect 100 557 115 563
rect 1501 557 1516 563
rect 804 537 867 543
rect 1396 537 1411 543
rect 1469 537 1484 543
rect 1972 537 1992 543
rect 45 517 60 523
rect 1949 517 1964 523
rect 2414 517 2451 523
rect 1405 497 1443 503
rect 2029 497 2067 503
rect 666 414 678 416
rect 651 406 653 414
rect 661 406 663 414
rect 671 406 673 414
rect 681 406 683 414
rect 691 406 693 414
rect 666 404 678 406
rect 1965 317 1987 323
rect 45 297 82 303
rect 484 297 499 303
rect 509 283 515 303
rect 2013 297 2028 303
rect 509 277 531 283
rect 1028 277 1059 283
rect 2029 277 2051 283
rect 2493 277 2540 283
rect 957 257 995 263
rect 1005 257 1043 263
rect 1866 214 1878 216
rect 1851 206 1853 214
rect 1861 206 1863 214
rect 1871 206 1873 214
rect 1881 206 1883 214
rect 1891 206 1893 214
rect 1866 204 1878 206
rect 429 157 467 163
rect 1197 157 1212 163
rect 1908 157 1987 163
rect 493 137 524 143
rect 1133 137 1155 143
rect 2029 137 2067 143
rect 45 117 82 123
rect 1101 117 1116 123
rect 1997 117 2012 123
rect 2525 97 2540 103
rect 666 14 678 16
rect 651 6 653 14
rect 661 6 663 14
rect 671 6 673 14
rect 681 6 683 14
rect 691 6 693 14
rect 666 4 678 6
<< m2contact >>
rect 1843 1806 1851 1814
rect 1853 1806 1861 1814
rect 1863 1806 1871 1814
rect 1873 1806 1881 1814
rect 1883 1806 1891 1814
rect 1893 1806 1901 1814
rect 476 1776 484 1784
rect 524 1776 532 1784
rect 1020 1776 1028 1784
rect 1036 1776 1044 1784
rect 1468 1776 1476 1784
rect 1516 1776 1524 1784
rect 1980 1776 1988 1784
rect 2380 1776 2388 1784
rect 76 1756 84 1764
rect 236 1756 244 1764
rect 412 1756 420 1764
rect 796 1756 804 1764
rect 1260 1756 1268 1764
rect 1692 1756 1700 1764
rect 2156 1756 2164 1764
rect 2396 1756 2404 1764
rect 268 1736 276 1744
rect 492 1736 500 1744
rect 764 1736 772 1744
rect 1292 1736 1300 1744
rect 1660 1736 1668 1744
rect 2124 1736 2132 1744
rect 2428 1736 2436 1744
rect 2476 1736 2484 1744
rect 348 1716 356 1724
rect 444 1716 452 1724
rect 508 1716 516 1724
rect 556 1716 564 1724
rect 668 1716 676 1724
rect 1388 1716 1396 1724
rect 1436 1716 1444 1724
rect 1484 1716 1492 1724
rect 1660 1716 1668 1724
rect 1948 1716 1956 1724
rect 2028 1716 2036 1724
rect 2444 1716 2452 1724
rect 2492 1716 2500 1724
rect 364 1696 372 1704
rect 700 1700 708 1708
rect 1356 1700 1364 1708
rect 1596 1700 1604 1708
rect 2028 1696 2036 1704
rect 2444 1696 2452 1704
rect 12 1676 20 1684
rect 2540 1676 2548 1684
rect 700 1654 708 1662
rect 1596 1654 1604 1662
rect 364 1636 372 1644
rect 956 1636 964 1644
rect 1100 1636 1108 1644
rect 1356 1636 1364 1644
rect 2028 1636 2036 1644
rect 2316 1636 2324 1644
rect 2412 1636 2420 1644
rect 643 1606 651 1614
rect 653 1606 661 1614
rect 663 1606 671 1614
rect 673 1606 681 1614
rect 683 1606 691 1614
rect 693 1606 701 1614
rect 364 1576 372 1584
rect 476 1576 484 1584
rect 908 1576 916 1584
rect 1164 1576 1172 1584
rect 1228 1576 1236 1584
rect 1356 1576 1364 1584
rect 1772 1576 1780 1584
rect 1836 1576 1844 1584
rect 1484 1558 1492 1566
rect 2444 1536 2452 1544
rect 364 1516 372 1524
rect 476 1516 484 1524
rect 1404 1516 1412 1524
rect 1484 1512 1492 1520
rect 348 1496 356 1504
rect 476 1496 484 1504
rect 860 1496 868 1504
rect 12 1476 20 1484
rect 74 1476 82 1484
rect 268 1476 276 1484
rect 572 1476 580 1484
rect 780 1476 788 1484
rect 972 1496 980 1504
rect 1036 1496 1044 1504
rect 236 1456 244 1464
rect 412 1456 420 1464
rect 604 1456 612 1464
rect 988 1476 996 1484
rect 1068 1476 1076 1484
rect 1116 1496 1124 1504
rect 1212 1496 1220 1504
rect 1276 1496 1284 1504
rect 1324 1496 1332 1504
rect 1468 1496 1476 1504
rect 1660 1496 1668 1504
rect 1804 1496 1812 1504
rect 1836 1496 1844 1504
rect 1948 1516 1956 1524
rect 2044 1516 2052 1524
rect 2028 1496 2036 1504
rect 2108 1496 2116 1504
rect 2124 1496 2132 1504
rect 2156 1516 2164 1524
rect 2364 1516 2372 1524
rect 2396 1516 2404 1524
rect 2428 1516 2436 1524
rect 2332 1496 2340 1504
rect 2364 1496 2372 1504
rect 2508 1496 2516 1504
rect 1260 1476 1268 1484
rect 1372 1476 1380 1484
rect 1548 1476 1556 1484
rect 1820 1476 1828 1484
rect 1980 1476 1988 1484
rect 924 1456 932 1464
rect 1020 1456 1028 1464
rect 1084 1456 1092 1464
rect 1116 1456 1124 1464
rect 1180 1456 1188 1464
rect 1308 1456 1316 1464
rect 1580 1456 1588 1464
rect 2076 1476 2084 1484
rect 2092 1476 2100 1484
rect 2188 1476 2196 1484
rect 2204 1476 2212 1484
rect 2300 1476 2308 1484
rect 2316 1476 2324 1484
rect 2348 1476 2356 1484
rect 2380 1476 2388 1484
rect 2028 1456 2036 1464
rect 2476 1456 2484 1464
rect 428 1436 436 1444
rect 764 1436 772 1444
rect 1004 1436 1012 1444
rect 1388 1436 1396 1444
rect 1740 1436 1748 1444
rect 2060 1436 2068 1444
rect 2236 1436 2244 1444
rect 2492 1436 2500 1444
rect 1843 1406 1851 1414
rect 1853 1406 1861 1414
rect 1863 1406 1871 1414
rect 1873 1406 1881 1414
rect 1883 1406 1891 1414
rect 1893 1406 1901 1414
rect 748 1376 756 1384
rect 780 1376 788 1384
rect 1148 1376 1156 1384
rect 1196 1376 1204 1384
rect 1548 1376 1556 1384
rect 1612 1376 1620 1384
rect 1932 1376 1940 1384
rect 2076 1376 2084 1384
rect 2188 1376 2196 1384
rect 2364 1376 2372 1384
rect 76 1356 84 1364
rect 236 1356 244 1364
rect 412 1356 420 1364
rect 684 1356 692 1364
rect 988 1356 996 1364
rect 1356 1356 1364 1364
rect 1628 1356 1636 1364
rect 1660 1356 1668 1364
rect 1948 1356 1956 1364
rect 1964 1356 1972 1364
rect 2156 1356 2164 1364
rect 2172 1356 2180 1364
rect 2236 1356 2244 1364
rect 2380 1356 2388 1364
rect 2412 1356 2420 1364
rect 268 1336 276 1344
rect 476 1336 484 1344
rect 508 1336 516 1344
rect 556 1336 564 1344
rect 588 1336 596 1344
rect 700 1336 708 1344
rect 764 1336 772 1344
rect 956 1336 964 1344
rect 1388 1336 1396 1344
rect 1596 1336 1604 1344
rect 1644 1336 1652 1344
rect 1708 1336 1716 1344
rect 1756 1336 1764 1344
rect 1772 1336 1780 1344
rect 1804 1336 1812 1344
rect 1916 1336 1924 1344
rect 1996 1336 2004 1344
rect 2124 1336 2132 1344
rect 2204 1336 2212 1344
rect 2268 1336 2276 1344
rect 2316 1336 2324 1344
rect 348 1316 356 1324
rect 460 1316 468 1324
rect 492 1316 500 1324
rect 540 1316 548 1324
rect 572 1316 580 1324
rect 620 1316 628 1324
rect 748 1316 756 1324
rect 812 1316 820 1324
rect 1068 1316 1076 1324
rect 1468 1316 1476 1324
rect 1580 1316 1588 1324
rect 1660 1316 1668 1324
rect 1772 1316 1780 1324
rect 1820 1316 1828 1324
rect 1900 1316 1908 1324
rect 1996 1316 2004 1324
rect 2012 1316 2020 1324
rect 2060 1316 2068 1324
rect 364 1296 372 1304
rect 892 1300 900 1308
rect 1452 1300 1460 1308
rect 1868 1296 1876 1304
rect 2060 1296 2068 1304
rect 2108 1316 2116 1324
rect 2220 1316 2228 1324
rect 2268 1316 2276 1324
rect 2332 1316 2340 1324
rect 2380 1316 2388 1324
rect 2460 1316 2468 1324
rect 2364 1296 2372 1304
rect 2444 1296 2452 1304
rect 12 1276 20 1284
rect 1996 1276 2004 1284
rect 2476 1276 2484 1284
rect 892 1254 900 1262
rect 1452 1254 1460 1262
rect 364 1236 372 1244
rect 428 1236 436 1244
rect 780 1236 788 1244
rect 1740 1236 1748 1244
rect 2028 1236 2036 1244
rect 2140 1236 2148 1244
rect 2428 1236 2436 1244
rect 2492 1236 2500 1244
rect 643 1206 651 1214
rect 653 1206 661 1214
rect 663 1206 671 1214
rect 673 1206 681 1214
rect 683 1206 691 1214
rect 693 1206 701 1214
rect 364 1176 372 1184
rect 636 1176 644 1184
rect 988 1176 996 1184
rect 1276 1176 1284 1184
rect 1788 1176 1796 1184
rect 2156 1158 2164 1166
rect 652 1136 660 1144
rect 1756 1136 1764 1144
rect 2540 1136 2548 1144
rect 364 1116 372 1124
rect 572 1116 580 1124
rect 796 1116 804 1124
rect 988 1116 996 1124
rect 1356 1116 1364 1124
rect 1484 1116 1492 1124
rect 1644 1116 1652 1124
rect 2028 1116 2036 1124
rect 2156 1112 2164 1120
rect 348 1096 356 1104
rect 364 1096 372 1104
rect 412 1096 420 1104
rect 508 1096 516 1104
rect 540 1096 548 1104
rect 556 1096 564 1104
rect 604 1096 612 1104
rect 892 1096 900 1104
rect 924 1096 932 1104
rect 1084 1096 1092 1104
rect 1196 1096 1204 1104
rect 1308 1096 1316 1104
rect 1340 1096 1348 1104
rect 1388 1096 1396 1104
rect 1404 1096 1412 1104
rect 1452 1096 1460 1104
rect 1484 1096 1492 1104
rect 1516 1096 1524 1104
rect 1548 1096 1556 1104
rect 1628 1096 1636 1104
rect 1660 1096 1668 1104
rect 1676 1096 1684 1104
rect 1740 1096 1748 1104
rect 1900 1096 1908 1104
rect 1964 1096 1972 1104
rect 2012 1096 2020 1104
rect 2060 1096 2068 1104
rect 2124 1096 2132 1104
rect 2428 1096 2436 1104
rect 2476 1096 2484 1104
rect 12 1076 20 1084
rect 268 1076 276 1084
rect 428 1076 436 1084
rect 76 1056 84 1064
rect 236 1056 244 1064
rect 524 1076 532 1084
rect 588 1076 596 1084
rect 764 1076 772 1084
rect 860 1076 868 1084
rect 876 1076 884 1084
rect 908 1076 916 1084
rect 940 1076 948 1084
rect 1084 1076 1092 1084
rect 1356 1076 1364 1084
rect 1420 1076 1428 1084
rect 1436 1076 1444 1084
rect 1500 1076 1508 1084
rect 1532 1076 1540 1084
rect 1564 1076 1572 1084
rect 1612 1076 1620 1084
rect 1692 1076 1700 1084
rect 1788 1076 1796 1084
rect 1836 1076 1844 1084
rect 2044 1076 2052 1084
rect 2076 1076 2084 1084
rect 2220 1076 2228 1084
rect 2444 1076 2452 1084
rect 476 1056 484 1064
rect 1116 1056 1124 1064
rect 1580 1056 1588 1064
rect 1708 1056 1716 1064
rect 1756 1056 1764 1064
rect 1820 1056 1828 1064
rect 1980 1056 1988 1064
rect 2252 1056 2260 1064
rect 444 1036 452 1044
rect 1596 1036 1604 1044
rect 1948 1036 1956 1044
rect 2412 1036 2420 1044
rect 1843 1006 1851 1014
rect 1853 1006 1861 1014
rect 1863 1006 1871 1014
rect 1873 1006 1881 1014
rect 1883 1006 1891 1014
rect 1893 1006 1901 1014
rect 540 976 548 984
rect 780 976 788 984
rect 1484 976 1492 984
rect 1628 976 1636 984
rect 1820 976 1828 984
rect 1964 976 1972 984
rect 2268 976 2276 984
rect 2476 976 2484 984
rect 236 956 244 964
rect 428 956 436 964
rect 268 936 276 944
rect 412 936 420 944
rect 476 936 484 944
rect 492 936 500 944
rect 588 936 596 944
rect 796 956 804 964
rect 988 956 996 964
rect 1324 956 1332 964
rect 1580 956 1588 964
rect 1644 956 1652 964
rect 1660 956 1668 964
rect 1708 956 1716 964
rect 1804 956 1812 964
rect 2140 956 2148 964
rect 2220 956 2228 964
rect 2284 956 2292 964
rect 2380 956 2388 964
rect 2460 956 2468 964
rect 620 936 628 944
rect 732 936 740 944
rect 1020 936 1028 944
rect 1292 936 1300 944
rect 1788 936 1796 944
rect 1996 936 2004 944
rect 2012 936 2020 944
rect 2124 936 2132 944
rect 2172 936 2180 944
rect 2252 936 2260 944
rect 2348 936 2356 944
rect 2412 936 2420 944
rect 2444 936 2452 944
rect 2492 936 2500 944
rect 364 916 372 924
rect 428 916 436 924
rect 460 916 468 924
rect 524 916 532 924
rect 716 916 724 924
rect 748 916 756 924
rect 908 916 916 924
rect 1132 916 1140 924
rect 1196 916 1204 924
rect 1516 916 1524 924
rect 1548 916 1556 924
rect 1692 916 1700 924
rect 1916 916 1924 924
rect 2028 916 2036 924
rect 2108 916 2116 924
rect 2188 916 2196 924
rect 2236 916 2244 924
rect 2300 916 2308 924
rect 2332 916 2340 924
rect 2428 916 2436 924
rect 2508 916 2516 924
rect 76 896 84 904
rect 364 896 372 904
rect 1116 896 1124 904
rect 1228 900 1236 908
rect 1500 896 1508 904
rect 1756 896 1764 904
rect 1964 896 1972 904
rect 2060 896 2068 904
rect 2076 896 2084 904
rect 2140 896 2148 904
rect 2348 896 2356 904
rect 2396 896 2404 904
rect 12 876 20 884
rect 1692 876 1700 884
rect 1932 876 1940 884
rect 2108 876 2116 884
rect 2172 876 2180 884
rect 364 836 372 844
rect 780 836 788 844
rect 1116 836 1124 844
rect 1228 836 1236 844
rect 1484 836 1492 844
rect 1612 836 1620 844
rect 1724 836 1732 844
rect 1916 836 1924 844
rect 2028 836 2036 844
rect 643 806 651 814
rect 653 806 661 814
rect 663 806 671 814
rect 673 806 681 814
rect 683 806 691 814
rect 693 806 701 814
rect 172 776 180 784
rect 764 776 772 784
rect 796 776 804 784
rect 876 776 884 784
rect 1164 776 1172 784
rect 1292 776 1300 784
rect 1788 776 1796 784
rect 2172 776 2180 784
rect 1916 758 1924 766
rect 2444 756 2452 764
rect 12 736 20 744
rect 364 736 372 744
rect 2460 736 2468 744
rect 876 716 884 724
rect 1484 716 1492 724
rect 1548 716 1556 724
rect 1612 716 1620 724
rect 1628 716 1636 724
rect 1916 712 1924 720
rect 2428 716 2436 724
rect 44 696 52 704
rect 396 696 404 704
rect 428 696 436 704
rect 460 696 468 704
rect 476 696 484 704
rect 524 696 532 704
rect 828 696 836 704
rect 908 696 916 704
rect 1084 696 1092 704
rect 1180 696 1188 704
rect 1228 696 1236 704
rect 1260 696 1268 704
rect 1452 696 1460 704
rect 1516 696 1524 704
rect 1548 696 1556 704
rect 1740 696 1748 704
rect 1772 696 1780 704
rect 1884 696 1892 704
rect 2092 696 2100 704
rect 2204 696 2212 704
rect 2268 696 2276 704
rect 2284 696 2292 704
rect 2444 696 2452 704
rect 2492 696 2500 704
rect 60 676 68 684
rect 204 676 212 684
rect 380 676 388 684
rect 444 676 452 684
rect 524 676 532 684
rect 556 676 564 684
rect 572 676 580 684
rect 652 676 660 684
rect 972 676 980 684
rect 1244 676 1252 684
rect 1356 676 1364 684
rect 1388 676 1396 684
rect 1420 676 1428 684
rect 1500 676 1508 684
rect 1564 676 1572 684
rect 1628 676 1636 684
rect 1660 676 1668 684
rect 1724 676 1732 684
rect 1980 676 1988 684
rect 2220 676 2228 684
rect 2252 676 2260 684
rect 2316 676 2324 684
rect 2412 676 2420 684
rect 348 656 356 664
rect 1004 656 1012 664
rect 1612 656 1620 664
rect 1676 656 1684 664
rect 1692 656 1700 664
rect 1740 656 1748 664
rect 2012 656 2020 664
rect 2300 656 2308 664
rect 2492 656 2500 664
rect 2524 656 2532 664
rect 316 636 324 644
rect 428 636 436 644
rect 476 636 484 644
rect 1484 636 1492 644
rect 1548 636 1556 644
rect 2172 636 2180 644
rect 2236 636 2244 644
rect 2348 636 2356 644
rect 1843 606 1851 614
rect 1853 606 1861 614
rect 1863 606 1871 614
rect 1873 606 1881 614
rect 1883 606 1891 614
rect 1893 606 1901 614
rect 76 576 84 584
rect 460 576 468 584
rect 908 576 916 584
rect 1436 576 1444 584
rect 1532 576 1540 584
rect 2412 576 2420 584
rect 2508 576 2516 584
rect 60 556 68 564
rect 92 556 100 564
rect 268 556 276 564
rect 620 556 628 564
rect 1036 556 1044 564
rect 1212 556 1220 564
rect 1372 556 1380 564
rect 1420 556 1428 564
rect 1484 556 1492 564
rect 1516 556 1524 564
rect 1692 556 1700 564
rect 2252 556 2260 564
rect 300 536 308 544
rect 652 536 660 544
rect 796 536 804 544
rect 1020 536 1028 544
rect 1180 536 1188 544
rect 1388 536 1396 544
rect 1484 536 1492 544
rect 1724 536 1732 544
rect 1932 536 1940 544
rect 1964 536 1972 544
rect 2044 536 2052 544
rect 2220 536 2228 544
rect 2524 536 2532 544
rect 60 516 68 524
rect 380 516 388 524
rect 396 516 404 524
rect 540 516 548 524
rect 748 516 756 524
rect 892 516 900 524
rect 940 516 948 524
rect 956 516 964 524
rect 1004 516 1012 524
rect 1084 516 1092 524
rect 1724 516 1732 524
rect 1964 516 1972 524
rect 2012 516 2020 524
rect 2140 516 2148 524
rect 396 496 404 504
rect 748 496 756 504
rect 1116 500 1124 508
rect 1788 500 1796 508
rect 1964 496 1972 504
rect 2076 496 2084 504
rect 2156 500 2164 508
rect 2492 496 2500 504
rect 12 476 20 484
rect 1996 476 2004 484
rect 2476 476 2484 484
rect 1116 454 1124 462
rect 1788 454 1796 462
rect 2156 454 2164 462
rect 396 436 404 444
rect 748 436 756 444
rect 988 436 996 444
rect 643 406 651 414
rect 653 406 661 414
rect 663 406 671 414
rect 673 406 681 414
rect 683 406 691 414
rect 693 406 701 414
rect 364 376 372 384
rect 1212 376 1220 384
rect 1516 376 1524 384
rect 2396 376 2404 384
rect 2428 376 2436 384
rect 700 358 708 366
rect 2204 356 2212 364
rect 364 316 372 324
rect 700 312 708 320
rect 1244 316 1252 324
rect 1516 316 1524 324
rect 2108 316 2116 324
rect 2140 312 2148 320
rect 364 296 372 304
rect 460 296 468 304
rect 476 296 484 304
rect 12 276 20 284
rect 268 276 276 284
rect 428 276 436 284
rect 444 276 452 284
rect 556 296 564 304
rect 652 296 660 304
rect 764 296 772 304
rect 1020 296 1028 304
rect 1084 296 1092 304
rect 1436 296 1444 304
rect 1516 296 1524 304
rect 1724 296 1732 304
rect 1932 296 1940 304
rect 2028 296 2036 304
rect 2204 296 2212 304
rect 2460 296 2468 304
rect 764 276 772 284
rect 1020 276 1028 284
rect 1068 276 1076 284
rect 1100 276 1108 284
rect 1276 276 1284 284
rect 1292 276 1300 284
rect 1468 276 1476 284
rect 1612 276 1620 284
rect 1806 276 1814 284
rect 2204 276 2212 284
rect 2540 276 2548 284
rect 76 256 84 264
rect 236 256 244 264
rect 412 256 420 264
rect 476 256 484 264
rect 796 256 804 264
rect 1644 256 1652 264
rect 1948 256 1956 264
rect 2060 256 2068 264
rect 2236 256 2244 264
rect 2444 256 2452 264
rect 524 236 532 244
rect 956 236 964 244
rect 1244 236 1252 244
rect 1404 236 1412 244
rect 1900 236 1908 244
rect 1980 236 1988 244
rect 1843 206 1851 214
rect 1853 206 1861 214
rect 1863 206 1871 214
rect 1873 206 1881 214
rect 1883 206 1891 214
rect 1893 206 1901 214
rect 1004 176 1012 184
rect 2028 176 2036 184
rect 2108 176 2116 184
rect 2524 176 2532 184
rect 236 156 244 164
rect 412 156 420 164
rect 476 156 484 164
rect 748 156 756 164
rect 1116 156 1124 164
rect 1212 156 1220 164
rect 1388 156 1396 164
rect 1724 156 1732 164
rect 1884 156 1892 164
rect 1900 156 1908 164
rect 2012 156 2020 164
rect 2284 156 2292 164
rect 74 136 82 144
rect 268 136 276 144
rect 524 136 532 144
rect 716 136 724 144
rect 910 136 918 144
rect 1052 136 1060 144
rect 1420 136 1428 144
rect 1692 136 1700 144
rect 2252 136 2260 144
rect 2476 136 2484 144
rect 364 116 372 124
rect 444 116 452 124
rect 508 116 516 124
rect 636 116 644 124
rect 940 116 948 124
rect 1116 116 1124 124
rect 1164 116 1172 124
rect 1226 116 1234 124
rect 1516 116 1524 124
rect 1596 116 1604 124
rect 2012 116 2020 124
rect 2044 116 2052 124
rect 2076 116 2084 124
rect 2156 116 2164 124
rect 2492 116 2500 124
rect 332 100 340 108
rect 652 100 660 108
rect 1196 96 1204 104
rect 1484 100 1492 108
rect 1628 100 1636 108
rect 2188 100 2196 108
rect 2444 96 2452 104
rect 2540 96 2548 104
rect 12 76 20 84
rect 652 54 660 62
rect 332 36 340 44
rect 972 36 980 44
rect 1068 36 1076 44
rect 1484 36 1492 44
rect 1628 36 1636 44
rect 2188 36 2196 44
rect 643 6 651 14
rect 653 6 661 14
rect 663 6 671 14
rect 673 6 681 14
rect 683 6 691 14
rect 693 6 701 14
<< metal2 >>
rect 525 1857 547 1863
rect 1005 1857 1027 1863
rect 525 1784 531 1857
rect 1021 1784 1027 1857
rect 1037 1857 1059 1863
rect 1149 1857 1171 1863
rect 1037 1784 1043 1857
rect 13 1684 19 1696
rect 13 1484 19 1496
rect 237 1464 243 1756
rect 269 1744 275 1776
rect 445 1724 451 1736
rect 349 1504 355 1716
rect 365 1644 371 1696
rect 365 1524 371 1576
rect 237 1364 243 1456
rect 269 1424 275 1476
rect 13 1284 19 1296
rect 13 1084 19 1096
rect 237 1064 243 1356
rect 349 1324 355 1496
rect 413 1464 419 1476
rect 429 1364 435 1436
rect 349 1104 355 1316
rect 365 1244 371 1296
rect 445 1244 451 1716
rect 477 1524 483 1576
rect 509 1504 515 1716
rect 557 1584 563 1716
rect 701 1662 707 1700
rect 666 1614 678 1616
rect 651 1606 653 1614
rect 661 1606 663 1614
rect 671 1606 673 1614
rect 681 1606 683 1614
rect 691 1606 693 1614
rect 666 1604 678 1606
rect 509 1364 515 1436
rect 573 1424 579 1476
rect 509 1344 515 1356
rect 557 1344 563 1416
rect 685 1384 691 1576
rect 685 1364 691 1376
rect 701 1344 707 1496
rect 749 1384 755 1416
rect 765 1384 771 1436
rect 781 1384 787 1476
rect 797 1344 803 1756
rect 909 1584 915 1736
rect 557 1317 572 1323
rect 365 1124 371 1176
rect 429 1104 435 1236
rect 237 964 243 1056
rect 269 1044 275 1076
rect 13 884 19 896
rect 237 824 243 956
rect 365 924 371 1096
rect 413 944 419 1096
rect 429 944 435 956
rect 365 844 371 896
rect 173 784 179 816
rect 413 744 419 936
rect 13 724 19 736
rect 45 624 51 696
rect 77 584 83 716
rect 381 684 387 716
rect 429 704 435 916
rect 429 684 435 696
rect 445 684 451 956
rect 461 924 467 1316
rect 493 1304 499 1316
rect 509 1104 515 1236
rect 509 1084 515 1096
rect 525 1084 531 1116
rect 557 1104 563 1317
rect 589 1184 595 1336
rect 749 1304 755 1316
rect 541 1084 547 1096
rect 541 984 547 1076
rect 573 1064 579 1116
rect 605 1104 611 1116
rect 461 704 467 716
rect 477 684 483 696
rect 317 604 323 636
rect 349 624 355 656
rect 269 564 275 596
rect 61 524 67 556
rect 13 484 19 496
rect 269 304 275 556
rect 301 544 307 556
rect 381 544 387 676
rect 429 564 435 636
rect 365 324 371 376
rect 381 303 387 516
rect 397 444 403 496
rect 445 324 451 676
rect 461 584 467 616
rect 477 544 483 636
rect 493 624 499 936
rect 525 864 531 916
rect 589 904 595 936
rect 509 683 515 736
rect 525 704 531 856
rect 605 744 611 1056
rect 621 944 627 1276
rect 666 1214 678 1216
rect 651 1206 653 1214
rect 661 1206 663 1214
rect 671 1206 673 1214
rect 681 1206 683 1214
rect 691 1206 693 1214
rect 666 1204 678 1206
rect 749 1104 755 1296
rect 765 1224 771 1336
rect 845 1163 851 1376
rect 861 1284 867 1496
rect 957 1484 963 1636
rect 1165 1584 1171 1857
rect 1341 1824 1347 1863
rect 1453 1857 1475 1863
rect 1501 1857 1523 1863
rect 1469 1784 1475 1857
rect 1517 1784 1523 1857
rect 1773 1857 1795 1863
rect 1965 1857 1987 1863
rect 2365 1857 2387 1863
rect 925 1464 931 1476
rect 973 1444 979 1496
rect 1117 1464 1123 1496
rect 1181 1464 1187 1636
rect 1293 1624 1299 1736
rect 1357 1644 1363 1700
rect 1229 1584 1235 1616
rect 1005 1404 1011 1436
rect 957 1344 963 1396
rect 1117 1384 1123 1456
rect 1197 1384 1203 1496
rect 1213 1484 1219 1496
rect 989 1304 995 1356
rect 893 1262 899 1300
rect 1069 1263 1075 1316
rect 1117 1304 1123 1356
rect 1069 1257 1091 1263
rect 845 1157 867 1163
rect 717 924 723 1096
rect 861 1084 867 1157
rect 749 924 755 1016
rect 765 1004 771 1076
rect 877 1044 883 1076
rect 781 984 787 1036
rect 925 1024 931 1096
rect 941 1084 947 1216
rect 989 1124 995 1176
rect 1085 1104 1091 1257
rect 1117 1064 1123 1296
rect 1277 1224 1283 1496
rect 1309 1464 1315 1636
rect 1357 1584 1363 1616
rect 1389 1564 1395 1716
rect 1437 1644 1443 1716
rect 1485 1704 1491 1716
rect 1373 1484 1379 1496
rect 1309 1404 1315 1456
rect 1389 1364 1395 1436
rect 1405 1404 1411 1516
rect 1469 1504 1475 1556
rect 1485 1520 1491 1558
rect 1357 1124 1363 1336
rect 1389 1104 1395 1336
rect 1469 1324 1475 1496
rect 1549 1424 1555 1476
rect 1581 1464 1587 1756
rect 1597 1662 1603 1700
rect 1661 1504 1667 1716
rect 1773 1584 1779 1857
rect 1866 1814 1878 1816
rect 1851 1806 1853 1814
rect 1861 1806 1863 1814
rect 1871 1806 1873 1814
rect 1881 1806 1883 1814
rect 1891 1806 1893 1814
rect 1866 1804 1878 1806
rect 1981 1784 1987 1857
rect 2381 1784 2387 1857
rect 1837 1584 1843 1736
rect 1949 1604 1955 1716
rect 2029 1644 2035 1696
rect 1741 1444 1747 1496
rect 1549 1384 1555 1396
rect 1613 1384 1619 1416
rect 1581 1324 1587 1376
rect 1709 1344 1715 1436
rect 1757 1344 1763 1456
rect 1805 1344 1811 1476
rect 1821 1464 1827 1476
rect 1866 1414 1878 1416
rect 1851 1406 1853 1414
rect 1861 1406 1863 1414
rect 1871 1406 1873 1414
rect 1881 1406 1883 1414
rect 1891 1406 1893 1414
rect 1866 1404 1878 1406
rect 1453 1262 1459 1300
rect 666 814 678 816
rect 651 806 653 814
rect 661 806 663 814
rect 671 806 673 814
rect 681 806 683 814
rect 691 806 693 814
rect 666 804 678 806
rect 573 684 579 736
rect 717 684 723 916
rect 749 864 755 916
rect 765 784 771 976
rect 797 964 803 996
rect 1117 984 1123 1056
rect 989 964 995 976
rect 509 677 524 683
rect 653 664 659 676
rect 621 564 627 596
rect 653 564 659 656
rect 461 304 467 536
rect 372 297 387 303
rect 13 284 19 296
rect 237 264 243 296
rect 237 164 243 256
rect 269 144 275 156
rect 365 124 371 296
rect 413 264 419 296
rect 413 144 419 156
rect 445 124 451 276
rect 509 124 515 316
rect 621 264 627 556
rect 749 444 755 496
rect 666 414 678 416
rect 651 406 653 414
rect 661 406 663 414
rect 671 406 673 414
rect 681 406 683 414
rect 691 406 693 414
rect 666 404 678 406
rect 701 320 707 358
rect 765 304 771 516
rect 781 384 787 836
rect 797 784 803 916
rect 877 724 883 776
rect 909 704 915 916
rect 989 843 995 956
rect 1117 844 1123 896
rect 989 837 1011 843
rect 797 524 803 536
rect 829 524 835 696
rect 909 584 915 696
rect 973 684 979 756
rect 1005 664 1011 837
rect 1165 784 1171 996
rect 1197 924 1203 1096
rect 1309 1064 1315 1096
rect 1341 1084 1347 1096
rect 1357 1084 1363 1096
rect 1293 944 1299 1036
rect 1405 1024 1411 1096
rect 1421 1063 1427 1076
rect 1421 1057 1443 1063
rect 1325 964 1331 976
rect 1229 844 1235 900
rect 1293 784 1299 916
rect 1165 724 1171 776
rect 1229 704 1235 716
rect 1037 544 1043 556
rect 957 524 963 536
rect 1085 524 1091 696
rect 525 144 531 236
rect 653 143 659 296
rect 797 204 803 256
rect 749 164 755 196
rect 941 184 947 516
rect 957 304 963 516
rect 989 304 995 436
rect 1085 304 1091 376
rect 1069 284 1075 296
rect 1101 284 1107 556
rect 1181 544 1187 696
rect 1245 684 1251 776
rect 1389 684 1395 716
rect 1421 684 1427 836
rect 1213 564 1219 656
rect 1389 604 1395 676
rect 1437 584 1443 1057
rect 1453 824 1459 1096
rect 1469 924 1475 1316
rect 1549 1104 1555 1196
rect 1485 984 1491 1076
rect 1501 1064 1507 1076
rect 1533 1064 1539 1076
rect 1549 1024 1555 1096
rect 1597 1083 1603 1336
rect 1645 1283 1651 1336
rect 1661 1304 1667 1316
rect 1645 1277 1667 1283
rect 1629 1104 1635 1136
rect 1613 1084 1619 1096
rect 1597 1077 1612 1083
rect 1645 1083 1651 1116
rect 1661 1104 1667 1277
rect 1629 1077 1651 1083
rect 1581 964 1587 996
rect 1501 904 1507 936
rect 1453 704 1459 816
rect 1517 764 1523 916
rect 1549 864 1555 916
rect 1597 884 1603 1016
rect 1613 964 1619 1076
rect 1629 984 1635 1077
rect 1661 964 1667 1076
rect 1677 984 1683 1096
rect 1709 1083 1715 1336
rect 1741 1204 1747 1236
rect 1757 1144 1763 1336
rect 1821 1324 1827 1396
rect 1933 1384 1939 1496
rect 1949 1484 1955 1516
rect 1981 1484 1987 1596
rect 1773 1104 1779 1316
rect 1869 1304 1875 1376
rect 1949 1364 1955 1396
rect 1917 1344 1923 1356
rect 1901 1324 1907 1336
rect 1965 1324 1971 1356
rect 1997 1344 2003 1456
rect 2029 1364 2035 1456
rect 2029 1324 2035 1356
rect 2045 1344 2051 1516
rect 2125 1504 2131 1736
rect 2077 1484 2083 1496
rect 2061 1384 2067 1436
rect 2077 1384 2083 1456
rect 2061 1324 2067 1376
rect 1789 1184 1795 1296
rect 1901 1104 1907 1316
rect 2013 1303 2019 1316
rect 1997 1297 2019 1303
rect 1997 1284 2003 1297
rect 2029 1264 2035 1316
rect 1700 1077 1715 1083
rect 1693 964 1699 1076
rect 1709 1004 1715 1056
rect 1757 984 1763 1056
rect 1773 1044 1779 1096
rect 1901 1064 1907 1096
rect 1821 984 1827 1056
rect 1949 1024 1955 1036
rect 1866 1014 1878 1016
rect 1851 1006 1853 1014
rect 1861 1006 1863 1014
rect 1871 1006 1873 1014
rect 1881 1006 1883 1014
rect 1891 1006 1893 1014
rect 1866 1004 1878 1006
rect 1709 964 1715 976
rect 1693 924 1699 956
rect 1981 944 1987 1056
rect 1997 944 2003 1256
rect 2029 1124 2035 1236
rect 2013 1104 2019 1116
rect 2061 1024 2067 1096
rect 2093 1083 2099 1476
rect 2109 1464 2115 1496
rect 2157 1484 2163 1516
rect 2317 1504 2323 1636
rect 2333 1504 2339 1536
rect 2189 1484 2195 1496
rect 2365 1484 2371 1496
rect 2189 1384 2195 1396
rect 2109 1324 2115 1376
rect 2205 1364 2211 1476
rect 2301 1464 2307 1476
rect 2237 1364 2243 1376
rect 2173 1344 2179 1356
rect 2269 1344 2275 1356
rect 2317 1344 2323 1356
rect 2141 1124 2147 1236
rect 2157 1120 2163 1158
rect 2349 1144 2355 1476
rect 2365 1384 2371 1476
rect 2381 1464 2387 1476
rect 2381 1364 2387 1436
rect 2413 1384 2419 1636
rect 2429 1564 2435 1736
rect 2452 1717 2467 1723
rect 2445 1564 2451 1696
rect 2461 1524 2467 1717
rect 2493 1684 2499 1716
rect 2541 1684 2547 1696
rect 2429 1504 2435 1516
rect 2509 1504 2515 1596
rect 2365 1304 2371 1356
rect 2445 1304 2451 1356
rect 2461 1324 2467 1376
rect 2084 1077 2099 1083
rect 2013 944 2019 976
rect 1693 884 1699 896
rect 1549 784 1555 856
rect 1549 744 1555 756
rect 1597 743 1603 876
rect 1725 844 1731 856
rect 1613 764 1619 836
rect 1597 737 1619 743
rect 1549 724 1555 736
rect 1613 724 1619 737
rect 1485 564 1491 636
rect 1517 564 1523 696
rect 1549 684 1555 696
rect 1725 684 1731 836
rect 1741 724 1747 936
rect 1789 784 1795 936
rect 1997 924 2003 936
rect 1741 704 1747 716
rect 1885 704 1891 916
rect 1933 884 1939 896
rect 1917 824 1923 836
rect 1917 720 1923 758
rect 1773 684 1779 696
rect 1981 684 1987 776
rect 2013 764 2019 936
rect 2029 924 2035 1016
rect 2077 984 2083 1076
rect 2125 1064 2131 1096
rect 2061 904 2067 956
rect 2077 884 2083 896
rect 2029 784 2035 836
rect 2013 664 2019 716
rect 2093 704 2099 1056
rect 2109 924 2115 976
rect 2125 944 2131 1036
rect 2381 1024 2387 1296
rect 2493 1283 2499 1436
rect 2484 1277 2499 1283
rect 2429 1104 2435 1236
rect 2269 984 2275 1016
rect 2173 944 2179 956
rect 2189 904 2195 916
rect 2141 884 2147 896
rect 2173 884 2179 896
rect 2221 784 2227 956
rect 2253 944 2259 976
rect 2285 964 2291 976
rect 2381 964 2387 1016
rect 2237 924 2243 936
rect 2301 924 2307 936
rect 2349 924 2355 936
rect 2333 903 2339 916
rect 2381 904 2387 956
rect 2397 904 2403 1036
rect 2413 1024 2419 1036
rect 2413 944 2419 956
rect 2429 944 2435 1096
rect 2445 1084 2451 1276
rect 2445 944 2451 1076
rect 2493 963 2499 1236
rect 2541 1144 2547 1516
rect 2477 957 2499 963
rect 2429 924 2435 936
rect 2445 924 2451 936
rect 2333 897 2348 903
rect 2221 684 2227 756
rect 2397 744 2403 896
rect 2429 724 2435 736
rect 2445 724 2451 756
rect 2477 723 2483 957
rect 2477 717 2499 723
rect 2269 704 2275 716
rect 2317 684 2323 696
rect 2253 664 2259 676
rect 2301 664 2307 676
rect 2413 664 2419 676
rect 1741 644 1747 656
rect 1533 584 1539 596
rect 1117 462 1123 500
rect 1213 384 1219 556
rect 1245 304 1251 316
rect 637 137 659 143
rect 525 124 531 136
rect 637 124 643 137
rect 13 84 19 96
rect 333 44 339 100
rect 653 62 659 100
rect 666 14 678 16
rect 651 6 653 14
rect 661 6 663 14
rect 671 6 673 14
rect 681 6 683 14
rect 691 6 693 14
rect 666 4 678 6
rect 717 -17 723 136
rect 957 123 963 236
rect 1005 184 1011 236
rect 948 117 963 123
rect 973 -17 979 36
rect 1053 24 1059 136
rect 1117 124 1123 156
rect 1165 124 1171 296
rect 1245 104 1251 236
rect 717 -23 755 -17
rect 957 -23 979 -17
rect 1069 -23 1075 36
rect 1101 -23 1107 16
rect 1277 -17 1283 276
rect 1405 244 1411 256
rect 1437 244 1443 296
rect 1469 284 1475 296
rect 1485 284 1491 536
rect 1549 484 1555 636
rect 1741 604 1747 636
rect 1866 614 1878 616
rect 1851 606 1853 614
rect 1861 606 1863 614
rect 1871 606 1873 614
rect 1881 606 1883 614
rect 1891 606 1893 614
rect 1866 604 1878 606
rect 1517 324 1523 376
rect 1405 203 1411 236
rect 1389 197 1411 203
rect 1389 164 1395 197
rect 1421 144 1427 156
rect 1517 124 1523 296
rect 1613 284 1619 556
rect 1693 424 1699 556
rect 1917 543 1923 636
rect 2237 603 2243 636
rect 2301 624 2307 656
rect 2221 597 2243 603
rect 2045 544 2051 596
rect 2221 544 2227 597
rect 1917 537 1932 543
rect 1645 264 1651 416
rect 1725 324 1731 516
rect 1789 462 1795 500
rect 1725 304 1731 316
rect 1933 304 1939 536
rect 2141 320 2147 516
rect 2157 462 2163 500
rect 2253 443 2259 556
rect 2349 504 2355 636
rect 2237 437 2259 443
rect 2205 304 2211 356
rect 1949 264 1955 276
rect 1725 164 1731 256
rect 1866 214 1878 216
rect 1851 206 1853 214
rect 1861 206 1863 214
rect 1871 206 1873 214
rect 1881 206 1883 214
rect 1891 206 1893 214
rect 1866 204 1878 206
rect 1901 144 1907 156
rect 1485 44 1491 100
rect 1629 44 1635 100
rect 1261 -23 1283 -17
rect 1933 -23 1939 236
rect 1981 144 1987 236
rect 2029 184 2035 296
rect 2061 123 2067 256
rect 2109 184 2115 276
rect 2237 264 2243 437
rect 2397 384 2403 596
rect 2413 584 2419 616
rect 2429 604 2435 716
rect 2477 704 2483 717
rect 2493 704 2499 717
rect 2429 384 2435 536
rect 2445 524 2451 696
rect 2461 304 2467 636
rect 2493 504 2499 656
rect 2509 584 2515 736
rect 2477 484 2483 496
rect 2237 204 2243 256
rect 2285 164 2291 196
rect 2525 184 2531 516
rect 2541 284 2547 296
rect 2061 117 2076 123
rect 2077 104 2083 116
rect 2541 104 2547 256
rect 2189 44 2195 100
<< m3contact >>
rect 268 1776 276 1784
rect 476 1776 484 1784
rect 76 1756 84 1764
rect 12 1696 20 1704
rect 12 1496 20 1504
rect 76 1476 82 1484
rect 82 1476 84 1484
rect 412 1756 420 1764
rect 796 1756 804 1764
rect 444 1736 452 1744
rect 492 1736 500 1744
rect 764 1736 772 1744
rect 348 1716 356 1724
rect 668 1716 676 1724
rect 348 1496 356 1504
rect 236 1456 244 1464
rect 268 1416 276 1424
rect 76 1356 84 1364
rect 12 1296 20 1304
rect 12 1096 20 1104
rect 268 1336 276 1344
rect 412 1476 420 1484
rect 412 1356 420 1364
rect 428 1356 436 1364
rect 643 1606 651 1614
rect 653 1606 661 1614
rect 663 1606 671 1614
rect 673 1606 681 1614
rect 683 1606 691 1614
rect 693 1606 701 1614
rect 556 1576 564 1584
rect 684 1576 692 1584
rect 476 1496 484 1504
rect 508 1496 516 1504
rect 508 1436 516 1444
rect 604 1456 612 1464
rect 556 1416 564 1424
rect 572 1416 580 1424
rect 508 1356 516 1364
rect 700 1496 708 1504
rect 684 1376 692 1384
rect 748 1416 756 1424
rect 764 1376 772 1384
rect 908 1736 916 1744
rect 1100 1636 1108 1644
rect 844 1376 852 1384
rect 476 1336 484 1344
rect 796 1336 804 1344
rect 460 1316 468 1324
rect 540 1316 548 1324
rect 444 1236 452 1244
rect 428 1096 436 1104
rect 76 1056 84 1064
rect 268 1036 276 1044
rect 12 896 20 904
rect 76 896 84 904
rect 268 936 276 944
rect 428 1076 436 1084
rect 444 1036 452 1044
rect 444 956 452 964
rect 428 936 436 944
rect 364 916 372 924
rect 172 816 180 824
rect 236 816 244 824
rect 364 736 372 744
rect 412 736 420 744
rect 12 716 20 724
rect 76 716 84 724
rect 380 716 388 724
rect 60 676 68 684
rect 44 616 52 624
rect 396 696 404 704
rect 492 1296 500 1304
rect 508 1236 516 1244
rect 524 1116 532 1124
rect 620 1316 628 1324
rect 748 1296 756 1304
rect 620 1276 628 1284
rect 588 1176 596 1184
rect 604 1116 612 1124
rect 508 1076 516 1084
rect 540 1076 548 1084
rect 476 1056 484 1064
rect 588 1076 596 1084
rect 572 1056 580 1064
rect 604 1056 612 1064
rect 476 936 484 944
rect 460 716 468 724
rect 204 676 212 684
rect 428 676 436 684
rect 476 676 484 684
rect 348 616 356 624
rect 268 596 276 604
rect 316 596 324 604
rect 60 556 68 564
rect 92 556 100 564
rect 300 556 308 564
rect 12 496 20 504
rect 428 556 436 564
rect 380 536 388 544
rect 396 516 404 524
rect 12 296 20 304
rect 236 296 244 304
rect 268 296 276 304
rect 460 616 468 624
rect 588 896 596 904
rect 524 856 532 864
rect 508 736 516 744
rect 643 1206 651 1214
rect 653 1206 661 1214
rect 663 1206 671 1214
rect 673 1206 681 1214
rect 683 1206 691 1214
rect 693 1206 701 1214
rect 636 1176 644 1184
rect 652 1136 660 1144
rect 812 1316 820 1324
rect 780 1236 788 1244
rect 764 1216 772 1224
rect 1340 1816 1348 1824
rect 1260 1756 1268 1764
rect 1580 1756 1588 1764
rect 1692 1756 1700 1764
rect 1180 1636 1188 1644
rect 1036 1496 1044 1504
rect 924 1476 932 1484
rect 956 1476 964 1484
rect 988 1476 996 1484
rect 1068 1476 1076 1484
rect 1308 1636 1316 1644
rect 1228 1616 1236 1624
rect 1292 1616 1300 1624
rect 1196 1496 1204 1504
rect 1020 1456 1028 1464
rect 1084 1456 1092 1464
rect 972 1436 980 1444
rect 956 1396 964 1404
rect 1004 1396 1012 1404
rect 1212 1476 1220 1484
rect 1260 1476 1268 1484
rect 1116 1376 1124 1384
rect 1148 1376 1156 1384
rect 1116 1356 1124 1364
rect 860 1276 868 1284
rect 988 1296 996 1304
rect 1116 1296 1124 1304
rect 940 1216 948 1224
rect 796 1116 804 1124
rect 716 1096 724 1104
rect 748 1096 756 1104
rect 620 936 628 944
rect 892 1096 900 1104
rect 908 1076 916 1084
rect 748 1016 756 1024
rect 732 936 740 944
rect 780 1036 788 1044
rect 876 1036 884 1044
rect 764 996 772 1004
rect 1084 1076 1092 1084
rect 1356 1616 1364 1624
rect 1484 1696 1492 1704
rect 1436 1636 1444 1644
rect 1388 1556 1396 1564
rect 1468 1556 1476 1564
rect 1324 1496 1332 1504
rect 1372 1496 1380 1504
rect 1308 1396 1316 1404
rect 1404 1396 1412 1404
rect 1356 1356 1364 1364
rect 1388 1356 1396 1364
rect 1356 1336 1364 1344
rect 1276 1216 1284 1224
rect 1276 1176 1284 1184
rect 1660 1736 1668 1744
rect 1660 1716 1668 1724
rect 1843 1806 1851 1814
rect 1853 1806 1861 1814
rect 1863 1806 1871 1814
rect 1873 1806 1881 1814
rect 1883 1806 1891 1814
rect 1893 1806 1901 1814
rect 2156 1756 2164 1764
rect 2396 1756 2404 1764
rect 1836 1736 1844 1744
rect 2476 1736 2484 1744
rect 2028 1716 2036 1724
rect 1948 1596 1956 1604
rect 1980 1596 1988 1604
rect 1740 1496 1748 1504
rect 1804 1496 1812 1504
rect 1836 1496 1844 1504
rect 1932 1496 1940 1504
rect 1804 1476 1812 1484
rect 1756 1456 1764 1464
rect 1708 1436 1716 1444
rect 1740 1436 1748 1444
rect 1548 1416 1556 1424
rect 1612 1416 1620 1424
rect 1548 1396 1556 1404
rect 1580 1376 1588 1384
rect 1628 1356 1636 1364
rect 1660 1356 1668 1364
rect 1820 1456 1828 1464
rect 1843 1406 1851 1414
rect 1853 1406 1861 1414
rect 1863 1406 1871 1414
rect 1873 1406 1881 1414
rect 1883 1406 1891 1414
rect 1893 1406 1901 1414
rect 1820 1396 1828 1404
rect 1772 1336 1780 1344
rect 1356 1096 1364 1104
rect 1452 1096 1460 1104
rect 924 1016 932 1024
rect 796 996 804 1004
rect 764 976 772 984
rect 643 806 651 814
rect 653 806 661 814
rect 663 806 671 814
rect 673 806 681 814
rect 683 806 691 814
rect 693 806 701 814
rect 572 736 580 744
rect 604 736 612 744
rect 524 696 532 704
rect 748 856 756 864
rect 1164 996 1172 1004
rect 988 976 996 984
rect 1116 976 1124 984
rect 796 916 804 924
rect 556 676 564 684
rect 716 676 724 684
rect 652 656 660 664
rect 492 616 500 624
rect 620 596 628 604
rect 652 556 660 564
rect 460 536 468 544
rect 476 536 484 544
rect 444 316 452 324
rect 540 516 548 524
rect 508 316 516 324
rect 412 296 420 304
rect 476 296 484 304
rect 268 276 276 284
rect 76 256 84 264
rect 268 156 276 164
rect 76 136 82 144
rect 82 136 84 144
rect 428 276 436 284
rect 412 136 420 144
rect 476 256 484 264
rect 476 156 484 164
rect 556 296 564 304
rect 652 536 660 544
rect 748 516 756 524
rect 764 516 772 524
rect 643 406 651 414
rect 653 406 661 414
rect 663 406 671 414
rect 673 406 681 414
rect 683 406 691 414
rect 693 406 701 414
rect 1020 936 1028 944
rect 1132 916 1140 924
rect 972 756 980 764
rect 828 696 836 704
rect 1340 1076 1348 1084
rect 1308 1056 1316 1064
rect 1292 1036 1300 1044
rect 1436 1076 1444 1084
rect 1404 1016 1412 1024
rect 1324 976 1332 984
rect 1196 916 1204 924
rect 1292 916 1300 924
rect 1420 836 1428 844
rect 1244 776 1252 784
rect 1164 716 1172 724
rect 1228 716 1236 724
rect 1004 656 1012 664
rect 956 536 964 544
rect 1020 536 1028 544
rect 1036 536 1044 544
rect 1100 556 1108 564
rect 796 516 804 524
rect 828 516 836 524
rect 892 516 900 524
rect 940 516 948 524
rect 1004 516 1012 524
rect 780 376 788 384
rect 620 256 628 264
rect 764 276 772 284
rect 796 256 804 264
rect 748 196 756 204
rect 796 196 804 204
rect 1084 376 1092 384
rect 956 296 964 304
rect 988 296 996 304
rect 1020 296 1028 304
rect 1068 296 1076 304
rect 1388 716 1396 724
rect 1260 696 1268 704
rect 1356 676 1364 684
rect 1212 656 1220 664
rect 1388 596 1396 604
rect 1548 1196 1556 1204
rect 1484 1116 1492 1124
rect 1484 1096 1492 1104
rect 1516 1096 1524 1104
rect 1484 1076 1492 1084
rect 1500 1056 1508 1064
rect 1532 1056 1540 1064
rect 1564 1076 1572 1084
rect 1660 1296 1668 1304
rect 1628 1136 1636 1144
rect 1644 1116 1652 1124
rect 1612 1096 1620 1104
rect 1580 1056 1588 1064
rect 1596 1036 1604 1044
rect 1548 1016 1556 1024
rect 1596 1016 1604 1024
rect 1580 996 1588 1004
rect 1500 936 1508 944
rect 1468 916 1476 924
rect 1484 836 1492 844
rect 1452 816 1460 824
rect 1660 1076 1668 1084
rect 1740 1196 1748 1204
rect 2028 1496 2036 1504
rect 1948 1476 1956 1484
rect 1996 1456 2004 1464
rect 1948 1396 1956 1404
rect 1868 1376 1876 1384
rect 1772 1316 1780 1324
rect 1916 1356 1924 1364
rect 1900 1336 1908 1344
rect 2028 1356 2036 1364
rect 2076 1496 2084 1504
rect 2092 1476 2100 1484
rect 2076 1456 2084 1464
rect 2060 1376 2068 1384
rect 2044 1336 2052 1344
rect 1964 1316 1972 1324
rect 1996 1316 2004 1324
rect 2028 1316 2036 1324
rect 1788 1296 1796 1304
rect 2060 1296 2068 1304
rect 1996 1256 2004 1264
rect 2028 1256 2036 1264
rect 1740 1096 1748 1104
rect 1772 1096 1780 1104
rect 1964 1096 1972 1104
rect 1676 976 1684 984
rect 1708 996 1716 1004
rect 1788 1076 1796 1084
rect 1836 1076 1844 1084
rect 1900 1056 1908 1064
rect 1980 1056 1988 1064
rect 1772 1036 1780 1044
rect 1948 1016 1956 1024
rect 1843 1006 1851 1014
rect 1853 1006 1861 1014
rect 1863 1006 1871 1014
rect 1873 1006 1881 1014
rect 1883 1006 1891 1014
rect 1893 1006 1901 1014
rect 1708 976 1716 984
rect 1756 976 1764 984
rect 1964 976 1972 984
rect 1612 956 1620 964
rect 1644 956 1652 964
rect 1692 956 1700 964
rect 1804 956 1812 964
rect 2012 1116 2020 1124
rect 2044 1076 2052 1084
rect 2332 1536 2340 1544
rect 2364 1516 2372 1524
rect 2396 1516 2404 1524
rect 2188 1496 2196 1504
rect 2316 1496 2324 1504
rect 2156 1476 2164 1484
rect 2204 1476 2212 1484
rect 2316 1476 2324 1484
rect 2364 1476 2372 1484
rect 2108 1456 2116 1464
rect 2188 1396 2196 1404
rect 2108 1376 2116 1384
rect 2300 1456 2308 1464
rect 2236 1436 2244 1444
rect 2236 1376 2244 1384
rect 2156 1356 2164 1364
rect 2204 1356 2212 1364
rect 2268 1356 2276 1364
rect 2316 1356 2324 1364
rect 2124 1336 2132 1344
rect 2172 1336 2180 1344
rect 2204 1336 2212 1344
rect 2220 1316 2228 1324
rect 2268 1316 2276 1324
rect 2332 1316 2340 1324
rect 2140 1116 2148 1124
rect 2380 1456 2388 1464
rect 2380 1436 2388 1444
rect 2428 1556 2436 1564
rect 2444 1556 2452 1564
rect 2444 1536 2452 1544
rect 2540 1696 2548 1704
rect 2492 1676 2500 1684
rect 2508 1596 2516 1604
rect 2460 1516 2468 1524
rect 2540 1516 2548 1524
rect 2428 1496 2436 1504
rect 2508 1496 2516 1504
rect 2476 1456 2484 1464
rect 2412 1376 2420 1384
rect 2460 1376 2468 1384
rect 2364 1356 2372 1364
rect 2412 1356 2420 1364
rect 2444 1356 2452 1364
rect 2380 1316 2388 1324
rect 2380 1296 2388 1304
rect 2348 1136 2356 1144
rect 2028 1016 2036 1024
rect 2060 1016 2068 1024
rect 2012 976 2020 984
rect 1740 936 1748 944
rect 1980 936 1988 944
rect 1692 896 1700 904
rect 1596 876 1604 884
rect 1548 856 1556 864
rect 1548 776 1556 784
rect 1516 756 1524 764
rect 1548 756 1556 764
rect 1548 736 1556 744
rect 1724 856 1732 864
rect 1612 756 1620 764
rect 1484 716 1492 724
rect 1628 716 1636 724
rect 1500 676 1508 684
rect 1756 896 1764 904
rect 1884 916 1892 924
rect 1916 916 1924 924
rect 1996 916 2004 924
rect 1740 716 1748 724
rect 1932 896 1940 904
rect 1964 896 1972 904
rect 1916 816 1924 824
rect 1980 776 1988 784
rect 2220 1076 2228 1084
rect 2092 1056 2100 1064
rect 2124 1056 2132 1064
rect 2252 1056 2260 1064
rect 2076 976 2084 984
rect 2060 956 2068 964
rect 2076 876 2084 884
rect 2028 776 2036 784
rect 2012 756 2020 764
rect 2012 716 2020 724
rect 1548 676 1556 684
rect 1564 676 1572 684
rect 1628 676 1636 684
rect 1660 676 1668 684
rect 1772 676 1780 684
rect 2124 1036 2132 1044
rect 2108 976 2116 984
rect 2444 1276 2452 1284
rect 2396 1036 2404 1044
rect 2268 1016 2276 1024
rect 2380 1016 2388 1024
rect 2252 976 2260 984
rect 2284 976 2292 984
rect 2140 956 2148 964
rect 2172 956 2180 964
rect 2220 956 2228 964
rect 2172 896 2180 904
rect 2188 896 2196 904
rect 2108 876 2116 884
rect 2140 876 2148 884
rect 2236 936 2244 944
rect 2252 936 2260 944
rect 2300 936 2308 944
rect 2348 916 2356 924
rect 2412 1016 2420 1024
rect 2412 956 2420 964
rect 2476 1096 2484 1104
rect 2476 976 2484 984
rect 2460 956 2468 964
rect 2428 936 2436 944
rect 2444 916 2452 924
rect 2380 896 2388 904
rect 2172 776 2180 784
rect 2220 776 2228 784
rect 2220 756 2228 764
rect 2204 696 2212 704
rect 2396 736 2404 744
rect 2428 736 2436 744
rect 2460 736 2468 744
rect 2268 716 2276 724
rect 2444 716 2452 724
rect 2492 936 2500 944
rect 2508 916 2516 924
rect 2508 736 2516 744
rect 2284 696 2292 704
rect 2316 696 2324 704
rect 2300 676 2308 684
rect 1612 656 1620 664
rect 1676 656 1684 664
rect 1692 656 1700 664
rect 2252 656 2260 664
rect 2412 656 2420 664
rect 1740 636 1748 644
rect 1916 636 1924 644
rect 2172 636 2180 644
rect 1532 596 1540 604
rect 1372 556 1380 564
rect 1420 556 1428 564
rect 1388 536 1396 544
rect 1164 296 1172 304
rect 1244 296 1252 304
rect 1468 296 1476 304
rect 1020 276 1028 284
rect 1100 276 1108 284
rect 1004 236 1012 244
rect 940 176 948 184
rect 908 136 910 144
rect 910 136 916 144
rect 444 116 452 124
rect 524 116 532 124
rect 12 96 20 104
rect 643 6 651 14
rect 653 6 661 14
rect 663 6 671 14
rect 673 6 681 14
rect 683 6 691 14
rect 693 6 701 14
rect 1004 176 1012 184
rect 1292 276 1300 284
rect 1212 156 1220 164
rect 1116 116 1124 124
rect 1228 116 1234 124
rect 1234 116 1236 124
rect 1196 96 1204 104
rect 1244 96 1252 104
rect 1052 16 1060 24
rect 1100 16 1108 24
rect 1404 256 1412 264
rect 1843 606 1851 614
rect 1853 606 1861 614
rect 1863 606 1871 614
rect 1873 606 1881 614
rect 1883 606 1891 614
rect 1893 606 1901 614
rect 1740 596 1748 604
rect 1612 556 1620 564
rect 1548 476 1556 484
rect 1516 296 1524 304
rect 1484 276 1492 284
rect 1436 236 1444 244
rect 1420 156 1428 164
rect 1724 536 1732 544
rect 2044 596 2052 604
rect 2300 616 2308 624
rect 1964 536 1972 544
rect 1644 416 1652 424
rect 1692 416 1700 424
rect 1724 316 1732 324
rect 1964 516 1972 524
rect 2012 516 2020 524
rect 1964 496 1972 504
rect 2076 496 2084 504
rect 1996 476 2004 484
rect 2108 316 2116 324
rect 2412 616 2420 624
rect 2396 596 2404 604
rect 2348 496 2356 504
rect 1804 276 1806 284
rect 1806 276 1812 284
rect 1948 276 1956 284
rect 1644 256 1652 264
rect 1724 256 1732 264
rect 1900 236 1908 244
rect 1932 236 1940 244
rect 1843 206 1851 214
rect 1853 206 1861 214
rect 1863 206 1871 214
rect 1873 206 1881 214
rect 1883 206 1891 214
rect 1893 206 1901 214
rect 1884 156 1892 164
rect 1692 136 1700 144
rect 1900 136 1908 144
rect 1516 116 1524 124
rect 1596 116 1604 124
rect 2108 276 2116 284
rect 2204 276 2212 284
rect 2012 156 2020 164
rect 1980 136 1988 144
rect 2012 116 2020 124
rect 2044 116 2052 124
rect 2476 696 2484 704
rect 2428 596 2436 604
rect 2428 536 2436 544
rect 2460 636 2468 644
rect 2444 516 2452 524
rect 2524 656 2532 664
rect 2524 536 2532 544
rect 2524 516 2532 524
rect 2476 496 2484 504
rect 2236 256 2244 264
rect 2444 256 2452 264
rect 2236 196 2244 204
rect 2284 196 2292 204
rect 2540 296 2548 304
rect 2540 256 2548 264
rect 2252 136 2260 144
rect 2476 136 2484 144
rect 2156 116 2164 124
rect 2492 116 2500 124
rect 2076 96 2084 104
rect 2444 96 2452 104
rect 2540 96 2548 104
<< metal3 >>
rect 1348 1817 1356 1823
rect 1842 1814 1902 1816
rect 1842 1806 1843 1814
rect 1852 1806 1853 1814
rect 1891 1806 1892 1814
rect 1901 1806 1902 1814
rect 1842 1804 1902 1806
rect 276 1777 476 1783
rect 84 1757 412 1763
rect 804 1757 1260 1763
rect 1268 1757 1580 1763
rect 1588 1757 1692 1763
rect 1700 1757 2156 1763
rect 2164 1757 2188 1763
rect 2404 1757 2444 1763
rect 452 1737 492 1743
rect 772 1737 908 1743
rect 1668 1737 1836 1743
rect 2292 1737 2476 1743
rect 2484 1737 2579 1743
rect 356 1717 668 1723
rect 1668 1717 2028 1723
rect -35 1697 12 1703
rect 2548 1697 2579 1703
rect 2356 1677 2492 1683
rect 1108 1637 1180 1643
rect 1316 1637 1436 1643
rect 1236 1617 1292 1623
rect 642 1614 702 1616
rect 642 1606 643 1614
rect 652 1606 653 1614
rect 691 1606 692 1614
rect 701 1606 702 1614
rect 642 1604 702 1606
rect 1956 1597 1980 1603
rect 2516 1597 2579 1603
rect 564 1577 684 1583
rect 1396 1557 1468 1563
rect 2388 1557 2428 1563
rect 2452 1557 2476 1563
rect 2484 1557 2579 1563
rect 2340 1537 2444 1543
rect 2372 1517 2396 1523
rect 2468 1517 2540 1523
rect 2548 1517 2579 1523
rect -35 1497 12 1503
rect 356 1497 476 1503
rect 516 1497 700 1503
rect 884 1497 1036 1503
rect 1204 1497 1324 1503
rect 1332 1497 1372 1503
rect 1748 1497 1804 1503
rect 1844 1497 1932 1503
rect 2036 1497 2076 1503
rect 2084 1497 2188 1503
rect 2196 1497 2316 1503
rect 2436 1497 2508 1503
rect 84 1477 412 1483
rect 932 1477 956 1483
rect 996 1477 1068 1483
rect 1076 1477 1212 1483
rect 1220 1477 1260 1483
rect 1812 1477 1948 1483
rect 1997 1477 2092 1483
rect 1997 1464 2003 1477
rect 2100 1477 2156 1483
rect 2212 1477 2316 1483
rect 2324 1477 2364 1483
rect 2477 1477 2579 1483
rect 2477 1464 2483 1477
rect 244 1457 604 1463
rect 1028 1457 1084 1463
rect 1764 1457 1820 1463
rect 1828 1457 1996 1463
rect 2084 1457 2108 1463
rect 2308 1457 2380 1463
rect 2388 1457 2476 1463
rect 516 1437 972 1443
rect 1716 1437 1740 1443
rect 1780 1437 2236 1443
rect 2388 1437 2476 1443
rect 276 1417 556 1423
rect 580 1417 748 1423
rect 1556 1417 1612 1423
rect 1842 1414 1902 1416
rect 1842 1406 1843 1414
rect 1852 1406 1853 1414
rect 1891 1406 1892 1414
rect 1901 1406 1902 1414
rect 1842 1404 1902 1406
rect 964 1397 1004 1403
rect 1316 1397 1324 1403
rect 1412 1397 1548 1403
rect 1556 1397 1820 1403
rect 1956 1397 2188 1403
rect 692 1377 764 1383
rect 772 1377 844 1383
rect 1124 1377 1148 1383
rect 1588 1377 1772 1383
rect 1876 1377 2060 1383
rect 2116 1377 2236 1383
rect 2244 1377 2284 1383
rect 2365 1377 2412 1383
rect 2365 1364 2371 1377
rect 2420 1377 2460 1383
rect 84 1357 412 1363
rect 436 1357 508 1363
rect 1124 1357 1356 1363
rect 1373 1357 1388 1363
rect 276 1337 476 1343
rect 788 1337 796 1343
rect 1373 1343 1379 1357
rect 1636 1357 1660 1363
rect 1924 1357 2028 1363
rect 2164 1357 2204 1363
rect 2276 1357 2316 1363
rect 2388 1357 2412 1363
rect 2420 1357 2444 1363
rect 1364 1337 1379 1343
rect 1908 1337 2044 1343
rect 2052 1337 2124 1343
rect 2132 1337 2172 1343
rect 2381 1343 2387 1356
rect 2212 1337 2387 1343
rect 468 1317 540 1323
rect 548 1317 620 1323
rect 820 1317 876 1323
rect 1780 1317 1964 1323
rect 2004 1317 2028 1323
rect 2228 1317 2268 1323
rect 2340 1317 2380 1323
rect -35 1297 12 1303
rect 500 1297 748 1303
rect 996 1297 1116 1303
rect 1668 1297 1788 1303
rect 2068 1297 2348 1303
rect 2356 1297 2380 1303
rect 628 1277 860 1283
rect 2004 1257 2028 1263
rect 452 1237 508 1243
rect 516 1237 780 1243
rect 772 1217 940 1223
rect 948 1217 1276 1223
rect 642 1214 702 1216
rect 642 1206 643 1214
rect 652 1206 653 1214
rect 691 1206 692 1214
rect 701 1206 702 1214
rect 642 1204 702 1206
rect 1556 1197 1740 1203
rect 596 1177 636 1183
rect 1284 1177 1324 1183
rect -35 1137 652 1143
rect 1636 1137 2348 1143
rect 532 1117 604 1123
rect 612 1117 796 1123
rect 1492 1117 1644 1123
rect 2020 1117 2140 1123
rect -35 1097 12 1103
rect 724 1097 748 1103
rect 756 1097 892 1103
rect 1364 1097 1452 1103
rect 1492 1097 1516 1103
rect 1620 1097 1740 1103
rect 1748 1097 1772 1103
rect 1972 1097 2476 1103
rect 436 1077 508 1083
rect 548 1077 588 1083
rect 916 1077 1084 1083
rect 1348 1077 1436 1083
rect 1444 1077 1484 1083
rect 1492 1077 1564 1083
rect 1572 1077 1660 1083
rect 1796 1077 1836 1083
rect 2052 1077 2220 1083
rect 84 1057 476 1063
rect 580 1057 604 1063
rect 1316 1057 1500 1063
rect 1540 1057 1580 1063
rect 1908 1057 1980 1063
rect 2100 1057 2124 1063
rect 2196 1057 2252 1063
rect 276 1037 444 1043
rect 788 1037 876 1043
rect 1300 1037 1596 1043
rect 1780 1037 2124 1043
rect 2132 1037 2396 1043
rect 756 1017 924 1023
rect 932 1017 1004 1023
rect 1012 1017 1404 1023
rect 1412 1017 1548 1023
rect 1556 1017 1596 1023
rect 1956 1017 2028 1023
rect 2068 1017 2268 1023
rect 2388 1017 2412 1023
rect 1842 1014 1902 1016
rect 1842 1006 1843 1014
rect 1852 1006 1853 1014
rect 1891 1006 1892 1014
rect 1901 1006 1902 1014
rect 1842 1004 1902 1006
rect 772 997 796 1003
rect 1172 997 1580 1003
rect 1588 997 1708 1003
rect 1716 997 1772 1003
rect 772 977 780 983
rect 996 977 1116 983
rect 1124 977 1324 983
rect 1684 977 1708 983
rect 1716 977 1756 983
rect 1764 977 1964 983
rect 2020 977 2076 983
rect 2116 977 2252 983
rect 2292 977 2476 983
rect 436 957 444 963
rect 1620 957 1644 963
rect 1700 957 1804 963
rect 2068 957 2140 963
rect 2180 957 2220 963
rect 2420 957 2460 963
rect 276 937 428 943
rect 484 937 620 943
rect 740 937 1020 943
rect 1508 937 1740 943
rect 1748 937 1980 943
rect 1988 937 2236 943
rect 2260 937 2300 943
rect 2436 937 2492 943
rect 372 917 796 923
rect 1140 917 1196 923
rect 1300 917 1468 923
rect 1476 917 1884 923
rect 1924 917 1996 923
rect 2004 917 2348 923
rect 2452 917 2508 923
rect 2516 917 2579 923
rect -35 897 12 903
rect 84 897 588 903
rect 1700 897 1756 903
rect 1940 897 1964 903
rect 1972 897 2172 903
rect 2196 897 2380 903
rect 1604 877 2076 883
rect 2116 877 2140 883
rect 532 857 748 863
rect 1556 857 1724 863
rect 1428 837 1484 843
rect 180 817 236 823
rect 1460 817 1916 823
rect 642 814 702 816
rect 642 806 643 814
rect 652 806 653 814
rect 691 806 692 814
rect 701 806 702 814
rect 642 804 702 806
rect 1252 777 1548 783
rect 1988 777 2028 783
rect 2180 777 2220 783
rect 980 757 1516 763
rect 1556 757 1612 763
rect 1972 757 2012 763
rect 2020 757 2220 763
rect 372 737 412 743
rect 420 737 508 743
rect 580 737 604 743
rect 612 737 1548 743
rect 2404 737 2428 743
rect 2468 737 2508 743
rect -35 717 12 723
rect 84 717 380 723
rect 388 717 460 723
rect 1172 717 1228 723
rect 1396 717 1484 723
rect 1636 717 1740 723
rect 2020 717 2188 723
rect 2276 717 2444 723
rect 404 697 524 703
rect 836 697 1260 703
rect 2212 697 2284 703
rect 2324 697 2444 703
rect 2452 697 2476 703
rect -35 677 60 683
rect 68 677 204 683
rect 436 677 476 683
rect 484 677 556 683
rect 564 677 716 683
rect 1364 677 1500 683
rect 1508 677 1548 683
rect 1572 677 1628 683
rect 1668 677 1772 683
rect 1780 677 2300 683
rect 205 663 211 676
rect 205 657 652 663
rect 1012 657 1212 663
rect 1620 657 1676 663
rect 1700 657 2252 663
rect 2420 657 2476 663
rect 2484 657 2524 663
rect 2532 657 2579 663
rect 1748 637 1916 643
rect 2180 637 2460 643
rect 52 617 348 623
rect 356 617 460 623
rect 468 617 492 623
rect 2308 617 2412 623
rect 1842 614 1902 616
rect 1842 606 1843 614
rect 1852 606 1853 614
rect 1891 606 1892 614
rect 1901 606 1902 614
rect 1842 604 1902 606
rect 276 597 316 603
rect 324 597 620 603
rect 1396 597 1532 603
rect 1540 597 1740 603
rect 2052 597 2396 603
rect 2404 597 2428 603
rect 68 557 92 563
rect 308 557 428 563
rect 660 557 1100 563
rect 1380 557 1420 563
rect 1428 557 1612 563
rect 388 537 460 543
rect 484 537 652 543
rect 884 537 956 543
rect 964 537 1020 543
rect 1044 537 1388 543
rect 1732 537 1964 543
rect 2436 537 2524 543
rect 404 517 540 523
rect 756 517 764 523
rect 772 517 796 523
rect 836 517 892 523
rect 900 517 940 523
rect 1972 517 2012 523
rect 2452 517 2524 523
rect -35 497 12 503
rect 2084 497 2348 503
rect 2484 497 2579 503
rect 1556 477 1996 483
rect 1652 417 1692 423
rect 642 414 702 416
rect 642 406 643 414
rect 652 406 653 414
rect 691 406 692 414
rect 701 406 702 414
rect 642 404 702 406
rect 788 377 1084 383
rect 452 317 508 323
rect 1732 317 2108 323
rect 2116 317 2156 323
rect -35 297 12 303
rect 244 297 268 303
rect 420 297 476 303
rect 564 297 956 303
rect 996 297 1020 303
rect 1028 297 1068 303
rect 1076 297 1164 303
rect 1172 297 1244 303
rect 1476 297 1516 303
rect 2548 297 2579 303
rect 276 277 428 283
rect 772 277 1020 283
rect 1108 277 1292 283
rect 1492 277 1804 283
rect 1812 277 1948 283
rect 2116 277 2204 283
rect 84 257 476 263
rect 628 257 796 263
rect 1412 257 1644 263
rect 1652 257 1724 263
rect 1732 257 2236 263
rect 2452 257 2540 263
rect 1012 237 1436 243
rect 1908 237 1932 243
rect 1842 214 1902 216
rect 1842 206 1843 214
rect 1852 206 1853 214
rect 1891 206 1892 214
rect 1901 206 1902 214
rect 1842 204 1902 206
rect 756 197 796 203
rect 2244 197 2284 203
rect 948 177 1004 183
rect 276 157 476 163
rect 1220 157 1420 163
rect 1892 157 2012 163
rect 84 137 412 143
rect 916 137 1692 143
rect 1700 137 1900 143
rect 1988 137 2252 143
rect 452 117 524 123
rect 1124 117 1228 123
rect 1524 117 1596 123
rect 2020 117 2044 123
rect 2452 117 2492 123
rect -35 97 12 103
rect 1204 97 1244 103
rect 2084 97 2444 103
rect 2548 97 2579 103
rect 1060 17 1100 23
rect 642 14 702 16
rect 642 6 643 14
rect 652 6 653 14
rect 691 6 692 14
rect 701 6 702 14
rect 642 4 702 6
<< m4contact >>
rect 1356 1816 1364 1824
rect 1844 1806 1851 1814
rect 1851 1806 1852 1814
rect 1856 1806 1861 1814
rect 1861 1806 1863 1814
rect 1863 1806 1864 1814
rect 1868 1806 1871 1814
rect 1871 1806 1873 1814
rect 1873 1806 1876 1814
rect 1880 1806 1881 1814
rect 1881 1806 1883 1814
rect 1883 1806 1888 1814
rect 1892 1806 1893 1814
rect 1893 1806 1900 1814
rect 2188 1756 2196 1764
rect 2444 1756 2452 1764
rect 2284 1736 2292 1744
rect 1484 1696 1492 1704
rect 2348 1676 2356 1684
rect 1356 1616 1364 1624
rect 644 1606 651 1614
rect 651 1606 652 1614
rect 656 1606 661 1614
rect 661 1606 663 1614
rect 663 1606 664 1614
rect 668 1606 671 1614
rect 671 1606 673 1614
rect 673 1606 676 1614
rect 680 1606 681 1614
rect 681 1606 683 1614
rect 683 1606 688 1614
rect 692 1606 693 1614
rect 693 1606 700 1614
rect 2380 1556 2388 1564
rect 2476 1556 2484 1564
rect 876 1496 884 1504
rect 1772 1436 1780 1444
rect 2476 1436 2484 1444
rect 1844 1406 1851 1414
rect 1851 1406 1852 1414
rect 1856 1406 1861 1414
rect 1861 1406 1863 1414
rect 1863 1406 1864 1414
rect 1868 1406 1871 1414
rect 1871 1406 1873 1414
rect 1873 1406 1876 1414
rect 1880 1406 1881 1414
rect 1881 1406 1883 1414
rect 1883 1406 1888 1414
rect 1892 1406 1893 1414
rect 1893 1406 1900 1414
rect 1324 1396 1332 1404
rect 1772 1376 1780 1384
rect 2284 1376 2292 1384
rect 780 1336 788 1344
rect 2380 1356 2388 1364
rect 1772 1336 1780 1344
rect 876 1316 884 1324
rect 2348 1296 2356 1304
rect 2444 1276 2452 1284
rect 644 1206 651 1214
rect 651 1206 652 1214
rect 656 1206 661 1214
rect 661 1206 663 1214
rect 663 1206 664 1214
rect 668 1206 671 1214
rect 671 1206 673 1214
rect 673 1206 676 1214
rect 680 1206 681 1214
rect 681 1206 683 1214
rect 683 1206 688 1214
rect 692 1206 693 1214
rect 693 1206 700 1214
rect 1324 1176 1332 1184
rect 428 1096 436 1104
rect 1484 1076 1492 1084
rect 2188 1056 2196 1064
rect 1004 1016 1012 1024
rect 1844 1006 1851 1014
rect 1851 1006 1852 1014
rect 1856 1006 1861 1014
rect 1861 1006 1863 1014
rect 1863 1006 1864 1014
rect 1868 1006 1871 1014
rect 1871 1006 1873 1014
rect 1873 1006 1876 1014
rect 1880 1006 1881 1014
rect 1881 1006 1883 1014
rect 1883 1006 1888 1014
rect 1892 1006 1893 1014
rect 1893 1006 1900 1014
rect 1772 996 1780 1004
rect 780 976 788 984
rect 428 956 436 964
rect 644 806 651 814
rect 651 806 652 814
rect 656 806 661 814
rect 661 806 663 814
rect 663 806 664 814
rect 668 806 671 814
rect 671 806 673 814
rect 673 806 676 814
rect 680 806 681 814
rect 681 806 683 814
rect 683 806 688 814
rect 692 806 693 814
rect 693 806 700 814
rect 1964 756 1972 764
rect 2188 716 2196 724
rect 2444 696 2452 704
rect 2476 656 2484 664
rect 1844 606 1851 614
rect 1851 606 1852 614
rect 1856 606 1861 614
rect 1861 606 1863 614
rect 1863 606 1864 614
rect 1868 606 1871 614
rect 1871 606 1873 614
rect 1873 606 1876 614
rect 1880 606 1881 614
rect 1881 606 1883 614
rect 1883 606 1888 614
rect 1892 606 1893 614
rect 1893 606 1900 614
rect 876 536 884 544
rect 1004 516 1012 524
rect 1964 496 1972 504
rect 644 406 651 414
rect 651 406 652 414
rect 656 406 661 414
rect 661 406 663 414
rect 663 406 664 414
rect 668 406 671 414
rect 671 406 673 414
rect 673 406 676 414
rect 680 406 681 414
rect 681 406 683 414
rect 683 406 688 414
rect 692 406 693 414
rect 693 406 700 414
rect 2156 316 2164 324
rect 1844 206 1851 214
rect 1851 206 1852 214
rect 1856 206 1861 214
rect 1861 206 1863 214
rect 1863 206 1864 214
rect 1868 206 1871 214
rect 1871 206 1873 214
rect 1873 206 1876 214
rect 1880 206 1881 214
rect 1881 206 1883 214
rect 1883 206 1888 214
rect 1892 206 1893 214
rect 1893 206 1900 214
rect 2476 136 2484 144
rect 2156 116 2164 124
rect 2444 116 2452 124
rect 644 6 651 14
rect 651 6 652 14
rect 656 6 661 14
rect 661 6 663 14
rect 663 6 664 14
rect 668 6 671 14
rect 671 6 673 14
rect 673 6 676 14
rect 680 6 681 14
rect 681 6 683 14
rect 683 6 688 14
rect 692 6 693 14
rect 693 6 700 14
<< metal4 >>
rect 1354 1824 1366 1826
rect 1354 1816 1356 1824
rect 1364 1816 1366 1824
rect 640 1614 704 1816
rect 1354 1624 1366 1816
rect 1840 1814 1904 1816
rect 1840 1806 1844 1814
rect 1852 1806 1856 1814
rect 1864 1806 1868 1814
rect 1876 1806 1880 1814
rect 1888 1806 1892 1814
rect 1900 1806 1904 1814
rect 1354 1616 1356 1624
rect 1364 1616 1366 1624
rect 1354 1614 1366 1616
rect 1482 1704 1494 1706
rect 1482 1696 1484 1704
rect 1492 1696 1494 1704
rect 640 1606 644 1614
rect 652 1606 656 1614
rect 664 1606 668 1614
rect 676 1606 680 1614
rect 688 1606 692 1614
rect 700 1606 704 1614
rect 640 1214 704 1606
rect 874 1504 886 1506
rect 874 1496 876 1504
rect 884 1496 886 1504
rect 640 1206 644 1214
rect 652 1206 656 1214
rect 664 1206 668 1214
rect 676 1206 680 1214
rect 688 1206 692 1214
rect 700 1206 704 1214
rect 426 1104 438 1106
rect 426 1096 428 1104
rect 436 1096 438 1104
rect 426 964 438 1096
rect 426 956 428 964
rect 436 956 438 964
rect 426 954 438 956
rect 640 814 704 1206
rect 778 1344 790 1346
rect 778 1336 780 1344
rect 788 1336 790 1344
rect 778 984 790 1336
rect 778 976 780 984
rect 788 976 790 984
rect 778 974 790 976
rect 874 1324 886 1496
rect 874 1316 876 1324
rect 884 1316 886 1324
rect 640 806 644 814
rect 652 806 656 814
rect 664 806 668 814
rect 676 806 680 814
rect 688 806 692 814
rect 700 806 704 814
rect 640 414 704 806
rect 874 544 886 1316
rect 1322 1404 1334 1406
rect 1322 1396 1324 1404
rect 1332 1396 1334 1404
rect 1322 1184 1334 1396
rect 1322 1176 1324 1184
rect 1332 1176 1334 1184
rect 1322 1174 1334 1176
rect 1482 1084 1494 1696
rect 1770 1444 1782 1446
rect 1770 1436 1772 1444
rect 1780 1436 1782 1444
rect 1770 1384 1782 1436
rect 1770 1376 1772 1384
rect 1780 1376 1782 1384
rect 1770 1374 1782 1376
rect 1840 1414 1904 1806
rect 1840 1406 1844 1414
rect 1852 1406 1856 1414
rect 1864 1406 1868 1414
rect 1876 1406 1880 1414
rect 1888 1406 1892 1414
rect 1900 1406 1904 1414
rect 1482 1076 1484 1084
rect 1492 1076 1494 1084
rect 1482 1074 1494 1076
rect 1770 1344 1782 1346
rect 1770 1336 1772 1344
rect 1780 1336 1782 1344
rect 874 536 876 544
rect 884 536 886 544
rect 874 534 886 536
rect 1002 1024 1014 1026
rect 1002 1016 1004 1024
rect 1012 1016 1014 1024
rect 1002 524 1014 1016
rect 1770 1004 1782 1336
rect 1770 996 1772 1004
rect 1780 996 1782 1004
rect 1770 994 1782 996
rect 1840 1014 1904 1406
rect 1840 1006 1844 1014
rect 1852 1006 1856 1014
rect 1864 1006 1868 1014
rect 1876 1006 1880 1014
rect 1888 1006 1892 1014
rect 1900 1006 1904 1014
rect 1002 516 1004 524
rect 1012 516 1014 524
rect 1002 514 1014 516
rect 1840 614 1904 1006
rect 2186 1764 2198 1766
rect 2186 1756 2188 1764
rect 2196 1756 2198 1764
rect 2186 1064 2198 1756
rect 2442 1764 2454 1766
rect 2442 1756 2444 1764
rect 2452 1756 2454 1764
rect 2282 1744 2294 1746
rect 2282 1736 2284 1744
rect 2292 1736 2294 1744
rect 2282 1384 2294 1736
rect 2282 1376 2284 1384
rect 2292 1376 2294 1384
rect 2282 1374 2294 1376
rect 2346 1684 2358 1686
rect 2346 1676 2348 1684
rect 2356 1676 2358 1684
rect 2346 1304 2358 1676
rect 2378 1564 2390 1566
rect 2378 1556 2380 1564
rect 2388 1556 2390 1564
rect 2378 1364 2390 1556
rect 2378 1356 2380 1364
rect 2388 1356 2390 1364
rect 2378 1354 2390 1356
rect 2346 1296 2348 1304
rect 2356 1296 2358 1304
rect 2346 1294 2358 1296
rect 2442 1284 2454 1756
rect 2474 1564 2486 1566
rect 2474 1556 2476 1564
rect 2484 1556 2486 1564
rect 2474 1444 2486 1556
rect 2474 1436 2476 1444
rect 2484 1436 2486 1444
rect 2474 1434 2486 1436
rect 2442 1276 2444 1284
rect 2452 1276 2454 1284
rect 2442 1274 2454 1276
rect 2186 1056 2188 1064
rect 2196 1056 2198 1064
rect 1840 606 1844 614
rect 1852 606 1856 614
rect 1864 606 1868 614
rect 1876 606 1880 614
rect 1888 606 1892 614
rect 1900 606 1904 614
rect 640 406 644 414
rect 652 406 656 414
rect 664 406 668 414
rect 676 406 680 414
rect 688 406 692 414
rect 700 406 704 414
rect 640 14 704 406
rect 640 6 644 14
rect 652 6 656 14
rect 664 6 668 14
rect 676 6 680 14
rect 688 6 692 14
rect 700 6 704 14
rect 640 -10 704 6
rect 1840 214 1904 606
rect 1962 764 1974 766
rect 1962 756 1964 764
rect 1972 756 1974 764
rect 1962 504 1974 756
rect 2186 724 2198 1056
rect 2186 716 2188 724
rect 2196 716 2198 724
rect 2186 714 2198 716
rect 1962 496 1964 504
rect 1972 496 1974 504
rect 1962 494 1974 496
rect 2442 704 2454 706
rect 2442 696 2444 704
rect 2452 696 2454 704
rect 1840 206 1844 214
rect 1852 206 1856 214
rect 1864 206 1868 214
rect 1876 206 1880 214
rect 1888 206 1892 214
rect 1900 206 1904 214
rect 1840 -10 1904 206
rect 2154 324 2166 326
rect 2154 316 2156 324
rect 2164 316 2166 324
rect 2154 124 2166 316
rect 2154 116 2156 124
rect 2164 116 2166 124
rect 2154 114 2166 116
rect 2442 124 2454 696
rect 2474 664 2486 666
rect 2474 656 2476 664
rect 2484 656 2486 664
rect 2474 144 2486 656
rect 2474 136 2476 144
rect 2484 136 2486 144
rect 2474 134 2486 136
rect 2442 116 2444 124
rect 2452 116 2454 124
rect 2442 114 2454 116
use BUFX2  _312_
timestamp 1618241807
transform -1 0 56 0 -1 210
box -4 -6 52 206
use DFFSR  _285_
timestamp 1618241807
transform -1 0 408 0 -1 210
box -4 -6 356 206
use BUFX2  _313_
timestamp 1618241807
transform -1 0 56 0 1 210
box -4 -6 52 206
use DFFSR  _286_
timestamp 1618241807
transform -1 0 408 0 1 210
box -4 -6 356 206
use FILL  SFILL5360x100
timestamp 1618241807
transform -1 0 552 0 -1 210
box -4 -6 20 206
use FILL  SFILL5200x100
timestamp 1618241807
transform -1 0 536 0 -1 210
box -4 -6 20 206
use BUFX2  BUFX2_insert12
timestamp 1618241807
transform -1 0 568 0 1 210
box -4 -6 52 206
use NOR2X1  _240_
timestamp 1618241807
transform 1 0 472 0 1 210
box -4 -6 52 206
use AOI21X1  _241_
timestamp 1618241807
transform -1 0 472 0 1 210
box -4 -6 68 206
use AOI21X1  _238_
timestamp 1618241807
transform -1 0 520 0 -1 210
box -4 -6 68 206
use NOR2X1  _237_
timestamp 1618241807
transform 1 0 408 0 -1 210
box -4 -6 52 206
use FILL  SFILL6160x2100
timestamp 1618241807
transform 1 0 616 0 1 210
box -4 -6 20 206
use FILL  SFILL6000x2100
timestamp 1618241807
transform 1 0 600 0 1 210
box -4 -6 20 206
use FILL  SFILL5840x2100
timestamp 1618241807
transform 1 0 584 0 1 210
box -4 -6 20 206
use FILL  SFILL5680x2100
timestamp 1618241807
transform 1 0 568 0 1 210
box -4 -6 20 206
use FILL  SFILL5680x100
timestamp 1618241807
transform -1 0 584 0 -1 210
box -4 -6 20 206
use FILL  SFILL5520x100
timestamp 1618241807
transform -1 0 568 0 -1 210
box -4 -6 20 206
use DFFSR  _289_
timestamp 1618241807
transform 1 0 632 0 1 210
box -4 -6 356 206
use DFFSR  _273_
timestamp 1618241807
transform 1 0 584 0 -1 210
box -4 -6 356 206
use BUFX2  _316_
timestamp 1618241807
transform 1 0 936 0 -1 210
box -4 -6 52 206
use INVX8  _141_
timestamp 1618241807
transform -1 0 1064 0 -1 210
box -4 -6 84 206
use BUFX2  _310_
timestamp 1618241807
transform -1 0 1112 0 -1 210
box -4 -6 52 206
use NOR2X1  _249_
timestamp 1618241807
transform 1 0 984 0 1 210
box -4 -6 52 206
use AOI21X1  _250_
timestamp 1618241807
transform -1 0 1096 0 1 210
box -4 -6 68 206
use INVX1  _228_
timestamp 1618241807
transform 1 0 1112 0 -1 210
box -4 -6 36 206
use OAI21X1  _232_
timestamp 1618241807
transform 1 0 1144 0 -1 210
box -4 -6 68 206
use DFFSR  _283_
timestamp 1618241807
transform -1 0 1560 0 -1 210
box -4 -6 356 206
use CLKBUF1  CLKBUF1_insert1
timestamp 1618241807
transform 1 0 1096 0 1 210
box -4 -6 148 206
use NAND2X1  _231_
timestamp 1618241807
transform -1 0 1288 0 1 210
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert0
timestamp 1618241807
transform 1 0 1288 0 1 210
box -4 -6 148 206
use BUFX2  BUFX2_insert5
timestamp 1618241807
transform 1 0 1432 0 1 210
box -4 -6 52 206
use DFFSR  _274_
timestamp 1618241807
transform 1 0 1560 0 -1 210
box -4 -6 356 206
use DFFSR  _272_
timestamp 1618241807
transform 1 0 1480 0 1 210
box -4 -6 356 206
use FILL  SFILL18320x2100
timestamp 1618241807
transform 1 0 1832 0 1 210
box -4 -6 20 206
use FILL  SFILL18480x2100
timestamp 1618241807
transform 1 0 1848 0 1 210
box -4 -6 20 206
use FILL  SFILL18640x2100
timestamp 1618241807
transform 1 0 1864 0 1 210
box -4 -6 20 206
use FILL  SFILL18800x2100
timestamp 1618241807
transform 1 0 1880 0 1 210
box -4 -6 20 206
use BUFX2  _307_
timestamp 1618241807
transform -1 0 1944 0 1 210
box -4 -6 52 206
use INVX1  _152_
timestamp 1618241807
transform 1 0 1944 0 1 210
box -4 -6 36 206
use FILL  SFILL19120x100
timestamp 1618241807
transform -1 0 1928 0 -1 210
box -4 -6 20 206
use FILL  SFILL19280x100
timestamp 1618241807
transform -1 0 1944 0 -1 210
box -4 -6 20 206
use FILL  SFILL19440x100
timestamp 1618241807
transform -1 0 1960 0 -1 210
box -4 -6 20 206
use INVX1  _154_
timestamp 1618241807
transform 1 0 1976 0 -1 210
box -4 -6 36 206
use OAI21X1  _156_
timestamp 1618241807
transform -1 0 2040 0 1 210
box -4 -6 68 206
use FILL  SFILL19600x100
timestamp 1618241807
transform -1 0 1976 0 -1 210
box -4 -6 20 206
use INVX1  _153_
timestamp 1618241807
transform -1 0 2072 0 1 210
box -4 -6 36 206
use AND2X2  _157_
timestamp 1618241807
transform 1 0 2056 0 -1 210
box -4 -6 68 206
use NOR2X1  _155_
timestamp 1618241807
transform 1 0 2008 0 -1 210
box -4 -6 52 206
use DFFSR  _268_
timestamp 1618241807
transform 1 0 2072 0 1 210
box -4 -6 356 206
use DFFSR  _269_
timestamp 1618241807
transform 1 0 2120 0 -1 210
box -4 -6 356 206
use OAI21X1  _219_
timestamp 1618241807
transform 1 0 2472 0 -1 210
box -4 -6 68 206
use INVX1  _220_
timestamp 1618241807
transform -1 0 2456 0 1 210
box -4 -6 36 206
use BUFX2  _304_
timestamp 1618241807
transform 1 0 2456 0 1 210
box -4 -6 52 206
use FILL  FILL23760x2100
timestamp 1618241807
transform 1 0 2504 0 1 210
box -4 -6 20 206
use FILL  FILL23920x2100
timestamp 1618241807
transform 1 0 2520 0 1 210
box -4 -6 20 206
use BUFX2  _321_
timestamp 1618241807
transform -1 0 56 0 -1 610
box -4 -6 52 206
use INVX1  _239_
timestamp 1618241807
transform 1 0 56 0 -1 610
box -4 -6 36 206
use DFFSR  _295_
timestamp 1618241807
transform -1 0 440 0 -1 610
box -4 -6 356 206
use DFFSR  _296_
timestamp 1618241807
transform -1 0 792 0 -1 610
box -4 -6 356 206
use BUFX2  BUFX2_insert8
timestamp 1618241807
transform -1 0 904 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert9
timestamp 1618241807
transform -1 0 952 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert13
timestamp 1618241807
transform 1 0 952 0 -1 610
box -4 -6 52 206
use NOR2X1  _230_
timestamp 1618241807
transform -1 0 1048 0 -1 610
box -4 -6 52 206
use DFFSR  _270_
timestamp 1618241807
transform 1 0 1048 0 -1 610
box -4 -6 356 206
use FILL  SFILL7920x4100
timestamp 1618241807
transform -1 0 808 0 -1 610
box -4 -6 20 206
use FILL  SFILL8080x4100
timestamp 1618241807
transform -1 0 824 0 -1 610
box -4 -6 20 206
use FILL  SFILL8240x4100
timestamp 1618241807
transform -1 0 840 0 -1 610
box -4 -6 20 206
use FILL  SFILL8400x4100
timestamp 1618241807
transform -1 0 856 0 -1 610
box -4 -6 20 206
use INVX1  _229_
timestamp 1618241807
transform -1 0 1432 0 -1 610
box -4 -6 36 206
use NAND2X1  _257_
timestamp 1618241807
transform -1 0 1480 0 -1 610
box -4 -6 52 206
use INVX1  _215_
timestamp 1618241807
transform 1 0 1480 0 -1 610
box -4 -6 36 206
use DFFSR  _281_
timestamp 1618241807
transform -1 0 1864 0 -1 610
box -4 -6 356 206
use NAND2X1  _212_
timestamp 1618241807
transform 1 0 1928 0 -1 610
box -4 -6 52 206
use NAND3X1  _217_
timestamp 1618241807
transform -1 0 2040 0 -1 610
box -4 -6 68 206
use NAND2X1  _211_
timestamp 1618241807
transform 1 0 2040 0 -1 610
box -4 -6 52 206
use DFFSR  _282_
timestamp 1618241807
transform 1 0 2088 0 -1 610
box -4 -6 356 206
use FILL  SFILL18640x4100
timestamp 1618241807
transform -1 0 1880 0 -1 610
box -4 -6 20 206
use FILL  SFILL18800x4100
timestamp 1618241807
transform -1 0 1896 0 -1 610
box -4 -6 20 206
use FILL  SFILL18960x4100
timestamp 1618241807
transform -1 0 1912 0 -1 610
box -4 -6 20 206
use FILL  SFILL19120x4100
timestamp 1618241807
transform -1 0 1928 0 -1 610
box -4 -6 20 206
use BUFX2  _308_
timestamp 1618241807
transform 1 0 2440 0 -1 610
box -4 -6 52 206
use NAND2X1  _222_
timestamp 1618241807
transform -1 0 2536 0 -1 610
box -4 -6 52 206
use BUFX2  _322_
timestamp 1618241807
transform -1 0 56 0 1 610
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert4
timestamp 1618241807
transform 1 0 56 0 1 610
box -4 -6 148 206
use CLKBUF1  CLKBUF1_insert3
timestamp 1618241807
transform 1 0 200 0 1 610
box -4 -6 148 206
use INVX1  _242_
timestamp 1618241807
transform 1 0 344 0 1 610
box -4 -6 36 206
use OAI22X1  _267_
timestamp 1618241807
transform 1 0 376 0 1 610
box -4 -6 84 206
use OAI22X1  _136_
timestamp 1618241807
transform -1 0 536 0 1 610
box -4 -6 84 206
use INVX4  _265_
timestamp 1618241807
transform -1 0 584 0 1 610
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert2
timestamp 1618241807
transform 1 0 648 0 1 610
box -4 -6 148 206
use FILL  SFILL5840x6100
timestamp 1618241807
transform 1 0 584 0 1 610
box -4 -6 20 206
use FILL  SFILL6000x6100
timestamp 1618241807
transform 1 0 600 0 1 610
box -4 -6 20 206
use FILL  SFILL6160x6100
timestamp 1618241807
transform 1 0 616 0 1 610
box -4 -6 20 206
use FILL  SFILL6320x6100
timestamp 1618241807
transform 1 0 632 0 1 610
box -4 -6 20 206
use BUFX2  BUFX2_insert6
timestamp 1618241807
transform -1 0 840 0 1 610
box -4 -6 52 206
use DFFSR  _271_
timestamp 1618241807
transform 1 0 840 0 1 610
box -4 -6 356 206
use AND2X2  _158_
timestamp 1618241807
transform -1 0 1256 0 1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert7
timestamp 1618241807
transform 1 0 1256 0 1 610
box -4 -6 52 206
use NOR3X1  _213_
timestamp 1618241807
transform -1 0 1432 0 1 610
box -4 -6 132 206
use OAI21X1  _214_
timestamp 1618241807
transform 1 0 1432 0 1 610
box -4 -6 68 206
use OAI21X1  _216_
timestamp 1618241807
transform 1 0 1496 0 1 610
box -4 -6 68 206
use OAI21X1  _225_
timestamp 1618241807
transform 1 0 1560 0 1 610
box -4 -6 68 206
use NAND2X1  _224_
timestamp 1618241807
transform -1 0 1672 0 1 610
box -4 -6 52 206
use AOI21X1  _226_
timestamp 1618241807
transform -1 0 1736 0 1 610
box -4 -6 68 206
use NOR2X1  _147_
timestamp 1618241807
transform 1 0 1736 0 1 610
box -4 -6 52 206
use FILL  SFILL17840x6100
timestamp 1618241807
transform 1 0 1784 0 1 610
box -4 -6 20 206
use FILL  SFILL18000x6100
timestamp 1618241807
transform 1 0 1800 0 1 610
box -4 -6 20 206
use DFFSR  _278_
timestamp 1618241807
transform 1 0 1848 0 1 610
box -4 -6 356 206
use FILL  SFILL18160x6100
timestamp 1618241807
transform 1 0 1816 0 1 610
box -4 -6 20 206
use FILL  SFILL18320x6100
timestamp 1618241807
transform 1 0 1832 0 1 610
box -4 -6 20 206
use AOI22X1  _227_
timestamp 1618241807
transform 1 0 2200 0 1 610
box -4 -6 84 206
use INVX1  _218_
timestamp 1618241807
transform -1 0 2312 0 1 610
box -4 -6 36 206
use XOR2X1  _210_
timestamp 1618241807
transform 1 0 2312 0 1 610
box -4 -6 116 206
use NAND3X1  _223_
timestamp 1618241807
transform 1 0 2424 0 1 610
box -4 -6 68 206
use NOR2X1  _221_
timestamp 1618241807
transform -1 0 2536 0 1 610
box -4 -6 52 206
use BUFX2  _323_
timestamp 1618241807
transform -1 0 56 0 -1 1010
box -4 -6 52 206
use DFFSR  _297_
timestamp 1618241807
transform -1 0 408 0 -1 1010
box -4 -6 356 206
use OAI22X1  _137_
timestamp 1618241807
transform -1 0 488 0 -1 1010
box -4 -6 84 206
use XOR2X1  _261_
timestamp 1618241807
transform -1 0 600 0 -1 1010
box -4 -6 116 206
use INVX1  _245_
timestamp 1618241807
transform 1 0 600 0 -1 1010
box -4 -6 36 206
use OAI22X1  _138_
timestamp 1618241807
transform -1 0 776 0 -1 1010
box -4 -6 84 206
use FILL  SFILL6320x8100
timestamp 1618241807
transform -1 0 648 0 -1 1010
box -4 -6 20 206
use FILL  SFILL6480x8100
timestamp 1618241807
transform -1 0 664 0 -1 1010
box -4 -6 20 206
use FILL  SFILL6640x8100
timestamp 1618241807
transform -1 0 680 0 -1 1010
box -4 -6 20 206
use FILL  SFILL6800x8100
timestamp 1618241807
transform -1 0 696 0 -1 1010
box -4 -6 20 206
use INVX1  _248_
timestamp 1618241807
transform -1 0 808 0 -1 1010
box -4 -6 36 206
use DFFSR  _298_
timestamp 1618241807
transform -1 0 1160 0 -1 1010
box -4 -6 356 206
use DFFSR  _280_
timestamp 1618241807
transform 1 0 1160 0 -1 1010
box -4 -6 356 206
use OAI21X1  _151_
timestamp 1618241807
transform -1 0 1576 0 -1 1010
box -4 -6 68 206
use INVX1  _142_
timestamp 1618241807
transform 1 0 1576 0 -1 1010
box -4 -6 36 206
use NOR2X1  _196_
timestamp 1618241807
transform -1 0 1656 0 -1 1010
box -4 -6 52 206
use NOR2X1  _148_
timestamp 1618241807
transform 1 0 1656 0 -1 1010
box -4 -6 52 206
use NOR2X1  _150_
timestamp 1618241807
transform 1 0 1704 0 -1 1010
box -4 -6 52 206
use NAND2X1  _149_
timestamp 1618241807
transform -1 0 1800 0 -1 1010
box -4 -6 52 206
use INVX1  _194_
timestamp 1618241807
transform 1 0 1800 0 -1 1010
box -4 -6 36 206
use NAND3X1  _204_
timestamp 1618241807
transform 1 0 1896 0 -1 1010
box -4 -6 68 206
use NAND2X1  _146_
timestamp 1618241807
transform -1 0 2008 0 -1 1010
box -4 -6 52 206
use OAI21X1  _192_
timestamp 1618241807
transform 1 0 2008 0 -1 1010
box -4 -6 68 206
use OAI21X1  _183_
timestamp 1618241807
transform -1 0 2136 0 -1 1010
box -4 -6 68 206
use NAND2X1  _184_
timestamp 1618241807
transform -1 0 2184 0 -1 1010
box -4 -6 52 206
use FILL  SFILL18320x8100
timestamp 1618241807
transform -1 0 1848 0 -1 1010
box -4 -6 20 206
use FILL  SFILL18480x8100
timestamp 1618241807
transform -1 0 1864 0 -1 1010
box -4 -6 20 206
use FILL  SFILL18640x8100
timestamp 1618241807
transform -1 0 1880 0 -1 1010
box -4 -6 20 206
use FILL  SFILL18800x8100
timestamp 1618241807
transform -1 0 1896 0 -1 1010
box -4 -6 20 206
use NOR2X1  _145_
timestamp 1618241807
transform -1 0 2232 0 -1 1010
box -4 -6 52 206
use AOI21X1  _180_
timestamp 1618241807
transform 1 0 2232 0 -1 1010
box -4 -6 68 206
use AND2X2  _179_
timestamp 1618241807
transform -1 0 2360 0 -1 1010
box -4 -6 68 206
use INVX1  _178_
timestamp 1618241807
transform -1 0 2392 0 -1 1010
box -4 -6 36 206
use OAI21X1  _176_
timestamp 1618241807
transform -1 0 2456 0 -1 1010
box -4 -6 68 206
use AOI21X1  _177_
timestamp 1618241807
transform -1 0 2520 0 -1 1010
box -4 -6 68 206
use FILL  FILL23920x8100
timestamp 1618241807
transform -1 0 2536 0 -1 1010
box -4 -6 20 206
use BUFX2  _314_
timestamp 1618241807
transform -1 0 56 0 1 1010
box -4 -6 52 206
use DFFSR  _287_
timestamp 1618241807
transform -1 0 408 0 1 1010
box -4 -6 356 206
use AOI21X1  _244_
timestamp 1618241807
transform 1 0 408 0 1 1010
box -4 -6 68 206
use NOR2X1  _243_
timestamp 1618241807
transform 1 0 472 0 1 1010
box -4 -6 52 206
use OAI21X1  _263_
timestamp 1618241807
transform 1 0 520 0 1 1010
box -4 -6 68 206
use AND2X2  _262_
timestamp 1618241807
transform 1 0 584 0 1 1010
box -4 -6 68 206
use BUFX2  _324_
timestamp 1618241807
transform -1 0 760 0 1 1010
box -4 -6 52 206
use FILL  SFILL6480x10100
timestamp 1618241807
transform 1 0 648 0 1 1010
box -4 -6 20 206
use FILL  SFILL6640x10100
timestamp 1618241807
transform 1 0 664 0 1 1010
box -4 -6 20 206
use FILL  SFILL6800x10100
timestamp 1618241807
transform 1 0 680 0 1 1010
box -4 -6 20 206
use FILL  SFILL6960x10100
timestamp 1618241807
transform 1 0 696 0 1 1010
box -4 -6 20 206
use XNOR2X1  _260_
timestamp 1618241807
transform -1 0 872 0 1 1010
box -4 -6 116 206
use OAI22X1  _139_
timestamp 1618241807
transform -1 0 952 0 1 1010
box -4 -6 84 206
use DFFSR  _299_
timestamp 1618241807
transform 1 0 952 0 1 1010
box -4 -6 356 206
use AND2X2  _205_
timestamp 1618241807
transform -1 0 1368 0 1 1010
box -4 -6 68 206
use OAI21X1  _259_
timestamp 1618241807
transform -1 0 1432 0 1 1010
box -4 -6 68 206
use OAI21X1  _206_
timestamp 1618241807
transform 1 0 1432 0 1 1010
box -4 -6 68 206
use OAI22X1  _207_
timestamp 1618241807
transform -1 0 1576 0 1 1010
box -4 -6 84 206
use AOI21X1  _208_
timestamp 1618241807
transform -1 0 1640 0 1 1010
box -4 -6 68 206
use OAI21X1  _197_
timestamp 1618241807
transform -1 0 1704 0 1 1010
box -4 -6 68 206
use NOR2X1  _159_
timestamp 1618241807
transform 1 0 1704 0 1 1010
box -4 -6 52 206
use INVX1  _185_
timestamp 1618241807
transform 1 0 1752 0 1 1010
box -4 -6 36 206
use NOR2X1  _195_
timestamp 1618241807
transform -1 0 1832 0 1 1010
box -4 -6 52 206
use AOI22X1  _191_
timestamp 1618241807
transform 1 0 1896 0 1 1010
box -4 -6 84 206
use NOR2X1  _190_
timestamp 1618241807
transform 1 0 1976 0 1 1010
box -4 -6 52 206
use OAI21X1  _181_
timestamp 1618241807
transform -1 0 2088 0 1 1010
box -4 -6 68 206
use DFFSR  _277_
timestamp 1618241807
transform 1 0 2088 0 1 1010
box -4 -6 356 206
use FILL  SFILL18320x10100
timestamp 1618241807
transform 1 0 1832 0 1 1010
box -4 -6 20 206
use FILL  SFILL18480x10100
timestamp 1618241807
transform 1 0 1848 0 1 1010
box -4 -6 20 206
use FILL  SFILL18640x10100
timestamp 1618241807
transform 1 0 1864 0 1 1010
box -4 -6 20 206
use FILL  SFILL18800x10100
timestamp 1618241807
transform 1 0 1880 0 1 1010
box -4 -6 20 206
use OAI21X1  _186_
timestamp 1618241807
transform 1 0 2440 0 1 1010
box -4 -6 68 206
use FILL  FILL23760x10100
timestamp 1618241807
transform 1 0 2504 0 1 1010
box -4 -6 20 206
use FILL  FILL23920x10100
timestamp 1618241807
transform 1 0 2520 0 1 1010
box -4 -6 20 206
use BUFX2  _320_
timestamp 1618241807
transform -1 0 56 0 -1 1410
box -4 -6 52 206
use DFFSR  _294_
timestamp 1618241807
transform -1 0 408 0 -1 1410
box -4 -6 356 206
use INVX1  _236_
timestamp 1618241807
transform 1 0 408 0 -1 1410
box -4 -6 36 206
use OAI22X1  _266_
timestamp 1618241807
transform 1 0 440 0 -1 1410
box -4 -6 84 206
use OAI22X1  _264_
timestamp 1618241807
transform 1 0 520 0 -1 1410
box -4 -6 84 206
use INVX1  _254_
timestamp 1618241807
transform -1 0 632 0 -1 1410
box -4 -6 36 206
use OAI22X1  _140_
timestamp 1618241807
transform 1 0 696 0 -1 1410
box -4 -6 84 206
use FILL  SFILL6320x12100
timestamp 1618241807
transform -1 0 648 0 -1 1410
box -4 -6 20 206
use FILL  SFILL6480x12100
timestamp 1618241807
transform -1 0 664 0 -1 1410
box -4 -6 20 206
use FILL  SFILL6640x12100
timestamp 1618241807
transform -1 0 680 0 -1 1410
box -4 -6 20 206
use FILL  SFILL6800x12100
timestamp 1618241807
transform -1 0 696 0 -1 1410
box -4 -6 20 206
use BUFX2  BUFX2_insert11
timestamp 1618241807
transform -1 0 824 0 -1 1410
box -4 -6 52 206
use DFFSR  _284_
timestamp 1618241807
transform 1 0 824 0 -1 1410
box -4 -6 356 206
use DFFSR  _292_
timestamp 1618241807
transform -1 0 1528 0 -1 1410
box -4 -6 356 206
use INVX4  _143_
timestamp 1618241807
transform -1 0 1576 0 -1 1410
box -4 -6 52 206
use AOI21X1  _199_
timestamp 1618241807
transform 1 0 1576 0 -1 1410
box -4 -6 68 206
use OAI22X1  _198_
timestamp 1618241807
transform -1 0 1720 0 -1 1410
box -4 -6 84 206
use INVX4  _182_
timestamp 1618241807
transform -1 0 1768 0 -1 1410
box -4 -6 52 206
use OAI21X1  _164_
timestamp 1618241807
transform 1 0 1768 0 -1 1410
box -4 -6 68 206
use FILL  SFILL18800x12100
timestamp 1618241807
transform -1 0 1896 0 -1 1410
box -4 -6 20 206
use FILL  SFILL18640x12100
timestamp 1618241807
transform -1 0 1880 0 -1 1410
box -4 -6 20 206
use FILL  SFILL18480x12100
timestamp 1618241807
transform -1 0 1864 0 -1 1410
box -4 -6 20 206
use FILL  SFILL18320x12100
timestamp 1618241807
transform -1 0 1848 0 -1 1410
box -4 -6 20 206
use AOI21X1  _171_
timestamp 1618241807
transform 1 0 1896 0 -1 1410
box -4 -6 68 206
use OAI21X1  _174_
timestamp 1618241807
transform 1 0 2008 0 -1 1410
box -4 -6 68 206
use NOR2X1  _173_
timestamp 1618241807
transform 1 0 1960 0 -1 1410
box -4 -6 52 206
use OAI21X1  _161_
timestamp 1618241807
transform -1 0 2136 0 -1 1410
box -4 -6 68 206
use AOI21X1  _170_
timestamp 1618241807
transform -1 0 2232 0 -1 1410
box -4 -6 68 206
use INVX1  _189_
timestamp 1618241807
transform -1 0 2168 0 -1 1410
box -4 -6 36 206
use INVX1  _166_
timestamp 1618241807
transform 1 0 2232 0 -1 1410
box -4 -6 36 206
use NAND2X1  _168_
timestamp 1618241807
transform 1 0 2264 0 -1 1410
box -4 -6 52 206
use OAI21X1  _188_
timestamp 1618241807
transform 1 0 2312 0 -1 1410
box -4 -6 68 206
use INVX1  _167_
timestamp 1618241807
transform 1 0 2376 0 -1 1410
box -4 -6 36 206
use INVX1  _175_
timestamp 1618241807
transform 1 0 2408 0 -1 1410
box -4 -6 36 206
use NAND3X1  _209_
timestamp 1618241807
transform 1 0 2440 0 -1 1410
box -4 -6 68 206
use FILL  FILL23760x12100
timestamp 1618241807
transform -1 0 2520 0 -1 1410
box -4 -6 20 206
use FILL  FILL23920x12100
timestamp 1618241807
transform -1 0 2536 0 -1 1410
box -4 -6 20 206
use BUFX2  _319_
timestamp 1618241807
transform -1 0 56 0 1 1410
box -4 -6 52 206
use DFFSR  _293_
timestamp 1618241807
transform -1 0 408 0 1 1410
box -4 -6 356 206
use INVX1  _233_
timestamp 1618241807
transform 1 0 408 0 1 1410
box -4 -6 36 206
use DFFSR  _300_
timestamp 1618241807
transform 1 0 440 0 1 1410
box -4 -6 356 206
use AOI21X1  _247_
timestamp 1618241807
transform 1 0 856 0 1 1410
box -4 -6 68 206
use NOR2X1  _246_
timestamp 1618241807
transform 1 0 920 0 1 1410
box -4 -6 52 206
use AOI21X1  _235_
timestamp 1618241807
transform 1 0 968 0 1 1410
box -4 -6 68 206
use BUFX2  BUFX2_insert10
timestamp 1618241807
transform 1 0 1032 0 1 1410
box -4 -6 52 206
use NOR2X1  _234_
timestamp 1618241807
transform -1 0 1128 0 1 1410
box -4 -6 52 206
use FILL  SFILL7920x14100
timestamp 1618241807
transform 1 0 792 0 1 1410
box -4 -6 20 206
use FILL  SFILL8080x14100
timestamp 1618241807
transform 1 0 808 0 1 1410
box -4 -6 20 206
use FILL  SFILL8240x14100
timestamp 1618241807
transform 1 0 824 0 1 1410
box -4 -6 20 206
use FILL  SFILL8400x14100
timestamp 1618241807
transform 1 0 840 0 1 1410
box -4 -6 20 206
use BUFX2  _311_
timestamp 1618241807
transform 1 0 1128 0 1 1410
box -4 -6 52 206
use NOR2X1  _252_
timestamp 1618241807
transform 1 0 1176 0 1 1410
box -4 -6 52 206
use AOI21X1  _253_
timestamp 1618241807
transform -1 0 1288 0 1 1410
box -4 -6 68 206
use INVX1  _251_
timestamp 1618241807
transform -1 0 1320 0 1 1410
box -4 -6 36 206
use BUFX2  _309_
timestamp 1618241807
transform 1 0 1320 0 1 1410
box -4 -6 52 206
use NAND2X1  _258_
timestamp 1618241807
transform 1 0 1368 0 1 1410
box -4 -6 52 206
use DFFSR  _279_
timestamp 1618241807
transform 1 0 1416 0 1 1410
box -4 -6 356 206
use BUFX2  _305_
timestamp 1618241807
transform -1 0 1816 0 1 1410
box -4 -6 52 206
use FILL  SFILL18800x14100
timestamp 1618241807
transform 1 0 1880 0 1 1410
box -4 -6 20 206
use OAI21X1  _172_
timestamp 1618241807
transform 1 0 1816 0 1 1410
box -4 -6 68 206
use FILL  SFILL19280x14100
timestamp 1618241807
transform 1 0 1928 0 1 1410
box -4 -6 20 206
use FILL  SFILL19120x14100
timestamp 1618241807
transform 1 0 1912 0 1 1410
box -4 -6 20 206
use FILL  SFILL18960x14100
timestamp 1618241807
transform 1 0 1896 0 1 1410
box -4 -6 20 206
use NAND2X1  _165_
timestamp 1618241807
transform -1 0 1992 0 1 1410
box -4 -6 52 206
use NOR2X1  _144_
timestamp 1618241807
transform 1 0 1992 0 1 1410
box -4 -6 52 206
use OAI21X1  _163_
timestamp 1618241807
transform 1 0 2088 0 1 1410
box -4 -6 68 206
use NAND2X1  _160_
timestamp 1618241807
transform -1 0 2088 0 1 1410
box -4 -6 52 206
use NAND2X1  _162_
timestamp 1618241807
transform -1 0 2200 0 1 1410
box -4 -6 52 206
use XNOR2X1  _193_
timestamp 1618241807
transform 1 0 2200 0 1 1410
box -4 -6 116 206
use OAI21X1  _203_
timestamp 1618241807
transform 1 0 2312 0 1 1410
box -4 -6 68 206
use OAI21X1  _200_
timestamp 1618241807
transform 1 0 2376 0 1 1410
box -4 -6 68 206
use INVX1  _202_
timestamp 1618241807
transform -1 0 2472 0 1 1410
box -4 -6 36 206
use NOR2X1  _201_
timestamp 1618241807
transform 1 0 2472 0 1 1410
box -4 -6 52 206
use FILL  FILL23920x14100
timestamp 1618241807
transform 1 0 2520 0 1 1410
box -4 -6 20 206
use BUFX2  _318_
timestamp 1618241807
transform -1 0 56 0 -1 1810
box -4 -6 52 206
use DFFSR  _291_
timestamp 1618241807
transform -1 0 408 0 -1 1810
box -4 -6 356 206
use NOR2X1  _255_
timestamp 1618241807
transform 1 0 408 0 -1 1810
box -4 -6 52 206
use AOI21X1  _256_
timestamp 1618241807
transform -1 0 520 0 -1 1810
box -4 -6 68 206
use BUFX2  _326_
timestamp 1618241807
transform -1 0 568 0 -1 1810
box -4 -6 52 206
use DFFSR  _288_
timestamp 1618241807
transform 1 0 632 0 -1 1810
box -4 -6 356 206
use FILL  SFILL5680x16100
timestamp 1618241807
transform -1 0 584 0 -1 1810
box -4 -6 20 206
use FILL  SFILL5840x16100
timestamp 1618241807
transform -1 0 600 0 -1 1810
box -4 -6 20 206
use FILL  SFILL6000x16100
timestamp 1618241807
transform -1 0 616 0 -1 1810
box -4 -6 20 206
use FILL  SFILL6160x16100
timestamp 1618241807
transform -1 0 632 0 -1 1810
box -4 -6 20 206
use BUFX2  _315_
timestamp 1618241807
transform 1 0 984 0 -1 1810
box -4 -6 52 206
use BUFX2  _317_
timestamp 1618241807
transform -1 0 1080 0 -1 1810
box -4 -6 52 206
use DFFSR  _290_
timestamp 1618241807
transform -1 0 1432 0 -1 1810
box -4 -6 356 206
use BUFX2  _325_
timestamp 1618241807
transform 1 0 1432 0 -1 1810
box -4 -6 52 206
use BUFX2  _306_
timestamp 1618241807
transform 1 0 1480 0 -1 1810
box -4 -6 52 206
use DFFSR  _276_
timestamp 1618241807
transform 1 0 1528 0 -1 1810
box -4 -6 356 206
use BUFX2  _302_
timestamp 1618241807
transform 1 0 1944 0 -1 1810
box -4 -6 52 206
use DFFSR  _275_
timestamp 1618241807
transform 1 0 1992 0 -1 1810
box -4 -6 356 206
use FILL  SFILL18800x16100
timestamp 1618241807
transform -1 0 1896 0 -1 1810
box -4 -6 20 206
use FILL  SFILL18960x16100
timestamp 1618241807
transform -1 0 1912 0 -1 1810
box -4 -6 20 206
use FILL  SFILL19120x16100
timestamp 1618241807
transform -1 0 1928 0 -1 1810
box -4 -6 20 206
use FILL  SFILL19280x16100
timestamp 1618241807
transform -1 0 1944 0 -1 1810
box -4 -6 20 206
use BUFX2  _301_
timestamp 1618241807
transform 1 0 2344 0 -1 1810
box -4 -6 52 206
use NOR2X1  _187_
timestamp 1618241807
transform 1 0 2392 0 -1 1810
box -4 -6 52 206
use NAND2X1  _169_
timestamp 1618241807
transform -1 0 2488 0 -1 1810
box -4 -6 52 206
use BUFX2  _303_
timestamp 1618241807
transform 1 0 2488 0 -1 1810
box -4 -6 52 206
<< labels >>
flabel metal4 s 1840 -10 1904 0 7 FreeSans 24 270 0 0 gnd
port 0 nsew
flabel metal4 s 640 -10 704 0 7 FreeSans 24 270 0 0 vdd
port 1 nsew
flabel metal3 s 2573 97 2579 103 3 FreeSans 24 0 0 0 N[8]
port 2 nsew
flabel metal3 s 2573 657 2579 663 3 FreeSans 24 0 0 0 N[7]
port 3 nsew
flabel metal3 s 2573 1597 2579 1603 3 FreeSans 24 0 0 0 N[6]
port 4 nsew
flabel metal3 s 2573 1477 2579 1483 3 FreeSans 24 0 0 0 N[5]
port 5 nsew
flabel metal3 s 2573 1517 2579 1523 3 FreeSans 24 0 0 0 N[4]
port 6 nsew
flabel metal3 s 2573 917 2579 923 3 FreeSans 24 0 0 0 N[3]
port 7 nsew
flabel metal3 s 2573 1557 2579 1563 3 FreeSans 24 0 0 0 N[2]
port 8 nsew
flabel metal3 s 2573 1737 2579 1743 3 FreeSans 24 0 0 0 N[1]
port 9 nsew
flabel metal2 s 1261 -23 1267 -17 7 FreeSans 24 270 0 0 N[0]
port 10 nsew
flabel metal3 s -35 677 -29 683 7 FreeSans 24 0 0 0 clock
port 11 nsew
flabel metal3 s 2573 497 2579 503 3 FreeSans 24 0 0 0 counter[7]
port 12 nsew
flabel metal2 s 1933 -23 1939 -17 7 FreeSans 24 270 0 0 counter[6]
port 13 nsew
flabel metal2 s 1501 1857 1507 1863 3 FreeSans 24 90 0 0 counter[5]
port 14 nsew
flabel metal2 s 1789 1857 1795 1863 3 FreeSans 24 90 0 0 counter[4]
port 15 nsew
flabel metal3 s 2573 297 2579 303 3 FreeSans 24 0 0 0 counter[3]
port 16 nsew
flabel metal3 s 2573 1697 2579 1703 3 FreeSans 24 0 0 0 counter[2]
port 17 nsew
flabel metal2 s 1965 1857 1971 1863 3 FreeSans 24 90 0 0 counter[1]
port 18 nsew
flabel metal2 s 2365 1857 2371 1863 3 FreeSans 24 90 0 0 counter[0]
port 19 nsew
flabel metal2 s 1341 1857 1347 1863 3 FreeSans 24 90 0 0 done
port 20 nsew
flabel metal3 s -35 1697 -29 1703 7 FreeSans 24 0 0 0 dp[8]
port 21 nsew
flabel metal2 s 1053 1857 1059 1863 3 FreeSans 24 90 0 0 dp[7]
port 22 nsew
flabel metal2 s 957 -23 963 -17 7 FreeSans 24 270 0 0 dp[6]
port 23 nsew
flabel metal2 s 1005 1857 1011 1863 3 FreeSans 24 90 0 0 dp[5]
port 24 nsew
flabel metal3 s -35 1097 -29 1103 7 FreeSans 24 0 0 0 dp[4]
port 25 nsew
flabel metal3 s -35 297 -29 303 7 FreeSans 24 0 0 0 dp[3]
port 26 nsew
flabel metal3 s -35 97 -29 103 7 FreeSans 24 0 0 0 dp[2]
port 27 nsew
flabel metal2 s 1149 1857 1155 1863 3 FreeSans 24 90 0 0 dp[1]
port 28 nsew
flabel metal2 s 1069 -23 1075 -17 7 FreeSans 24 270 0 0 dp[0]
port 29 nsew
flabel metal2 s 1101 -23 1107 -17 7 FreeSans 24 270 0 0 reset
port 30 nsew
flabel metal2 s 541 1857 547 1863 3 FreeSans 24 90 0 0 sr[7]
port 31 nsew
flabel metal2 s 1453 1857 1459 1863 3 FreeSans 24 90 0 0 sr[6]
port 32 nsew
flabel metal3 s -35 1137 -29 1143 7 FreeSans 24 0 0 0 sr[5]
port 33 nsew
flabel metal3 s -35 897 -29 903 7 FreeSans 24 0 0 0 sr[4]
port 34 nsew
flabel metal3 s -35 717 -29 723 7 FreeSans 24 0 0 0 sr[3]
port 35 nsew
flabel metal3 s -35 497 -29 503 7 FreeSans 24 0 0 0 sr[2]
port 36 nsew
flabel metal3 s -35 1297 -29 1303 7 FreeSans 24 0 0 0 sr[1]
port 37 nsew
flabel metal3 s -35 1497 -29 1503 7 FreeSans 24 0 0 0 sr[0]
port 38 nsew
flabel metal2 s 749 -23 755 -17 7 FreeSans 24 270 0 0 start
port 39 nsew
<< end >>
