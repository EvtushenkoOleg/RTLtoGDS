magic
tech scmos
magscale 1 2
timestamp 1618002947
<< metal1 >>
rect 2746 3814 2758 3816
rect 2731 3806 2733 3814
rect 2741 3806 2743 3814
rect 2751 3806 2753 3814
rect 2761 3806 2763 3814
rect 2771 3806 2773 3814
rect 2746 3804 2758 3806
rect 3805 3757 3843 3763
rect 2221 3737 2243 3743
rect 2372 3737 2387 3743
rect 3380 3737 3395 3743
rect 3156 3717 3171 3723
rect 3204 3717 3219 3723
rect 3828 3717 3859 3723
rect 2228 3697 2243 3703
rect 3245 3697 3260 3703
rect 20 3677 35 3683
rect 1805 3677 1820 3683
rect 2330 3676 2332 3684
rect 2404 3677 2420 3683
rect 2932 3677 2948 3683
rect 3108 3677 3123 3683
rect 5076 3677 5091 3683
rect 1242 3614 1254 3616
rect 4250 3614 4262 3616
rect 1227 3606 1229 3614
rect 1237 3606 1239 3614
rect 1247 3606 1249 3614
rect 1257 3606 1259 3614
rect 1267 3606 1269 3614
rect 4235 3606 4237 3614
rect 4245 3606 4247 3614
rect 4255 3606 4257 3614
rect 4265 3606 4267 3614
rect 4275 3606 4277 3614
rect 1242 3604 1254 3606
rect 4250 3604 4262 3606
rect 3610 3576 3612 3584
rect 3690 3576 3692 3584
rect 4804 3576 4806 3584
rect 5050 3576 5052 3584
rect 4740 3556 4742 3564
rect 3396 3537 3427 3543
rect 3754 3536 3756 3544
rect 4500 3536 4502 3544
rect 365 3497 403 3503
rect 525 3497 563 3503
rect 932 3497 947 3503
rect 3085 3497 3100 3503
rect 3581 3503 3587 3523
rect 4644 3516 4652 3524
rect 4893 3517 4915 3523
rect 3549 3497 3587 3503
rect 4333 3497 4364 3503
rect 4628 3497 4643 3503
rect 3165 3477 3180 3483
rect 3460 3477 3491 3483
rect 3501 3477 3516 3483
rect 509 3457 524 3463
rect 909 3457 940 3463
rect 3501 3457 3507 3477
rect 4221 3477 4323 3483
rect 4061 3457 4076 3463
rect 2746 3414 2758 3416
rect 2731 3406 2733 3414
rect 2741 3406 2743 3414
rect 2751 3406 2753 3414
rect 2761 3406 2763 3414
rect 2771 3406 2773 3414
rect 2746 3404 2758 3406
rect 3828 3376 3830 3384
rect 756 3356 764 3364
rect 2125 3344 2131 3363
rect 3581 3357 3603 3363
rect 4141 3357 4163 3363
rect 4173 3357 4188 3363
rect 4196 3357 4236 3363
rect 4244 3357 4275 3363
rect 5197 3357 5212 3363
rect 5252 3357 5267 3363
rect 685 3337 723 3343
rect 781 3337 819 3343
rect 1700 3337 1715 3343
rect 1805 3337 1843 3343
rect 1940 3337 1955 3343
rect 2132 3337 2163 3343
rect 3444 3337 3459 3343
rect 3709 3337 3731 3343
rect 3748 3337 3779 3343
rect 3789 3337 3804 3343
rect 3821 3337 3859 3343
rect 4180 3337 4291 3343
rect 413 3317 451 3323
rect 445 3297 451 3317
rect 621 3317 636 3323
rect 1789 3317 1804 3323
rect 2173 3317 2210 3323
rect 3693 3317 3708 3323
rect 4093 3323 4099 3336
rect 4525 3324 4531 3343
rect 4973 3337 4995 3343
rect 5277 3337 5299 3343
rect 4093 3317 4115 3323
rect 4148 3317 4163 3323
rect 4532 3317 4547 3323
rect 4957 3317 4972 3323
rect 5117 3317 5148 3323
rect 1837 3297 1859 3303
rect 3988 3297 4003 3303
rect 4013 3297 4051 3303
rect 4980 3297 4995 3303
rect 5380 3296 5388 3304
rect 5405 3297 5427 3303
rect 52 3277 67 3283
rect 3421 3277 3436 3283
rect 4074 3256 4076 3264
rect 3690 3236 3692 3244
rect 1242 3214 1254 3216
rect 4250 3214 4262 3216
rect 1227 3206 1229 3214
rect 1237 3206 1239 3214
rect 1247 3206 1249 3214
rect 1257 3206 1259 3214
rect 1267 3206 1269 3214
rect 4235 3206 4237 3214
rect 4245 3206 4247 3214
rect 4255 3206 4257 3214
rect 4265 3206 4267 3214
rect 4275 3206 4277 3214
rect 1242 3204 1254 3206
rect 4250 3204 4262 3206
rect 298 3176 300 3184
rect 452 3176 454 3184
rect 692 3176 694 3184
rect 1412 3176 1414 3184
rect 1946 3176 1948 3184
rect 2452 3176 2454 3184
rect 540 3137 595 3143
rect 540 3132 548 3137
rect 3354 3136 3356 3144
rect 4084 3137 4115 3143
rect 205 3117 220 3123
rect 948 3116 956 3124
rect 676 3097 691 3103
rect 973 3103 979 3123
rect 932 3097 947 3103
rect 973 3097 1011 3103
rect 1133 3097 1148 3103
rect 1181 3097 1204 3103
rect 1196 3092 1204 3097
rect 1372 3103 1380 3108
rect 1372 3097 1395 3103
rect 1389 3077 1395 3097
rect 1716 3097 1747 3103
rect 1853 3103 1859 3123
rect 1853 3097 1891 3103
rect 2045 3103 2051 3123
rect 2228 3117 2243 3123
rect 3492 3116 3500 3124
rect 2045 3097 2083 3103
rect 3517 3103 3523 3123
rect 3885 3117 3916 3123
rect 4372 3117 4387 3123
rect 5380 3116 5388 3124
rect 3517 3097 3555 3103
rect 3661 3097 3683 3103
rect 3741 3097 3756 3103
rect 3796 3097 3811 3103
rect 4328 3096 4332 3104
rect 5181 3097 5196 3103
rect 1773 3077 1827 3083
rect 1972 3077 1987 3083
rect 2004 3077 2019 3083
rect 2221 3077 2259 3083
rect 2317 3077 2339 3083
rect 2388 3077 2403 3083
rect 2413 3077 2435 3083
rect 20 3057 35 3063
rect 1133 3057 1155 3063
rect 1165 3057 1180 3063
rect 2397 3057 2403 3077
rect 3389 3077 3404 3083
rect 3908 3077 3923 3083
rect 4132 3077 4163 3083
rect 4173 3077 4291 3083
rect 4173 3064 4179 3077
rect 5053 3077 5084 3083
rect 5101 3077 5107 3096
rect 5277 3077 5292 3083
rect 5453 3077 5516 3083
rect 3764 3056 3772 3064
rect 4125 3057 4140 3063
rect 4196 3057 4275 3063
rect 4733 3057 4771 3063
rect 104 3036 108 3044
rect 173 3037 188 3043
rect 580 3037 595 3043
rect 1245 3037 1260 3043
rect 1341 3037 1356 3043
rect 1844 3036 1846 3044
rect 2036 3036 2038 3044
rect 5434 3036 5436 3044
rect 2746 3014 2758 3016
rect 2731 3006 2733 3014
rect 2741 3006 2743 3014
rect 2751 3006 2753 3014
rect 2761 3006 2763 3014
rect 2771 3006 2773 3014
rect 2746 3004 2758 3006
rect 1668 2976 1670 2984
rect 2020 2976 2022 2984
rect 2212 2976 2214 2984
rect 2669 2977 2700 2983
rect 3261 2977 3276 2983
rect 3586 2977 3628 2983
rect 4068 2976 4070 2984
rect 5098 2976 5100 2984
rect 93 2957 108 2963
rect 148 2957 163 2963
rect 1092 2956 1100 2964
rect 3501 2957 3539 2963
rect 3620 2957 3651 2963
rect 317 2937 332 2943
rect 1117 2937 1139 2943
rect 1300 2937 1315 2943
rect 1389 2937 1411 2943
rect 1789 2937 1804 2943
rect 1853 2937 1875 2943
rect 2109 2937 2140 2943
rect 2605 2937 2627 2943
rect 3325 2937 3347 2943
rect 3453 2937 3475 2943
rect 3485 2937 3516 2943
rect 3469 2924 3475 2937
rect 3540 2937 3555 2943
rect 4004 2937 4019 2943
rect 4036 2937 4051 2943
rect 4125 2937 4179 2943
rect 4397 2937 4451 2943
rect 4477 2943 4483 2963
rect 5140 2957 5155 2963
rect 4468 2937 4483 2943
rect 1268 2917 1331 2923
rect 1341 2917 1372 2923
rect 1684 2917 1715 2923
rect 1805 2917 1843 2923
rect 2157 2917 2195 2923
rect 2477 2917 2492 2923
rect 2509 2917 2531 2923
rect 3389 2917 3427 2923
rect 1860 2897 1875 2903
rect 3389 2897 3395 2917
rect 3844 2917 3859 2923
rect 3869 2917 3907 2923
rect 4196 2917 4211 2923
rect 4973 2917 4988 2923
rect 29 2877 83 2883
rect 173 2877 188 2883
rect 1229 2877 1292 2883
rect 3261 2877 3308 2883
rect 1242 2814 1254 2816
rect 4250 2814 4262 2816
rect 1227 2806 1229 2814
rect 1237 2806 1239 2814
rect 1247 2806 1249 2814
rect 1257 2806 1259 2814
rect 1267 2806 1269 2814
rect 4235 2806 4237 2814
rect 4245 2806 4247 2814
rect 4255 2806 4257 2814
rect 4265 2806 4267 2814
rect 4275 2806 4277 2814
rect 1242 2804 1254 2806
rect 4250 2804 4262 2806
rect 2084 2776 2086 2784
rect 388 2736 390 2744
rect 1684 2737 1699 2743
rect 1708 2737 1740 2743
rect 1708 2732 1716 2737
rect 1866 2736 1868 2744
rect 4157 2737 4172 2743
rect 589 2717 604 2723
rect 509 2697 524 2703
rect 740 2697 787 2703
rect 1869 2697 1884 2703
rect 2148 2697 2179 2703
rect 2237 2697 2268 2703
rect 5436 2703 5444 2706
rect 797 2683 803 2696
rect 5436 2697 5459 2703
rect 797 2677 819 2683
rect 1230 2677 1324 2683
rect 1373 2677 1388 2683
rect 1437 2677 1459 2683
rect 1501 2677 1539 2683
rect 1597 2677 1635 2683
rect 2205 2677 2227 2683
rect 2285 2677 2307 2683
rect 2461 2677 2483 2683
rect 4317 2677 4332 2683
rect 5364 2676 5366 2684
rect 5485 2677 5516 2683
rect 3357 2657 3395 2663
rect 4509 2657 4547 2663
rect 458 2636 460 2644
rect 618 2636 620 2644
rect 2746 2614 2758 2616
rect 2731 2606 2733 2614
rect 2741 2606 2743 2614
rect 2751 2606 2753 2614
rect 2761 2606 2763 2614
rect 2771 2606 2773 2614
rect 2746 2604 2758 2606
rect 2426 2576 2428 2584
rect 1245 2557 1324 2563
rect 1917 2557 1939 2563
rect 2045 2557 2060 2563
rect 3869 2557 3884 2563
rect 3892 2557 3907 2563
rect 637 2543 643 2556
rect 621 2537 643 2543
rect 29 2517 44 2523
rect 221 2517 236 2523
rect 324 2517 339 2523
rect 605 2517 636 2523
rect 669 2517 684 2523
rect 781 2517 796 2523
rect 1332 2517 1347 2523
rect 1837 2523 1843 2543
rect 1981 2537 2012 2543
rect 2445 2537 2482 2543
rect 3421 2537 3443 2543
rect 1837 2517 1875 2523
rect 1965 2517 1980 2523
rect 3261 2517 3299 2523
rect 3325 2517 3356 2523
rect 3293 2504 3299 2517
rect 5324 2504 5332 2514
rect 3821 2477 3836 2483
rect 772 2456 774 2464
rect 394 2436 396 2444
rect 660 2436 662 2444
rect 1242 2414 1254 2416
rect 4250 2414 4262 2416
rect 1227 2406 1229 2414
rect 1237 2406 1239 2414
rect 1247 2406 1249 2414
rect 1257 2406 1259 2414
rect 1267 2406 1269 2414
rect 4235 2406 4237 2414
rect 4245 2406 4247 2414
rect 4255 2406 4257 2414
rect 4265 2406 4267 2414
rect 4275 2406 4277 2414
rect 1242 2404 1254 2406
rect 4250 2404 4262 2406
rect 1946 2376 1948 2384
rect 3220 2376 3222 2384
rect 3572 2376 3574 2384
rect 5501 2377 5516 2383
rect 701 2343 707 2363
rect 701 2337 716 2343
rect 1677 2337 1708 2343
rect 1757 2337 1772 2343
rect 2052 2337 2067 2343
rect 4228 2337 4316 2343
rect 4404 2337 4435 2343
rect 452 2316 460 2324
rect 1556 2316 1564 2324
rect 4205 2317 4268 2323
rect 4397 2317 4412 2323
rect 4468 2317 4483 2323
rect 4900 2317 4915 2323
rect 1565 2297 1580 2303
rect 1885 2297 1916 2303
rect 3380 2297 3411 2303
rect 3492 2297 3507 2303
rect 3741 2297 3772 2303
rect 5428 2297 5443 2303
rect 516 2277 531 2283
rect 893 2283 899 2296
rect 836 2277 883 2283
rect 893 2277 915 2283
rect 1668 2277 1683 2283
rect 3444 2277 3459 2283
rect 4141 2277 4163 2283
rect 4708 2277 4723 2283
rect 4804 2277 4819 2283
rect 5348 2277 5372 2283
rect 628 2256 636 2264
rect 2029 2257 2044 2263
rect 2404 2257 2419 2263
rect 2772 2257 2819 2263
rect 676 2236 680 2244
rect 2746 2214 2758 2216
rect 2731 2206 2733 2214
rect 2741 2206 2743 2214
rect 2751 2206 2753 2214
rect 2761 2206 2763 2214
rect 2771 2206 2773 2214
rect 2746 2204 2758 2206
rect 154 2176 156 2184
rect 562 2176 572 2184
rect 1085 2177 1132 2183
rect 2100 2176 2102 2184
rect 792 2157 819 2163
rect 1524 2157 1539 2163
rect 1700 2156 1708 2164
rect 2381 2157 2403 2163
rect 2868 2157 2883 2163
rect 4397 2157 4412 2163
rect 77 2137 115 2143
rect 29 2117 60 2123
rect 109 2117 115 2137
rect 157 2137 172 2143
rect 196 2137 211 2143
rect 909 2137 940 2143
rect 980 2137 995 2143
rect 1684 2137 1699 2143
rect 1725 2137 1740 2143
rect 1869 2137 1907 2143
rect 2132 2137 2156 2143
rect 2317 2137 2355 2143
rect 3277 2137 3299 2143
rect 3405 2137 3420 2143
rect 3773 2137 3788 2143
rect 4164 2137 4179 2143
rect 4221 2137 4236 2143
rect 4292 2137 4323 2143
rect 1486 2117 1516 2123
rect 1661 2117 1683 2123
rect 1661 2104 1667 2117
rect 2237 2117 2268 2123
rect 2381 2117 2396 2123
rect 2429 2117 2460 2123
rect 3341 2117 3379 2123
rect 3341 2097 3347 2117
rect 3757 2117 3772 2123
rect 4205 2117 4284 2123
rect 4532 2117 4579 2123
rect 4701 2117 4716 2123
rect 260 2077 300 2083
rect 1924 2076 1926 2084
rect 4442 2076 4444 2084
rect 4500 2076 4502 2084
rect 5469 2077 5500 2083
rect 4010 2036 4012 2044
rect 4138 2036 4140 2044
rect 1242 2014 1254 2016
rect 4250 2014 4262 2016
rect 1227 2006 1229 2014
rect 1237 2006 1239 2014
rect 1247 2006 1249 2014
rect 1257 2006 1259 2014
rect 1267 2006 1269 2014
rect 4235 2006 4237 2014
rect 4245 2006 4247 2014
rect 4255 2006 4257 2014
rect 4265 2006 4267 2014
rect 4275 2006 4277 2014
rect 1242 2004 1254 2006
rect 4250 2004 4262 2006
rect 4212 1976 4214 1984
rect 4650 1976 4652 1984
rect 5082 1976 5084 1984
rect 5156 1976 5158 1984
rect 5428 1976 5430 1984
rect 4236 1937 4300 1943
rect 4573 1937 4604 1943
rect 2253 1917 2275 1923
rect 228 1897 243 1903
rect 2173 1897 2188 1903
rect 2397 1903 2403 1923
rect 3812 1917 3827 1923
rect 4317 1917 4332 1923
rect 2365 1897 2403 1903
rect 4180 1897 4211 1903
rect 5316 1897 5331 1903
rect 5453 1903 5459 1923
rect 5453 1897 5491 1903
rect 125 1877 163 1883
rect 356 1877 372 1883
rect 364 1876 372 1877
rect 1805 1877 1820 1883
rect 2429 1877 2451 1883
rect 2461 1877 2483 1883
rect 2525 1877 2563 1883
rect 2573 1877 2668 1883
rect 2445 1864 2451 1877
rect 3389 1877 3411 1883
rect 4572 1877 4588 1883
rect 4572 1876 4580 1877
rect 2589 1857 2636 1863
rect 3812 1857 3827 1863
rect 3956 1856 3964 1864
rect 74 1836 76 1844
rect 2746 1814 2758 1816
rect 2731 1806 2733 1814
rect 2741 1806 2743 1814
rect 2751 1806 2753 1814
rect 2761 1806 2763 1814
rect 2771 1806 2773 1814
rect 2746 1804 2758 1806
rect 360 1776 364 1784
rect 522 1776 524 1784
rect 2538 1776 2540 1784
rect 4872 1776 4876 1784
rect 109 1757 124 1763
rect 173 1757 188 1763
rect 1892 1757 1923 1763
rect 4116 1757 4195 1763
rect 989 1737 1043 1743
rect 1949 1737 1987 1743
rect 2397 1737 2435 1743
rect 3357 1737 3379 1743
rect 3549 1737 3587 1743
rect 4589 1737 4604 1743
rect 5005 1737 5020 1743
rect 29 1717 51 1723
rect 61 1717 92 1723
rect 941 1717 972 1723
rect 1012 1717 1027 1723
rect 1085 1717 1100 1723
rect 2749 1717 2812 1723
rect 2932 1717 2962 1723
rect 3421 1717 3459 1723
rect 3469 1717 3484 1723
rect 308 1697 323 1703
rect 500 1697 515 1703
rect 3421 1697 3427 1717
rect 4564 1717 4595 1723
rect 5229 1717 5235 1736
rect 4780 1712 4788 1716
rect 4036 1697 4051 1703
rect 269 1677 300 1683
rect 308 1677 316 1683
rect 324 1677 355 1683
rect 4020 1677 4044 1683
rect 4074 1636 4076 1644
rect 4538 1636 4540 1644
rect 1242 1614 1254 1616
rect 4250 1614 4262 1616
rect 1227 1606 1229 1614
rect 1237 1606 1239 1614
rect 1247 1606 1249 1614
rect 1257 1606 1259 1614
rect 1267 1606 1269 1614
rect 4235 1606 4237 1614
rect 4245 1606 4247 1614
rect 4255 1606 4257 1614
rect 4265 1606 4267 1614
rect 4275 1606 4277 1614
rect 1242 1604 1254 1606
rect 4250 1604 4262 1606
rect 3546 1576 3548 1584
rect 4970 1576 4972 1584
rect 84 1537 99 1543
rect 1908 1537 1923 1543
rect 4580 1537 4636 1543
rect 5124 1537 5139 1543
rect 292 1497 307 1503
rect 637 1503 643 1523
rect 2564 1517 2579 1523
rect 2861 1517 2883 1523
rect 3245 1517 3260 1523
rect 3892 1517 3907 1523
rect 4589 1517 4604 1523
rect 596 1497 611 1503
rect 637 1497 675 1503
rect 2141 1497 2179 1503
rect 3549 1497 3580 1503
rect 3661 1497 3676 1503
rect 4413 1497 4444 1503
rect 5229 1497 5244 1503
rect 221 1477 275 1483
rect 221 1457 227 1477
rect 452 1477 499 1483
rect 580 1477 595 1483
rect 637 1477 652 1483
rect 685 1477 722 1483
rect 1092 1477 1107 1483
rect 1117 1477 1139 1483
rect 1806 1477 1843 1483
rect 1885 1477 1907 1483
rect 1940 1477 1971 1483
rect 1981 1477 2035 1483
rect 2084 1477 2099 1483
rect 2628 1477 2643 1483
rect 2804 1477 2819 1483
rect 2925 1477 2962 1483
rect 3341 1477 3363 1483
rect 3572 1477 3587 1483
rect 3780 1477 3795 1483
rect 4141 1477 4179 1483
rect 4276 1477 4356 1483
rect 5485 1477 5516 1483
rect 372 1457 387 1463
rect 1085 1457 1091 1476
rect 4524 1472 4532 1476
rect 4548 1456 4552 1464
rect 84 1437 99 1443
rect 2746 1414 2758 1416
rect 2731 1406 2733 1414
rect 2741 1406 2743 1414
rect 2751 1406 2753 1414
rect 2761 1406 2763 1414
rect 2771 1406 2773 1414
rect 2746 1404 2758 1406
rect 1754 1376 1756 1384
rect 2637 1377 2652 1383
rect 1805 1357 1820 1363
rect 3549 1357 3564 1363
rect 125 1343 131 1356
rect 109 1337 131 1343
rect 141 1337 172 1343
rect 1485 1337 1507 1343
rect 1645 1337 1676 1343
rect 1773 1337 1795 1343
rect 2477 1337 2492 1343
rect 2532 1337 2563 1343
rect 877 1317 899 1323
rect 1732 1317 1747 1323
rect 1485 1297 1500 1303
rect 1741 1297 1747 1317
rect 2205 1317 2243 1323
rect 2253 1317 2268 1323
rect 2276 1317 2300 1323
rect 2340 1317 2355 1323
rect 2589 1323 2595 1343
rect 3117 1337 3139 1343
rect 3597 1337 3612 1343
rect 3773 1343 3779 1363
rect 5156 1357 5171 1363
rect 3773 1337 3811 1343
rect 3828 1337 3852 1343
rect 3885 1337 3923 1343
rect 4605 1337 4627 1343
rect 2580 1317 2595 1323
rect 4356 1317 4387 1323
rect 2397 1297 2451 1303
rect 3021 1297 3036 1303
rect 3156 1297 3171 1303
rect 445 1277 492 1283
rect 4461 1277 4515 1283
rect 5108 1277 5123 1283
rect 1380 1237 1411 1243
rect 2506 1236 2508 1244
rect 1242 1214 1254 1216
rect 4250 1214 4262 1216
rect 1227 1206 1229 1214
rect 1237 1206 1239 1214
rect 1247 1206 1249 1214
rect 1257 1206 1259 1214
rect 1267 1206 1269 1214
rect 4235 1206 4237 1214
rect 4245 1206 4247 1214
rect 4255 1206 4257 1214
rect 4265 1206 4267 1214
rect 4275 1206 4277 1214
rect 1242 1204 1254 1206
rect 4250 1204 4262 1206
rect 29 1137 60 1143
rect 52 1117 67 1123
rect 1684 1116 1692 1124
rect 349 1097 364 1103
rect 372 1097 403 1103
rect 1284 1097 1299 1103
rect 1453 1097 1484 1103
rect 1716 1097 1731 1103
rect 2260 1097 2291 1103
rect 2301 1097 2355 1103
rect 2532 1097 2563 1103
rect 2573 1097 2611 1103
rect 3149 1103 3155 1123
rect 4164 1116 4172 1124
rect 3117 1097 3155 1103
rect 3997 1097 4019 1103
rect 4109 1097 4124 1103
rect 4196 1097 4211 1103
rect 4365 1097 4380 1103
rect 4564 1097 4588 1103
rect 4605 1097 4636 1103
rect 4724 1097 4755 1103
rect 5037 1103 5043 1123
rect 5037 1097 5075 1103
rect 1556 1077 1571 1083
rect 1629 1077 1667 1083
rect 2164 1077 2179 1083
rect 2189 1077 2243 1083
rect 2317 1077 2332 1083
rect 3197 1077 3235 1083
rect 3805 1077 3827 1083
rect 3844 1077 3875 1083
rect 4676 1077 4691 1083
rect 4932 1077 4947 1083
rect 1213 1057 1292 1063
rect 1421 1057 1436 1063
rect 2148 1057 2163 1063
rect 2372 1057 2387 1063
rect 2653 1057 2668 1063
rect 3940 1057 3955 1063
rect 4509 1057 4540 1063
rect 100 1036 102 1044
rect 4708 1036 4710 1044
rect 2746 1014 2758 1016
rect 2731 1006 2733 1014
rect 2741 1006 2743 1014
rect 2751 1006 2753 1014
rect 2761 1006 2763 1014
rect 2771 1006 2773 1014
rect 2746 1004 2758 1006
rect 125 977 140 983
rect 4756 976 4758 984
rect 893 957 931 963
rect 1309 957 1372 963
rect 2260 956 2268 964
rect 2477 957 2492 963
rect 2612 957 2707 963
rect 3076 957 3091 963
rect 317 937 355 943
rect 861 937 876 943
rect 916 937 947 943
rect 1869 937 1907 943
rect 1940 937 1955 943
rect 2029 937 2051 943
rect 2109 937 2147 943
rect 2301 937 2316 943
rect 2452 937 2483 943
rect 4141 937 4179 943
rect 4701 937 4716 943
rect 4724 937 4755 943
rect 4781 937 4834 943
rect 29 917 67 923
rect 244 917 259 923
rect 269 917 300 923
rect 1485 917 1500 923
rect 1981 917 2019 923
rect 484 897 499 903
rect 1524 896 1532 904
rect 1981 897 1987 917
rect 2173 917 2211 923
rect 2132 897 2163 903
rect 2173 897 2179 917
rect 2372 917 2403 923
rect 2413 917 2460 923
rect 2484 917 2499 923
rect 3469 917 3507 923
rect 3469 897 3475 917
rect 3870 917 3900 923
rect 4061 917 4099 923
rect 3940 897 3955 903
rect 4093 897 4099 917
rect 4500 917 4515 923
rect 4564 917 4579 923
rect 781 877 796 883
rect 2221 877 2236 883
rect 3900 883 3908 888
rect 3892 877 3908 883
rect 4420 877 4435 883
rect 74 836 76 844
rect 4602 836 4604 844
rect 1242 814 1254 816
rect 4250 814 4262 816
rect 1227 806 1229 814
rect 1237 806 1239 814
rect 1247 806 1249 814
rect 1257 806 1259 814
rect 1267 806 1269 814
rect 4235 806 4237 814
rect 4245 806 4247 814
rect 4255 806 4257 814
rect 4265 806 4267 814
rect 4275 806 4277 814
rect 1242 804 1254 806
rect 4250 804 4262 806
rect 36 776 38 784
rect 154 776 156 784
rect 234 776 236 784
rect 4077 777 4108 783
rect 5018 776 5020 784
rect 404 717 419 723
rect 77 697 92 703
rect 132 697 147 703
rect 205 697 220 703
rect 573 703 579 723
rect 573 697 611 703
rect 780 703 788 708
rect 772 697 788 703
rect 892 703 900 708
rect 892 697 930 703
rect 2557 703 2563 723
rect 2557 697 2595 703
rect 2653 697 2732 703
rect 3133 703 3139 723
rect 3956 717 3971 723
rect 5092 717 5107 723
rect 3133 697 3171 703
rect 3837 697 3852 703
rect 4541 697 4556 703
rect 4653 697 4668 703
rect 4788 697 4803 703
rect 4861 697 4876 703
rect 4893 697 4924 703
rect 109 677 140 683
rect 308 677 339 683
rect 2493 677 2515 683
rect 3325 677 3347 683
rect 3853 677 3868 683
rect 4557 677 4579 683
rect 4596 677 4627 683
rect 4637 677 4652 683
rect 4701 677 4739 683
rect 4916 677 4931 683
rect 5085 677 5100 683
rect 5133 677 5148 683
rect 2676 657 2755 663
rect 3357 657 3395 663
rect 4826 656 4828 664
rect 5114 636 5116 644
rect 2746 614 2758 616
rect 2731 606 2733 614
rect 2741 606 2743 614
rect 2751 606 2753 614
rect 2761 606 2763 614
rect 2771 606 2773 614
rect 2746 604 2758 606
rect 356 576 358 584
rect 733 557 748 563
rect 1364 557 1379 563
rect 1437 557 1468 563
rect 2333 557 2348 563
rect 3565 557 3580 563
rect 4397 557 4435 563
rect 1492 537 1507 543
rect 1709 543 1715 556
rect 1709 537 1731 543
rect 2253 537 2291 543
rect 3613 537 3635 543
rect 4100 537 4115 543
rect 4973 537 4995 543
rect 1373 517 1411 523
rect 1492 517 1523 523
rect 1533 517 1571 523
rect 29 497 44 503
rect 77 497 115 503
rect 365 497 387 503
rect 1533 497 1539 517
rect 1636 517 1651 523
rect 1668 517 1683 523
rect 2173 517 2211 523
rect 2173 497 2179 517
rect 3518 517 3548 523
rect 3677 517 3715 523
rect 3677 497 3683 517
rect 4260 517 4307 523
rect 4900 517 4915 523
rect 4989 523 4995 537
rect 4989 517 5027 523
rect 5117 497 5132 503
rect 2093 477 2108 483
rect 2253 477 2268 483
rect 276 436 278 444
rect 1418 436 1420 444
rect 2733 437 2796 443
rect 1242 414 1254 416
rect 4250 414 4262 416
rect 1227 406 1229 414
rect 1237 406 1239 414
rect 1247 406 1249 414
rect 1257 406 1259 414
rect 1267 406 1269 414
rect 4235 406 4237 414
rect 4245 406 4247 414
rect 4255 406 4257 414
rect 4265 406 4267 414
rect 4275 406 4277 414
rect 1242 404 1254 406
rect 4250 404 4262 406
rect 2260 376 2262 384
rect 4093 377 4140 383
rect 2148 337 2163 343
rect 2061 303 2067 323
rect 2196 316 2204 324
rect 2285 317 2300 323
rect 2605 317 2620 323
rect 2061 297 2099 303
rect 2116 297 2140 303
rect 2157 297 2195 303
rect 2228 297 2259 303
rect 2733 303 2739 323
rect 2733 297 2835 303
rect 2845 297 2876 303
rect 5252 297 5267 303
rect 2669 277 2691 283
rect 4733 277 4755 283
rect 4556 263 4564 272
rect 4556 257 4588 263
rect 1741 237 1756 243
rect 2746 214 2758 216
rect 2731 206 2733 214
rect 2741 206 2743 214
rect 2751 206 2753 214
rect 2761 206 2763 214
rect 2771 206 2773 214
rect 2746 204 2758 206
rect 2356 176 2358 184
rect 2141 157 2179 163
rect 765 137 780 143
rect 2180 137 2211 143
rect 2749 137 2780 143
rect 2804 137 2835 143
rect 708 117 723 123
rect 1229 117 1331 123
rect 1341 117 1394 123
rect 1764 117 1779 123
rect 2260 117 2291 123
rect 2477 117 2515 123
rect 2509 97 2515 117
rect 2564 117 2595 123
rect 2605 117 2620 123
rect 2749 117 2812 123
rect 2749 104 2755 117
rect 2820 117 2851 123
rect 3757 117 3780 123
rect 3772 114 3780 117
rect 4556 117 4579 123
rect 4556 114 4564 117
rect 5374 117 5411 123
rect 2660 97 2691 103
rect 3197 97 3212 103
rect 2292 76 2294 84
rect 2404 76 2406 84
rect 2538 76 2540 84
rect 5485 77 5516 83
rect 1242 14 1254 16
rect 4250 14 4262 16
rect 1227 6 1229 14
rect 1237 6 1239 14
rect 1247 6 1249 14
rect 1257 6 1259 14
rect 1267 6 1269 14
rect 4235 6 4237 14
rect 4245 6 4247 14
rect 4255 6 4257 14
rect 4265 6 4267 14
rect 4275 6 4277 14
rect 1242 4 1254 6
rect 4250 4 4262 6
<< m2contact >>
rect 2723 3806 2731 3814
rect 2733 3806 2741 3814
rect 2743 3806 2751 3814
rect 2753 3806 2761 3814
rect 2763 3806 2771 3814
rect 2773 3806 2781 3814
rect 2188 3776 2196 3784
rect 3420 3776 3428 3784
rect 3884 3776 3892 3784
rect 188 3756 196 3764
rect 524 3756 532 3764
rect 892 3756 900 3764
rect 1308 3756 1316 3764
rect 1644 3756 1652 3764
rect 1996 3756 2004 3764
rect 2492 3756 2500 3764
rect 2700 3756 2708 3764
rect 3020 3756 3028 3764
rect 3148 3756 3156 3764
rect 3644 3756 3652 3764
rect 4108 3756 4116 3764
rect 4540 3756 4548 3764
rect 4876 3756 4884 3764
rect 5292 3756 5300 3764
rect 5484 3756 5492 3764
rect 220 3736 228 3744
rect 492 3736 500 3744
rect 924 3736 932 3744
rect 1340 3736 1348 3744
rect 1612 3736 1620 3744
rect 1964 3736 1972 3744
rect 2284 3736 2292 3744
rect 2348 3736 2356 3744
rect 2364 3736 2372 3744
rect 2396 3736 2404 3744
rect 2428 3736 2436 3744
rect 2460 3736 2468 3744
rect 2476 3736 2484 3744
rect 2732 3736 2740 3744
rect 2956 3736 2964 3744
rect 2988 3736 2996 3744
rect 3004 3736 3012 3744
rect 3068 3736 3076 3744
rect 3196 3736 3204 3744
rect 3356 3736 3364 3744
rect 3372 3736 3380 3744
rect 3404 3736 3412 3744
rect 3468 3736 3476 3744
rect 3612 3736 3620 3744
rect 3932 3736 3940 3744
rect 4076 3736 4084 3744
rect 4270 3736 4278 3744
rect 4572 3736 4580 3744
rect 4844 3736 4852 3744
rect 5068 3736 5076 3744
rect 5324 3736 5332 3744
rect 284 3716 292 3724
rect 316 3716 324 3724
rect 380 3716 388 3724
rect 604 3716 612 3724
rect 1004 3716 1012 3724
rect 1404 3716 1412 3724
rect 1532 3716 1540 3724
rect 1724 3716 1732 3724
rect 1868 3716 1876 3724
rect 2268 3716 2276 3724
rect 2332 3716 2340 3724
rect 2444 3716 2452 3724
rect 2812 3716 2820 3724
rect 2972 3716 2980 3724
rect 3100 3716 3108 3724
rect 3148 3716 3156 3724
rect 3180 3716 3188 3724
rect 3196 3716 3204 3724
rect 3228 3716 3236 3724
rect 3276 3716 3284 3724
rect 3452 3716 3460 3724
rect 3724 3716 3732 3724
rect 3820 3716 3828 3724
rect 3868 3716 3876 3724
rect 3916 3716 3924 3724
rect 3996 3716 4004 3724
rect 4378 3716 4386 3724
rect 4636 3716 4644 3724
rect 4748 3716 4756 3724
rect 4956 3716 4964 3724
rect 5212 3716 5220 3724
rect 5420 3716 5428 3724
rect 316 3696 324 3704
rect 428 3700 436 3708
rect 988 3700 996 3708
rect 1436 3696 1444 3704
rect 1548 3700 1556 3708
rect 1900 3700 1908 3708
rect 2156 3696 2164 3704
rect 2188 3696 2196 3704
rect 2220 3696 2228 3704
rect 2364 3696 2372 3704
rect 2508 3696 2516 3704
rect 2828 3696 2836 3704
rect 3036 3696 3044 3704
rect 3084 3696 3092 3704
rect 3260 3696 3268 3704
rect 3324 3696 3332 3704
rect 3340 3696 3348 3704
rect 3372 3696 3380 3704
rect 3516 3696 3524 3704
rect 3884 3696 3892 3704
rect 3980 3696 3988 3704
rect 4668 3696 4676 3704
rect 4780 3700 4788 3708
rect 5100 3696 5108 3704
rect 5388 3700 5396 3708
rect 12 3676 20 3684
rect 732 3676 740 3684
rect 1820 3676 1828 3684
rect 2300 3676 2308 3684
rect 2332 3676 2340 3684
rect 2396 3676 2404 3684
rect 2924 3676 2932 3684
rect 3100 3676 3108 3684
rect 3132 3676 3140 3684
rect 3292 3676 3300 3684
rect 5068 3676 5076 3684
rect 988 3654 996 3662
rect 1148 3656 1156 3664
rect 3276 3656 3284 3664
rect 3724 3654 3732 3662
rect 4780 3654 4788 3662
rect 316 3636 324 3644
rect 428 3636 436 3644
rect 684 3636 692 3644
rect 1436 3636 1444 3644
rect 1548 3636 1556 3644
rect 1900 3636 1908 3644
rect 2540 3636 2548 3644
rect 2828 3636 2836 3644
rect 3052 3636 3060 3644
rect 3804 3636 3812 3644
rect 3980 3636 3988 3644
rect 4668 3636 4676 3644
rect 5036 3636 5044 3644
rect 5132 3636 5140 3644
rect 5388 3636 5396 3644
rect 5468 3636 5476 3644
rect 1219 3606 1227 3614
rect 1229 3606 1237 3614
rect 1239 3606 1247 3614
rect 1249 3606 1257 3614
rect 1259 3606 1267 3614
rect 1269 3606 1277 3614
rect 4227 3606 4235 3614
rect 4237 3606 4245 3614
rect 4247 3606 4255 3614
rect 4257 3606 4265 3614
rect 4267 3606 4275 3614
rect 4277 3606 4285 3614
rect 316 3576 324 3584
rect 1436 3576 1444 3584
rect 2460 3576 2468 3584
rect 2524 3576 2532 3584
rect 2684 3576 2692 3584
rect 3036 3576 3044 3584
rect 3116 3576 3124 3584
rect 3196 3576 3204 3584
rect 3260 3576 3268 3584
rect 3612 3576 3620 3584
rect 3692 3576 3700 3584
rect 3884 3576 3892 3584
rect 4060 3576 4068 3584
rect 4460 3576 4468 3584
rect 4572 3576 4580 3584
rect 4796 3576 4804 3584
rect 5052 3576 5060 3584
rect 5084 3576 5092 3584
rect 5452 3576 5460 3584
rect 652 3558 660 3566
rect 1052 3558 1060 3566
rect 2028 3558 2036 3566
rect 2380 3558 2388 3566
rect 3788 3556 3796 3564
rect 4732 3556 4740 3564
rect 4924 3556 4932 3564
rect 4988 3556 4996 3564
rect 2476 3536 2484 3544
rect 2540 3536 2548 3544
rect 3020 3536 3028 3544
rect 3244 3536 3252 3544
rect 3372 3536 3380 3544
rect 3388 3536 3396 3544
rect 3756 3536 3764 3544
rect 4204 3536 4212 3544
rect 4444 3536 4452 3544
rect 4492 3536 4500 3544
rect 4940 3536 4948 3544
rect 5004 3536 5012 3544
rect 316 3516 324 3524
rect 572 3516 580 3524
rect 652 3512 660 3520
rect 1052 3512 1060 3520
rect 1436 3516 1444 3524
rect 2028 3512 2036 3520
rect 2380 3512 2388 3520
rect 2508 3516 2516 3524
rect 2572 3516 2580 3524
rect 2684 3516 2692 3524
rect 3052 3516 3060 3524
rect 3212 3516 3220 3524
rect 3276 3516 3284 3524
rect 3404 3516 3412 3524
rect 3564 3516 3572 3524
rect 284 3496 292 3504
rect 316 3496 324 3504
rect 444 3496 452 3504
rect 604 3496 612 3504
rect 828 3496 836 3504
rect 924 3496 932 3504
rect 1004 3496 1012 3504
rect 1228 3496 1236 3504
rect 1436 3496 1444 3504
rect 1532 3496 1540 3504
rect 2060 3496 2068 3504
rect 2204 3496 2212 3504
rect 2428 3496 2436 3504
rect 2492 3496 2500 3504
rect 2556 3496 2564 3504
rect 2684 3496 2692 3504
rect 2700 3496 2708 3504
rect 2974 3496 2982 3504
rect 3036 3496 3044 3504
rect 3068 3496 3076 3504
rect 3100 3496 3108 3504
rect 3148 3496 3156 3504
rect 3260 3496 3268 3504
rect 3308 3496 3316 3504
rect 3340 3496 3348 3504
rect 3388 3496 3396 3504
rect 3420 3496 3428 3504
rect 3468 3496 3476 3504
rect 3532 3496 3540 3504
rect 3724 3516 3732 3524
rect 4348 3516 4356 3524
rect 4396 3516 4404 3524
rect 4412 3516 4420 3524
rect 4524 3516 4532 3524
rect 4620 3516 4628 3524
rect 4652 3516 4660 3524
rect 4764 3516 4772 3524
rect 4828 3516 4836 3524
rect 4972 3516 4980 3524
rect 5452 3516 5460 3524
rect 3612 3496 3620 3504
rect 3660 3496 3668 3504
rect 3692 3496 3700 3504
rect 3756 3496 3764 3504
rect 3836 3496 3844 3504
rect 3932 3496 3940 3504
rect 3948 3496 3956 3504
rect 3980 3496 3988 3504
rect 4012 3496 4020 3504
rect 4124 3496 4132 3504
rect 4204 3496 4212 3504
rect 4364 3496 4372 3504
rect 4428 3496 4436 3504
rect 4492 3496 4500 3504
rect 4556 3496 4564 3504
rect 4588 3496 4596 3504
rect 4620 3496 4628 3504
rect 4652 3496 4660 3504
rect 4732 3496 4740 3504
rect 4796 3496 4804 3504
rect 4924 3496 4932 3504
rect 4988 3496 4996 3504
rect 5036 3496 5044 3504
rect 5132 3496 5140 3504
rect 5420 3496 5428 3504
rect 220 3476 228 3484
rect 540 3476 548 3484
rect 716 3476 724 3484
rect 1116 3476 1124 3484
rect 1532 3476 1540 3484
rect 1964 3476 1972 3484
rect 2316 3476 2324 3484
rect 2780 3476 2788 3484
rect 3180 3476 3188 3484
rect 3324 3476 3332 3484
rect 3372 3476 3380 3484
rect 3452 3476 3460 3484
rect 188 3456 196 3464
rect 380 3456 388 3464
rect 428 3456 436 3464
rect 476 3456 484 3464
rect 492 3456 500 3464
rect 524 3456 532 3464
rect 748 3456 756 3464
rect 940 3456 948 3464
rect 972 3456 980 3464
rect 1148 3456 1156 3464
rect 1564 3456 1572 3464
rect 1932 3456 1940 3464
rect 2284 3456 2292 3464
rect 2812 3456 2820 3464
rect 3100 3456 3108 3464
rect 3292 3456 3300 3464
rect 3452 3456 3460 3464
rect 3516 3476 3524 3484
rect 3628 3476 3636 3484
rect 3644 3476 3652 3484
rect 3708 3476 3716 3484
rect 3772 3476 3780 3484
rect 3820 3476 3828 3484
rect 3868 3476 3876 3484
rect 3916 3476 3924 3484
rect 3964 3476 3972 3484
rect 4028 3476 4036 3484
rect 4108 3476 4116 3484
rect 4364 3476 4372 3484
rect 4476 3476 4484 3484
rect 4540 3476 4548 3484
rect 4604 3476 4612 3484
rect 4668 3476 4676 3484
rect 4716 3476 4724 3484
rect 4780 3476 4788 3484
rect 5116 3476 5124 3484
rect 5356 3476 5364 3484
rect 3788 3456 3796 3464
rect 3852 3456 3860 3464
rect 3884 3456 3892 3464
rect 3996 3456 4004 3464
rect 4076 3456 4084 3464
rect 4092 3456 4100 3464
rect 4236 3456 4244 3464
rect 4684 3456 4692 3464
rect 4700 3456 4708 3464
rect 4844 3456 4852 3464
rect 4876 3456 4884 3464
rect 5068 3456 5076 3464
rect 5084 3456 5092 3464
rect 5324 3456 5332 3464
rect 28 3436 36 3444
rect 412 3436 420 3444
rect 460 3436 468 3444
rect 956 3436 964 3444
rect 1308 3436 1316 3444
rect 1724 3436 1732 3444
rect 1772 3436 1780 3444
rect 2124 3436 2132 3444
rect 4108 3436 4116 3444
rect 4396 3436 4404 3444
rect 4860 3436 4868 3444
rect 5164 3436 5172 3444
rect 2723 3406 2731 3414
rect 2733 3406 2741 3414
rect 2743 3406 2751 3414
rect 2753 3406 2761 3414
rect 2763 3406 2771 3414
rect 2773 3406 2781 3414
rect 444 3376 452 3384
rect 1756 3376 1764 3384
rect 1996 3376 2004 3384
rect 2092 3376 2100 3384
rect 2652 3376 2660 3384
rect 3516 3376 3524 3384
rect 3820 3376 3828 3384
rect 3884 3376 3892 3384
rect 3948 3376 3956 3384
rect 4124 3376 4132 3384
rect 4284 3376 4292 3384
rect 4508 3376 4516 3384
rect 5228 3376 5236 3384
rect 5340 3376 5348 3384
rect 12 3356 20 3364
rect 220 3356 228 3364
rect 748 3356 756 3364
rect 796 3356 804 3364
rect 924 3356 932 3364
rect 1116 3356 1124 3364
rect 1516 3356 1524 3364
rect 1820 3356 1828 3364
rect 1916 3356 1924 3364
rect 2140 3356 2148 3364
rect 2364 3356 2372 3364
rect 2908 3356 2916 3364
rect 3260 3356 3268 3364
rect 3564 3356 3572 3364
rect 3740 3356 3748 3364
rect 4188 3356 4196 3364
rect 4236 3356 4244 3364
rect 4572 3356 4580 3364
rect 4748 3356 4756 3364
rect 5068 3356 5076 3364
rect 5212 3356 5220 3364
rect 5244 3356 5252 3364
rect 5436 3356 5444 3364
rect 252 3336 260 3344
rect 396 3336 404 3344
rect 492 3336 500 3344
rect 636 3336 644 3344
rect 732 3336 740 3344
rect 1148 3336 1156 3344
rect 1484 3336 1492 3344
rect 1692 3336 1700 3344
rect 1932 3336 1940 3344
rect 2012 3336 2020 3344
rect 2124 3336 2132 3344
rect 2396 3336 2404 3344
rect 2540 3336 2548 3344
rect 2876 3336 2884 3344
rect 3228 3336 3236 3344
rect 3436 3336 3444 3344
rect 3484 3336 3492 3344
rect 3548 3336 3556 3344
rect 3644 3336 3652 3344
rect 3740 3336 3748 3344
rect 3804 3336 3812 3344
rect 3932 3336 3940 3344
rect 3980 3336 3988 3344
rect 4028 3336 4036 3344
rect 4092 3336 4100 3344
rect 4172 3336 4180 3344
rect 4492 3336 4500 3344
rect 316 3316 324 3324
rect 348 3296 356 3304
rect 428 3296 436 3304
rect 476 3316 484 3324
rect 524 3316 532 3324
rect 588 3316 596 3324
rect 636 3316 644 3324
rect 668 3316 676 3324
rect 828 3316 836 3324
rect 876 3316 884 3324
rect 908 3316 916 3324
rect 1228 3316 1236 3324
rect 1404 3316 1412 3324
rect 1596 3316 1604 3324
rect 1740 3316 1748 3324
rect 1804 3316 1812 3324
rect 1868 3316 1876 3324
rect 1964 3316 1972 3324
rect 2060 3316 2068 3324
rect 2284 3316 2292 3324
rect 2812 3316 2820 3324
rect 3116 3316 3124 3324
rect 3148 3316 3156 3324
rect 3532 3316 3540 3324
rect 3628 3316 3636 3324
rect 3708 3316 3716 3324
rect 3916 3316 3924 3324
rect 4076 3316 4084 3324
rect 4716 3336 4724 3344
rect 5036 3336 5044 3344
rect 5084 3336 5092 3344
rect 5148 3336 5156 3344
rect 5356 3336 5364 3344
rect 4140 3316 4148 3324
rect 4300 3316 4308 3324
rect 4396 3316 4404 3324
rect 4460 3316 4468 3324
rect 4476 3316 4484 3324
rect 4524 3316 4532 3324
rect 4556 3316 4564 3324
rect 4636 3316 4644 3324
rect 4652 3316 4660 3324
rect 4972 3316 4980 3324
rect 5020 3316 5028 3324
rect 5100 3316 5108 3324
rect 5148 3316 5156 3324
rect 5164 3316 5172 3324
rect 5180 3316 5188 3324
rect 5212 3316 5220 3324
rect 5308 3316 5316 3324
rect 5372 3316 5380 3324
rect 5484 3316 5492 3324
rect 508 3296 516 3304
rect 572 3296 580 3304
rect 636 3296 644 3304
rect 700 3296 708 3304
rect 748 3296 756 3304
rect 892 3296 900 3304
rect 1212 3300 1220 3308
rect 1420 3300 1428 3308
rect 1756 3296 1764 3304
rect 1996 3296 2004 3304
rect 2044 3296 2052 3304
rect 2460 3300 2468 3308
rect 2780 3296 2788 3304
rect 3164 3300 3172 3308
rect 3516 3296 3524 3304
rect 3596 3296 3604 3304
rect 3660 3296 3668 3304
rect 3756 3296 3764 3304
rect 3836 3296 3844 3304
rect 3884 3296 3892 3304
rect 3948 3296 3956 3304
rect 3980 3296 3988 3304
rect 4380 3296 4388 3304
rect 4444 3296 4452 3304
rect 4620 3296 4628 3304
rect 4940 3296 4948 3304
rect 4972 3296 4980 3304
rect 5132 3296 5140 3304
rect 5196 3296 5204 3304
rect 5340 3296 5348 3304
rect 5372 3296 5380 3304
rect 44 3276 52 3284
rect 540 3276 548 3284
rect 604 3276 612 3284
rect 860 3276 868 3284
rect 1884 3276 1892 3284
rect 3436 3276 3444 3284
rect 4412 3276 4420 3284
rect 5404 3276 5412 3284
rect 5452 3276 5460 3284
rect 524 3256 532 3264
rect 1212 3254 1220 3262
rect 2460 3254 2468 3262
rect 3164 3254 3172 3262
rect 4012 3256 4020 3264
rect 4076 3256 4084 3264
rect 28 3236 36 3244
rect 348 3236 356 3244
rect 876 3236 884 3244
rect 956 3236 964 3244
rect 1420 3236 1428 3244
rect 1676 3236 1684 3244
rect 1868 3236 1876 3244
rect 2028 3236 2036 3244
rect 2108 3236 2116 3244
rect 2204 3236 2212 3244
rect 2780 3236 2788 3244
rect 3068 3236 3076 3244
rect 3468 3236 3476 3244
rect 3692 3236 3700 3244
rect 3868 3236 3876 3244
rect 4396 3236 4404 3244
rect 4620 3236 4628 3244
rect 4908 3236 4916 3244
rect 5052 3236 5060 3244
rect 1219 3206 1227 3214
rect 1229 3206 1237 3214
rect 1239 3206 1247 3214
rect 1249 3206 1257 3214
rect 1259 3206 1267 3214
rect 1269 3206 1277 3214
rect 4227 3206 4235 3214
rect 4237 3206 4245 3214
rect 4247 3206 4255 3214
rect 4257 3206 4265 3214
rect 4267 3206 4275 3214
rect 4277 3206 4285 3214
rect 300 3176 308 3184
rect 444 3176 452 3184
rect 572 3176 580 3184
rect 636 3176 644 3184
rect 684 3176 692 3184
rect 1404 3176 1412 3184
rect 1564 3176 1572 3184
rect 1948 3176 1956 3184
rect 2444 3176 2452 3184
rect 2796 3176 2804 3184
rect 3308 3176 3316 3184
rect 3420 3176 3428 3184
rect 3596 3176 3604 3184
rect 3692 3176 3700 3184
rect 3996 3176 4004 3184
rect 4076 3176 4084 3184
rect 4444 3176 4452 3184
rect 4732 3176 4740 3184
rect 4780 3176 4788 3184
rect 4956 3176 4964 3184
rect 4988 3176 4996 3184
rect 5244 3176 5252 3184
rect 524 3156 532 3164
rect 3116 3156 3124 3164
rect 92 3136 100 3144
rect 124 3136 132 3144
rect 172 3136 180 3144
rect 236 3136 244 3144
rect 412 3136 420 3144
rect 1052 3136 1060 3144
rect 1340 3136 1348 3144
rect 3324 3136 3332 3144
rect 3356 3136 3364 3144
rect 3612 3136 3620 3144
rect 4012 3136 4020 3144
rect 4060 3136 4068 3144
rect 4076 3136 4084 3144
rect 60 3116 68 3124
rect 220 3116 228 3124
rect 252 3116 260 3124
rect 268 3116 276 3124
rect 540 3116 548 3124
rect 556 3116 564 3124
rect 652 3116 660 3124
rect 940 3116 948 3124
rect 12 3096 20 3104
rect 76 3096 84 3104
rect 188 3096 196 3104
rect 300 3096 308 3104
rect 364 3096 372 3104
rect 412 3096 420 3104
rect 444 3096 452 3104
rect 476 3096 484 3104
rect 572 3096 580 3104
rect 668 3096 676 3104
rect 716 3096 724 3104
rect 924 3096 932 3104
rect 988 3116 996 3124
rect 1100 3116 1108 3124
rect 1372 3116 1380 3124
rect 1436 3116 1444 3124
rect 1660 3116 1668 3124
rect 1724 3116 1732 3124
rect 1148 3096 1156 3104
rect 1212 3096 1220 3104
rect 1356 3096 1364 3104
rect 220 3076 228 3084
rect 316 3076 324 3084
rect 428 3076 436 3084
rect 492 3076 500 3084
rect 508 3076 516 3084
rect 620 3076 628 3084
rect 668 3076 676 3084
rect 732 3076 740 3084
rect 780 3076 788 3084
rect 908 3076 916 3084
rect 924 3076 932 3084
rect 1020 3076 1028 3084
rect 1036 3076 1044 3084
rect 1196 3076 1204 3084
rect 1404 3096 1412 3104
rect 1596 3096 1604 3104
rect 1644 3096 1652 3104
rect 1676 3096 1684 3104
rect 1692 3096 1700 3104
rect 1708 3096 1716 3104
rect 1756 3096 1764 3104
rect 1916 3116 1924 3124
rect 1900 3096 1908 3104
rect 1948 3096 1956 3104
rect 2060 3116 2068 3124
rect 2172 3116 2180 3124
rect 2188 3116 2196 3124
rect 2220 3116 2228 3124
rect 2284 3116 2292 3124
rect 2332 3116 2340 3124
rect 2476 3116 2484 3124
rect 2796 3116 2804 3124
rect 3180 3112 3188 3120
rect 3484 3116 3492 3124
rect 2092 3096 2100 3104
rect 2140 3096 2148 3104
rect 2364 3096 2372 3104
rect 2444 3096 2452 3104
rect 2700 3096 2708 3104
rect 2812 3096 2820 3104
rect 3116 3096 3124 3104
rect 3260 3096 3268 3104
rect 3356 3096 3364 3104
rect 3452 3096 3460 3104
rect 3484 3096 3492 3104
rect 3532 3116 3540 3124
rect 3580 3116 3588 3124
rect 3756 3116 3764 3124
rect 3916 3116 3924 3124
rect 3980 3116 3988 3124
rect 4092 3116 4100 3124
rect 4364 3116 4372 3124
rect 4444 3116 4452 3124
rect 5148 3116 5156 3124
rect 5340 3116 5348 3124
rect 5372 3116 5380 3124
rect 5404 3116 5412 3124
rect 5420 3116 5428 3124
rect 3596 3096 3604 3104
rect 3756 3096 3764 3104
rect 3788 3096 3796 3104
rect 3836 3096 3844 3104
rect 3868 3096 3876 3104
rect 3948 3096 3956 3104
rect 3996 3096 4004 3104
rect 4076 3096 4084 3104
rect 4140 3096 4148 3104
rect 4300 3096 4308 3104
rect 4332 3096 4340 3104
rect 4444 3096 4452 3104
rect 4652 3096 4660 3104
rect 5036 3096 5044 3104
rect 5100 3096 5108 3104
rect 5116 3096 5124 3104
rect 5196 3096 5204 3104
rect 5308 3096 5316 3104
rect 5372 3096 5380 3104
rect 1452 3076 1460 3084
rect 1612 3076 1620 3084
rect 1708 3076 1716 3084
rect 1964 3076 1972 3084
rect 1996 3076 2004 3084
rect 2108 3076 2116 3084
rect 2124 3076 2132 3084
rect 2268 3076 2276 3084
rect 2380 3076 2388 3084
rect 12 3056 20 3064
rect 44 3056 52 3064
rect 140 3056 148 3064
rect 332 3056 340 3064
rect 348 3056 356 3064
rect 380 3056 388 3064
rect 748 3056 756 3064
rect 764 3056 772 3064
rect 1084 3056 1092 3064
rect 1116 3056 1124 3064
rect 1180 3056 1188 3064
rect 1644 3056 1652 3064
rect 1788 3056 1796 3064
rect 1868 3056 1876 3064
rect 1996 3056 2004 3064
rect 2700 3076 2708 3084
rect 3116 3076 3124 3084
rect 3276 3076 3284 3084
rect 3372 3076 3380 3084
rect 3404 3076 3412 3084
rect 3468 3076 3476 3084
rect 3564 3076 3572 3084
rect 3692 3076 3700 3084
rect 3724 3076 3732 3084
rect 3788 3076 3796 3084
rect 3820 3076 3828 3084
rect 3852 3076 3860 3084
rect 3900 3076 3908 3084
rect 3964 3076 3972 3084
rect 4124 3076 4132 3084
rect 4540 3076 4548 3084
rect 4924 3076 4932 3084
rect 5084 3076 5092 3084
rect 5212 3076 5220 3084
rect 5292 3076 5300 3084
rect 5356 3076 5364 3084
rect 5516 3076 5524 3084
rect 2668 3056 2676 3064
rect 3084 3056 3092 3064
rect 3308 3056 3316 3064
rect 3404 3056 3412 3064
rect 3644 3056 3652 3064
rect 3756 3056 3764 3064
rect 3900 3056 3908 3064
rect 4140 3056 4148 3064
rect 4172 3056 4180 3064
rect 4188 3056 4196 3064
rect 4284 3056 4292 3064
rect 4396 3056 4404 3064
rect 4572 3056 4580 3064
rect 4940 3056 4948 3064
rect 5068 3056 5076 3064
rect 5164 3056 5172 3064
rect 5244 3056 5252 3064
rect 5260 3056 5268 3064
rect 108 3036 116 3044
rect 188 3036 196 3044
rect 572 3036 580 3044
rect 1260 3036 1268 3044
rect 1356 3036 1364 3044
rect 1836 3036 1844 3044
rect 2028 3036 2036 3044
rect 2172 3036 2180 3044
rect 2188 3036 2196 3044
rect 2284 3036 2292 3044
rect 2508 3036 2516 3044
rect 2924 3036 2932 3044
rect 4812 3036 4820 3044
rect 5148 3036 5156 3044
rect 5340 3036 5348 3044
rect 5436 3036 5444 3044
rect 2723 3006 2731 3014
rect 2733 3006 2741 3014
rect 2743 3006 2751 3014
rect 2753 3006 2761 3014
rect 2763 3006 2771 3014
rect 2773 3006 2781 3014
rect 284 2976 292 2984
rect 396 2976 404 2984
rect 1628 2976 1636 2984
rect 1660 2976 1668 2984
rect 1772 2976 1780 2984
rect 2012 2976 2020 2984
rect 2204 2976 2212 2984
rect 2300 2976 2308 2984
rect 2380 2976 2388 2984
rect 2556 2976 2564 2984
rect 2700 2976 2708 2984
rect 3276 2976 3284 2984
rect 3628 2976 3636 2984
rect 3708 2976 3716 2984
rect 3740 2976 3748 2984
rect 4060 2976 4068 2984
rect 4108 2976 4116 2984
rect 4300 2976 4308 2984
rect 4380 2976 4388 2984
rect 4876 2976 4884 2984
rect 5004 2976 5012 2984
rect 5100 2976 5108 2984
rect 108 2956 116 2964
rect 124 2956 132 2964
rect 140 2956 148 2964
rect 188 2956 196 2964
rect 204 2956 212 2964
rect 332 2956 340 2964
rect 556 2956 564 2964
rect 908 2956 916 2964
rect 1084 2956 1092 2964
rect 1196 2956 1204 2964
rect 1372 2956 1380 2964
rect 1564 2956 1572 2964
rect 1692 2956 1700 2964
rect 1980 2956 1988 2964
rect 2124 2956 2132 2964
rect 2492 2956 2500 2964
rect 2572 2956 2580 2964
rect 2588 2956 2596 2964
rect 2924 2956 2932 2964
rect 3308 2956 3316 2964
rect 3548 2956 3556 2964
rect 3612 2956 3620 2964
rect 3660 2956 3668 2964
rect 3756 2956 3764 2964
rect 3836 2956 3844 2964
rect 4092 2956 4100 2964
rect 4156 2956 4164 2964
rect 4188 2956 4196 2964
rect 332 2936 340 2944
rect 588 2936 596 2944
rect 940 2936 948 2944
rect 1180 2936 1188 2944
rect 1292 2936 1300 2944
rect 1436 2936 1444 2944
rect 1580 2936 1588 2944
rect 1644 2936 1652 2944
rect 1756 2936 1764 2944
rect 1804 2936 1812 2944
rect 1916 2936 1924 2944
rect 1964 2936 1972 2944
rect 2012 2936 2020 2944
rect 2044 2936 2052 2944
rect 2140 2936 2148 2944
rect 2172 2936 2180 2944
rect 2204 2936 2212 2944
rect 2236 2936 2244 2944
rect 2284 2936 2292 2944
rect 2316 2936 2324 2944
rect 2364 2936 2372 2944
rect 2396 2936 2404 2944
rect 2428 2936 2436 2944
rect 2540 2936 2548 2944
rect 2956 2936 2964 2944
rect 3228 2936 3236 2944
rect 3372 2936 3380 2944
rect 3516 2936 3524 2944
rect 3532 2936 3540 2944
rect 3676 2936 3684 2944
rect 3724 2936 3732 2944
rect 3772 2936 3780 2944
rect 3820 2936 3828 2944
rect 3916 2936 3924 2944
rect 3932 2936 3940 2944
rect 3996 2936 4004 2944
rect 4028 2936 4036 2944
rect 4364 2936 4372 2944
rect 4460 2936 4468 2944
rect 4684 2956 4692 2964
rect 4860 2956 4868 2964
rect 5036 2956 5044 2964
rect 5132 2956 5140 2964
rect 5308 2956 5316 2964
rect 4492 2936 4500 2944
rect 4716 2936 4724 2944
rect 4892 2936 4900 2944
rect 4924 2936 4932 2944
rect 4988 2936 4996 2944
rect 5020 2936 5028 2944
rect 5116 2936 5124 2944
rect 5340 2936 5348 2944
rect 44 2916 52 2924
rect 140 2916 148 2924
rect 236 2916 244 2924
rect 364 2916 372 2924
rect 476 2916 484 2924
rect 684 2916 692 2924
rect 828 2916 836 2924
rect 1036 2916 1044 2924
rect 1164 2916 1172 2924
rect 1228 2916 1236 2924
rect 1260 2916 1268 2924
rect 1372 2916 1380 2924
rect 1420 2916 1428 2924
rect 1500 2916 1508 2924
rect 1532 2916 1540 2924
rect 1548 2916 1556 2924
rect 1596 2916 1604 2924
rect 1676 2916 1684 2924
rect 1724 2916 1732 2924
rect 1740 2916 1748 2924
rect 1900 2916 1908 2924
rect 1996 2916 2004 2924
rect 2060 2916 2068 2924
rect 2252 2916 2260 2924
rect 2268 2916 2276 2924
rect 2332 2916 2340 2924
rect 2348 2916 2356 2924
rect 2412 2916 2420 2924
rect 2444 2916 2452 2924
rect 2492 2916 2500 2924
rect 2636 2916 2644 2924
rect 3052 2916 3060 2924
rect 3100 2916 3108 2924
rect 3276 2916 3284 2924
rect 3356 2916 3364 2924
rect 60 2896 68 2904
rect 220 2896 228 2904
rect 284 2896 292 2904
rect 652 2900 660 2908
rect 1004 2900 1012 2908
rect 1084 2896 1092 2904
rect 1132 2896 1140 2904
rect 1356 2896 1364 2904
rect 1452 2896 1460 2904
rect 1516 2896 1524 2904
rect 1628 2896 1636 2904
rect 1676 2896 1684 2904
rect 1820 2896 1828 2904
rect 1852 2896 1860 2904
rect 2076 2896 2084 2904
rect 2140 2896 2148 2904
rect 2668 2896 2676 2904
rect 3020 2900 3028 2908
rect 3292 2896 3300 2904
rect 3436 2916 3444 2924
rect 3468 2916 3476 2924
rect 3564 2916 3572 2924
rect 3692 2916 3700 2924
rect 3804 2916 3812 2924
rect 3836 2916 3844 2924
rect 3948 2916 3956 2924
rect 3964 2916 3972 2924
rect 4140 2916 4148 2924
rect 4188 2916 4196 2924
rect 4220 2916 4228 2924
rect 4332 2916 4340 2924
rect 4348 2916 4356 2924
rect 4412 2916 4420 2924
rect 4604 2916 4612 2924
rect 4796 2916 4804 2924
rect 4908 2916 4916 2924
rect 4940 2916 4948 2924
rect 4956 2916 4964 2924
rect 4988 2916 4996 2924
rect 5068 2916 5076 2924
rect 5228 2916 5236 2924
rect 3404 2896 3412 2904
rect 3772 2896 3780 2904
rect 3884 2896 3892 2904
rect 3980 2896 3988 2904
rect 3996 2896 4004 2904
rect 4076 2896 4084 2904
rect 4428 2896 4436 2904
rect 4780 2900 4788 2908
rect 5084 2896 5092 2904
rect 5404 2900 5412 2908
rect 188 2876 196 2884
rect 252 2876 260 2884
rect 1292 2876 1300 2884
rect 1484 2876 1492 2884
rect 3308 2876 3316 2884
rect 5068 2876 5076 2884
rect 652 2854 660 2862
rect 3020 2854 3028 2862
rect 4780 2854 4788 2862
rect 5404 2854 5412 2862
rect 44 2836 52 2844
rect 236 2836 244 2844
rect 364 2836 372 2844
rect 396 2836 404 2844
rect 748 2836 756 2844
rect 1004 2836 1012 2844
rect 1500 2836 1508 2844
rect 1932 2836 1940 2844
rect 2508 2836 2516 2844
rect 2764 2836 2772 2844
rect 4524 2836 4532 2844
rect 1219 2806 1227 2814
rect 1229 2806 1237 2814
rect 1239 2806 1247 2814
rect 1249 2806 1257 2814
rect 1259 2806 1267 2814
rect 1269 2806 1277 2814
rect 4227 2806 4235 2814
rect 4237 2806 4245 2814
rect 4247 2806 4255 2814
rect 4257 2806 4265 2814
rect 4267 2806 4275 2814
rect 4277 2806 4285 2814
rect 28 2776 36 2784
rect 316 2776 324 2784
rect 668 2776 676 2784
rect 1340 2776 1348 2784
rect 1740 2776 1748 2784
rect 1980 2776 1988 2784
rect 2076 2776 2084 2784
rect 2572 2776 2580 2784
rect 4540 2776 4548 2784
rect 4828 2776 4836 2784
rect 4892 2776 4900 2784
rect 5180 2776 5188 2784
rect 972 2758 980 2766
rect 2892 2756 2900 2764
rect 3164 2756 3172 2764
rect 3612 2756 3620 2764
rect 3900 2758 3908 2766
rect 380 2736 388 2744
rect 1676 2736 1684 2744
rect 1740 2736 1748 2744
rect 1756 2736 1764 2744
rect 1868 2736 1876 2744
rect 1996 2736 2004 2744
rect 2108 2736 2116 2744
rect 2380 2736 2388 2744
rect 3356 2736 3364 2744
rect 4172 2736 4180 2744
rect 316 2716 324 2724
rect 444 2716 452 2724
rect 604 2716 612 2724
rect 652 2716 660 2724
rect 700 2716 708 2724
rect 972 2712 980 2720
rect 1404 2716 1412 2724
rect 1452 2716 1460 2724
rect 1660 2716 1668 2724
rect 1708 2716 1716 2724
rect 1724 2716 1732 2724
rect 1788 2716 1796 2724
rect 1836 2716 1844 2724
rect 1900 2716 1908 2724
rect 1964 2716 1972 2724
rect 2204 2716 2212 2724
rect 2252 2716 2260 2724
rect 2348 2716 2356 2724
rect 2524 2716 2532 2724
rect 2956 2712 2964 2720
rect 3068 2716 3076 2724
rect 3548 2712 3556 2720
rect 3900 2712 3908 2720
rect 4380 2716 4388 2724
rect 4444 2716 4452 2724
rect 4828 2716 4836 2724
rect 5180 2716 5188 2724
rect 284 2696 292 2704
rect 300 2696 308 2704
rect 380 2696 388 2704
rect 412 2696 420 2704
rect 492 2696 500 2704
rect 524 2696 532 2704
rect 556 2696 564 2704
rect 732 2696 740 2704
rect 796 2696 804 2704
rect 828 2696 836 2704
rect 860 2696 868 2704
rect 1036 2696 1044 2704
rect 1148 2696 1156 2704
rect 1324 2696 1332 2704
rect 1388 2696 1396 2704
rect 1420 2696 1428 2704
rect 1484 2696 1492 2704
rect 1564 2696 1572 2704
rect 1612 2696 1620 2704
rect 1740 2696 1748 2704
rect 1884 2696 1892 2704
rect 1932 2696 1940 2704
rect 1980 2696 1988 2704
rect 2028 2696 2036 2704
rect 2092 2696 2100 2704
rect 2108 2696 2116 2704
rect 2140 2696 2148 2704
rect 2268 2696 2276 2704
rect 2316 2696 2324 2704
rect 2364 2696 2372 2704
rect 2428 2696 2436 2704
rect 2492 2696 2500 2704
rect 2556 2696 2564 2704
rect 2588 2696 2596 2704
rect 2892 2696 2900 2704
rect 3164 2696 3172 2704
rect 3436 2696 3444 2704
rect 3612 2696 3620 2704
rect 3868 2696 3876 2704
rect 4188 2696 4196 2704
rect 4348 2696 4356 2704
rect 4412 2696 4420 2704
rect 4428 2696 4436 2704
rect 4620 2696 4628 2704
rect 4796 2696 4804 2704
rect 4828 2696 4836 2704
rect 4972 2696 4980 2704
rect 5196 2696 5204 2704
rect 220 2676 228 2684
rect 364 2676 372 2684
rect 428 2676 436 2684
rect 476 2676 484 2684
rect 540 2676 548 2684
rect 636 2676 644 2684
rect 684 2676 692 2684
rect 748 2676 756 2684
rect 5308 2694 5316 2702
rect 1036 2676 1044 2684
rect 1324 2676 1332 2684
rect 1340 2676 1348 2684
rect 1388 2676 1396 2684
rect 1548 2676 1556 2684
rect 1676 2676 1684 2684
rect 1820 2676 1828 2684
rect 1884 2676 1892 2684
rect 1916 2676 1924 2684
rect 1948 2676 1956 2684
rect 2156 2676 2164 2684
rect 2380 2676 2388 2684
rect 2412 2676 2420 2684
rect 2540 2676 2548 2684
rect 2604 2676 2612 2684
rect 2698 2676 2706 2684
rect 2892 2676 2900 2684
rect 3164 2676 3172 2684
rect 3420 2676 3428 2684
rect 3612 2676 3620 2684
rect 3964 2676 3972 2684
rect 4332 2676 4340 2684
rect 4364 2676 4372 2684
rect 4396 2676 4404 2684
rect 4492 2676 4500 2684
rect 4732 2676 4740 2684
rect 5084 2676 5092 2684
rect 5276 2676 5284 2684
rect 5356 2676 5364 2684
rect 5516 2676 5524 2684
rect 188 2656 196 2664
rect 524 2656 532 2664
rect 764 2656 772 2664
rect 876 2656 884 2664
rect 1068 2656 1076 2664
rect 1516 2656 1524 2664
rect 1580 2656 1588 2664
rect 2044 2656 2052 2664
rect 2060 2656 2068 2664
rect 2140 2656 2148 2664
rect 2268 2656 2276 2664
rect 2444 2656 2452 2664
rect 2860 2656 2868 2664
rect 3196 2656 3204 2664
rect 3644 2656 3652 2664
rect 3996 2656 4004 2664
rect 4220 2656 4228 2664
rect 4300 2656 4308 2664
rect 4460 2656 4468 2664
rect 4700 2656 4708 2664
rect 5052 2656 5060 2664
rect 5244 2656 5252 2664
rect 460 2636 468 2644
rect 620 2636 628 2644
rect 700 2636 708 2644
rect 892 2636 900 2644
rect 1660 2636 1668 2644
rect 1788 2636 1796 2644
rect 2348 2636 2356 2644
rect 2524 2636 2532 2644
rect 3404 2636 3412 2644
rect 3468 2636 3476 2644
rect 3804 2636 3812 2644
rect 4204 2636 4212 2644
rect 4476 2636 4484 2644
rect 5228 2636 5236 2644
rect 2723 2606 2731 2614
rect 2733 2606 2741 2614
rect 2743 2606 2751 2614
rect 2753 2606 2761 2614
rect 2763 2606 2771 2614
rect 2773 2606 2781 2614
rect 300 2576 308 2584
rect 572 2576 580 2584
rect 1228 2576 1236 2584
rect 1372 2576 1380 2584
rect 1420 2576 1428 2584
rect 1772 2576 1780 2584
rect 1820 2576 1828 2584
rect 1884 2576 1892 2584
rect 1900 2576 1908 2584
rect 2076 2576 2084 2584
rect 2428 2576 2436 2584
rect 2892 2576 2900 2584
rect 3228 2576 3236 2584
rect 3372 2576 3380 2584
rect 3484 2576 3492 2584
rect 12 2556 20 2564
rect 44 2556 52 2564
rect 236 2556 244 2564
rect 412 2556 420 2564
rect 444 2556 452 2564
rect 636 2556 644 2564
rect 748 2556 756 2564
rect 812 2556 820 2564
rect 972 2556 980 2564
rect 1324 2556 1332 2564
rect 1436 2556 1444 2564
rect 1612 2556 1620 2564
rect 1996 2556 2004 2564
rect 2060 2556 2068 2564
rect 2236 2556 2244 2564
rect 2636 2556 2644 2564
rect 3052 2556 3060 2564
rect 3404 2556 3412 2564
rect 3660 2556 3668 2564
rect 3884 2556 3892 2564
rect 4060 2556 4068 2564
rect 4300 2556 4308 2564
rect 4508 2556 4516 2564
rect 4684 2556 4692 2564
rect 4780 2556 4788 2564
rect 4956 2556 4964 2564
rect 92 2536 100 2544
rect 140 2536 148 2544
rect 252 2536 260 2544
rect 316 2536 324 2544
rect 428 2536 436 2544
rect 540 2536 548 2544
rect 732 2536 740 2544
rect 1004 2536 1012 2544
rect 1228 2536 1236 2544
rect 1356 2536 1364 2544
rect 1388 2536 1396 2544
rect 1580 2536 1588 2544
rect 44 2516 52 2524
rect 76 2516 84 2524
rect 156 2516 164 2524
rect 204 2516 212 2524
rect 236 2516 244 2524
rect 268 2516 276 2524
rect 316 2516 324 2524
rect 348 2516 356 2524
rect 380 2516 388 2524
rect 492 2516 500 2524
rect 636 2516 644 2524
rect 684 2516 692 2524
rect 700 2516 708 2524
rect 716 2516 724 2524
rect 796 2516 804 2524
rect 1100 2516 1108 2524
rect 1212 2516 1220 2524
rect 1324 2516 1332 2524
rect 1404 2516 1412 2524
rect 1580 2516 1588 2524
rect 1852 2536 1860 2544
rect 2012 2536 2020 2544
rect 2268 2536 2276 2544
rect 2668 2536 2676 2544
rect 3084 2536 3092 2544
rect 3276 2536 3284 2544
rect 3292 2536 3300 2544
rect 3340 2536 3348 2544
rect 3388 2536 3396 2544
rect 3628 2536 3636 2544
rect 4092 2536 4100 2544
rect 4346 2536 4354 2544
rect 4540 2536 4548 2544
rect 4716 2536 4724 2544
rect 4764 2536 4772 2544
rect 4924 2536 4932 2544
rect 5148 2536 5156 2544
rect 5276 2536 5284 2544
rect 1980 2516 1988 2524
rect 2332 2516 2340 2524
rect 2556 2516 2564 2524
rect 2972 2516 2980 2524
rect 124 2496 132 2504
rect 364 2496 372 2504
rect 460 2496 468 2504
rect 476 2496 484 2504
rect 572 2496 580 2504
rect 588 2496 596 2504
rect 684 2496 692 2504
rect 1068 2500 1076 2508
rect 1516 2500 1524 2508
rect 3356 2516 3364 2524
rect 3452 2516 3460 2524
rect 3548 2516 3556 2524
rect 3628 2516 3636 2524
rect 4188 2516 4196 2524
rect 4428 2516 4436 2524
rect 4620 2516 4628 2524
rect 4700 2516 4708 2524
rect 4732 2516 4740 2524
rect 4748 2516 4756 2524
rect 4828 2516 4836 2524
rect 5118 2516 5126 2524
rect 5356 2516 5364 2524
rect 5420 2518 5428 2526
rect 1884 2496 1892 2504
rect 1932 2496 1940 2504
rect 2364 2496 2372 2504
rect 2412 2496 2420 2504
rect 2764 2496 2772 2504
rect 3180 2496 3188 2504
rect 3228 2496 3236 2504
rect 3292 2496 3300 2504
rect 3484 2496 3492 2504
rect 3564 2500 3572 2508
rect 4156 2500 4164 2508
rect 4604 2500 4612 2508
rect 4860 2500 4868 2508
rect 5324 2496 5332 2504
rect 108 2476 116 2484
rect 508 2476 516 2484
rect 3836 2476 3844 2484
rect 764 2456 772 2464
rect 1068 2454 1076 2462
rect 1516 2454 1524 2462
rect 2556 2454 2564 2462
rect 2972 2454 2980 2462
rect 3564 2454 3572 2462
rect 4316 2456 4324 2464
rect 4604 2454 4612 2462
rect 4860 2454 4868 2462
rect 76 2436 84 2444
rect 188 2436 196 2444
rect 300 2436 308 2444
rect 396 2436 404 2444
rect 524 2436 532 2444
rect 652 2436 660 2444
rect 2364 2436 2372 2444
rect 2476 2436 2484 2444
rect 3852 2436 3860 2444
rect 4156 2436 4164 2444
rect 1219 2406 1227 2414
rect 1229 2406 1237 2414
rect 1239 2406 1247 2414
rect 1249 2406 1257 2414
rect 1259 2406 1267 2414
rect 1269 2406 1277 2414
rect 4227 2406 4235 2414
rect 4237 2406 4245 2414
rect 4247 2406 4255 2414
rect 4257 2406 4265 2414
rect 4267 2406 4275 2414
rect 4277 2406 4285 2414
rect 316 2376 324 2384
rect 412 2376 420 2384
rect 1468 2376 1476 2384
rect 1756 2376 1764 2384
rect 1820 2376 1828 2384
rect 1948 2376 1956 2384
rect 2348 2376 2356 2384
rect 3212 2376 3220 2384
rect 3564 2376 3572 2384
rect 3612 2376 3620 2384
rect 3788 2376 3796 2384
rect 4412 2376 4420 2384
rect 4588 2376 4596 2384
rect 4652 2376 4660 2384
rect 5260 2376 5268 2384
rect 5516 2376 5524 2384
rect 396 2336 404 2344
rect 684 2336 692 2344
rect 1308 2358 1316 2366
rect 2668 2358 2676 2366
rect 3052 2356 3060 2364
rect 4044 2358 4052 2366
rect 4300 2356 4308 2364
rect 716 2336 724 2344
rect 780 2336 788 2344
rect 1500 2336 1508 2344
rect 1708 2336 1716 2344
rect 1772 2336 1780 2344
rect 2044 2336 2052 2344
rect 4220 2336 4228 2344
rect 4316 2336 4324 2344
rect 4396 2336 4404 2344
rect 4604 2336 4612 2344
rect 4668 2336 4676 2344
rect 316 2316 324 2324
rect 364 2316 372 2324
rect 444 2316 452 2324
rect 620 2316 628 2324
rect 716 2316 724 2324
rect 1308 2312 1316 2320
rect 1532 2316 1540 2324
rect 1564 2316 1572 2324
rect 1644 2316 1652 2324
rect 1660 2316 1668 2324
rect 1788 2316 1796 2324
rect 1804 2316 1812 2324
rect 1900 2316 1908 2324
rect 1916 2316 1924 2324
rect 2028 2316 2036 2324
rect 2348 2316 2356 2324
rect 2668 2312 2676 2320
rect 3116 2312 3124 2320
rect 3244 2316 3252 2324
rect 3308 2316 3316 2324
rect 3324 2316 3332 2324
rect 3388 2316 3396 2324
rect 3596 2316 3604 2324
rect 3660 2316 3668 2324
rect 3756 2316 3764 2324
rect 4044 2312 4052 2320
rect 4268 2316 4276 2324
rect 4284 2316 4292 2324
rect 4412 2316 4420 2324
rect 4460 2316 4468 2324
rect 4492 2316 4500 2324
rect 4556 2316 4564 2324
rect 4572 2316 4580 2324
rect 4636 2316 4644 2324
rect 4764 2316 4772 2324
rect 4876 2316 4884 2324
rect 4892 2316 4900 2324
rect 5260 2316 5268 2324
rect 5372 2316 5380 2324
rect 284 2296 292 2304
rect 380 2296 388 2304
rect 444 2296 452 2304
rect 476 2296 484 2304
rect 508 2296 516 2304
rect 588 2296 596 2304
rect 700 2296 708 2304
rect 748 2296 756 2304
rect 844 2296 852 2304
rect 892 2296 900 2304
rect 924 2296 932 2304
rect 1020 2296 1028 2304
rect 1050 2296 1058 2304
rect 1340 2296 1348 2304
rect 1580 2296 1588 2304
rect 1612 2296 1620 2304
rect 1628 2296 1636 2304
rect 1852 2296 1860 2304
rect 1916 2296 1924 2304
rect 1948 2296 1956 2304
rect 1996 2296 2004 2304
rect 2332 2296 2340 2304
rect 2348 2296 2356 2304
rect 2492 2296 2500 2304
rect 2700 2296 2708 2304
rect 3052 2296 3060 2304
rect 3212 2296 3220 2304
rect 3276 2296 3284 2304
rect 3356 2296 3364 2304
rect 3372 2296 3380 2304
rect 3420 2296 3428 2304
rect 3484 2296 3492 2304
rect 3564 2296 3572 2304
rect 3644 2296 3652 2304
rect 3676 2296 3684 2304
rect 3692 2296 3700 2304
rect 3772 2296 3780 2304
rect 3868 2296 3876 2304
rect 4172 2296 4180 2304
rect 4300 2296 4308 2304
rect 4348 2296 4356 2304
rect 4364 2296 4372 2304
rect 4412 2296 4420 2304
rect 4524 2296 4532 2304
rect 4540 2296 4548 2304
rect 4588 2296 4596 2304
rect 4652 2296 4660 2304
rect 4732 2296 4740 2304
rect 4780 2296 4788 2304
rect 4796 2296 4804 2304
rect 4844 2296 4852 2304
rect 5052 2296 5060 2304
rect 5356 2296 5364 2304
rect 5420 2296 5428 2304
rect 5452 2296 5460 2304
rect 5468 2296 5476 2304
rect 220 2276 228 2284
rect 428 2276 436 2284
rect 492 2276 500 2284
rect 508 2276 516 2284
rect 604 2276 612 2284
rect 652 2276 660 2284
rect 732 2276 740 2284
rect 828 2276 836 2284
rect 1004 2276 1012 2284
rect 1244 2276 1252 2284
rect 1452 2276 1460 2284
rect 1580 2276 1588 2284
rect 1596 2276 1604 2284
rect 1660 2276 1668 2284
rect 1692 2276 1700 2284
rect 1708 2276 1716 2284
rect 1724 2280 1732 2288
rect 1772 2276 1780 2284
rect 1868 2276 1876 2284
rect 1964 2276 1972 2284
rect 1980 2276 1988 2284
rect 2252 2276 2260 2284
rect 2604 2276 2612 2284
rect 2828 2276 2836 2284
rect 3052 2276 3060 2284
rect 3196 2276 3204 2284
rect 3260 2276 3268 2284
rect 3292 2276 3300 2284
rect 3324 2276 3332 2284
rect 3372 2276 3380 2284
rect 3436 2276 3444 2284
rect 3532 2276 3540 2284
rect 3548 2276 3556 2284
rect 3708 2276 3716 2284
rect 3724 2276 3732 2284
rect 3980 2276 3988 2284
rect 4188 2276 4196 2284
rect 4460 2276 4468 2284
rect 4508 2276 4516 2284
rect 4700 2276 4708 2284
rect 4796 2276 4804 2284
rect 4860 2276 4868 2284
rect 4940 2276 4948 2284
rect 4970 2276 4978 2284
rect 5164 2276 5172 2284
rect 5340 2276 5348 2284
rect 5372 2276 5380 2284
rect 5404 2276 5412 2284
rect 188 2256 196 2264
rect 540 2256 548 2264
rect 620 2256 628 2264
rect 796 2256 804 2264
rect 860 2256 868 2264
rect 972 2256 980 2264
rect 1212 2256 1220 2264
rect 1516 2256 1524 2264
rect 2044 2256 2052 2264
rect 2220 2256 2228 2264
rect 2396 2256 2404 2264
rect 2572 2256 2580 2264
rect 2764 2256 2772 2264
rect 3020 2256 3028 2264
rect 3788 2256 3796 2264
rect 3948 2256 3956 2264
rect 4124 2256 4132 2264
rect 4380 2256 4388 2264
rect 4700 2256 4708 2264
rect 4748 2256 4756 2264
rect 4844 2256 4852 2264
rect 5132 2256 5140 2264
rect 5308 2256 5316 2264
rect 5420 2256 5428 2264
rect 28 2236 36 2244
rect 396 2236 404 2244
rect 556 2236 564 2244
rect 668 2236 676 2244
rect 812 2236 820 2244
rect 956 2236 964 2244
rect 988 2236 996 2244
rect 1468 2236 1476 2244
rect 2060 2236 2068 2244
rect 2860 2236 2868 2244
rect 4140 2236 4148 2244
rect 4908 2236 4916 2244
rect 5324 2236 5332 2244
rect 5372 2236 5380 2244
rect 2723 2206 2731 2214
rect 2733 2206 2741 2214
rect 2743 2206 2751 2214
rect 2753 2206 2761 2214
rect 2763 2206 2771 2214
rect 2773 2206 2781 2214
rect 156 2176 164 2184
rect 572 2176 580 2184
rect 860 2176 868 2184
rect 956 2176 964 2184
rect 1132 2176 1140 2184
rect 1756 2176 1764 2184
rect 2092 2176 2100 2184
rect 2892 2176 2900 2184
rect 3436 2176 3444 2184
rect 3452 2176 3460 2184
rect 3884 2176 3892 2184
rect 4332 2176 4340 2184
rect 4812 2176 4820 2184
rect 60 2156 68 2164
rect 508 2156 516 2164
rect 972 2156 980 2164
rect 1324 2156 1332 2164
rect 1516 2156 1524 2164
rect 1548 2156 1556 2164
rect 1692 2156 1700 2164
rect 1772 2156 1780 2164
rect 1884 2156 1892 2164
rect 2636 2156 2644 2164
rect 2860 2156 2868 2164
rect 2924 2156 2932 2164
rect 3084 2156 3092 2164
rect 3260 2156 3268 2164
rect 3420 2156 3428 2164
rect 3788 2156 3796 2164
rect 4156 2156 4164 2164
rect 4380 2156 4388 2164
rect 4412 2156 4420 2164
rect 4460 2156 4468 2164
rect 4972 2156 4980 2164
rect 5308 2156 5316 2164
rect 44 2136 52 2144
rect 60 2116 68 2124
rect 92 2116 100 2124
rect 124 2136 132 2144
rect 172 2136 180 2144
rect 188 2136 196 2144
rect 220 2136 228 2144
rect 300 2136 308 2144
rect 364 2136 372 2144
rect 524 2136 532 2144
rect 828 2136 836 2144
rect 892 2136 900 2144
rect 940 2136 948 2144
rect 972 2136 980 2144
rect 1036 2136 1044 2144
rect 1292 2136 1300 2144
rect 1564 2136 1572 2144
rect 1580 2136 1588 2144
rect 1612 2136 1620 2144
rect 1644 2136 1652 2144
rect 1676 2136 1684 2144
rect 1740 2136 1748 2144
rect 1788 2136 1796 2144
rect 1964 2136 1972 2144
rect 2092 2136 2100 2144
rect 2124 2136 2132 2144
rect 2156 2136 2164 2144
rect 2188 2136 2196 2144
rect 2204 2136 2212 2144
rect 2268 2136 2276 2144
rect 2444 2136 2452 2144
rect 2668 2136 2676 2144
rect 3116 2136 3124 2144
rect 3324 2136 3332 2144
rect 3420 2136 3428 2144
rect 3612 2136 3620 2144
rect 3660 2136 3668 2144
rect 3692 2136 3700 2144
rect 3708 2136 3716 2144
rect 3740 2136 3748 2144
rect 3788 2136 3796 2144
rect 3804 2136 3812 2144
rect 3820 2136 3828 2144
rect 3852 2136 3860 2144
rect 3900 2136 3908 2144
rect 3948 2136 3956 2144
rect 3964 2136 3972 2144
rect 4028 2136 4036 2144
rect 4044 2136 4052 2144
rect 4076 2136 4084 2144
rect 4108 2136 4116 2144
rect 4156 2136 4164 2144
rect 4236 2136 4244 2144
rect 4284 2136 4292 2144
rect 4348 2136 4356 2144
rect 4476 2136 4484 2144
rect 4540 2136 4548 2144
rect 4556 2136 4564 2144
rect 4588 2136 4596 2144
rect 4620 2136 4628 2144
rect 4732 2136 4740 2144
rect 5004 2136 5012 2144
rect 5276 2136 5284 2144
rect 172 2116 180 2124
rect 268 2116 276 2124
rect 316 2116 324 2124
rect 348 2116 356 2124
rect 380 2116 388 2124
rect 460 2116 468 2124
rect 540 2116 548 2124
rect 636 2116 644 2124
rect 700 2116 708 2124
rect 764 2116 772 2124
rect 924 2116 932 2124
rect 1052 2116 1060 2124
rect 1292 2116 1300 2124
rect 1404 2116 1412 2124
rect 1516 2116 1524 2124
rect 1628 2116 1636 2124
rect 1740 2116 1748 2124
rect 1804 2116 1812 2124
rect 1836 2116 1844 2124
rect 1852 2116 1860 2124
rect 1916 2116 1924 2124
rect 1980 2116 1988 2124
rect 2044 2116 2052 2124
rect 2076 2116 2084 2124
rect 2140 2116 2148 2124
rect 2220 2116 2228 2124
rect 2268 2116 2276 2124
rect 2284 2116 2292 2124
rect 2332 2116 2340 2124
rect 2396 2116 2404 2124
rect 2460 2116 2468 2124
rect 2764 2116 2772 2124
rect 3004 2116 3012 2124
rect 3308 2116 3316 2124
rect 188 2096 196 2104
rect 284 2096 292 2104
rect 476 2096 484 2104
rect 620 2096 628 2104
rect 684 2096 692 2104
rect 748 2096 756 2104
rect 876 2096 884 2104
rect 1004 2096 1012 2104
rect 1020 2096 1028 2104
rect 1084 2096 1092 2104
rect 1196 2096 1204 2104
rect 1596 2096 1604 2104
rect 1660 2096 1668 2104
rect 1948 2096 1956 2104
rect 1996 2096 2004 2104
rect 2060 2096 2068 2104
rect 2156 2096 2164 2104
rect 2172 2096 2180 2104
rect 2252 2096 2260 2104
rect 2316 2096 2324 2104
rect 2396 2096 2404 2104
rect 2732 2100 2740 2108
rect 3180 2100 3188 2108
rect 3388 2116 3396 2124
rect 3580 2118 3588 2126
rect 3676 2116 3684 2124
rect 3724 2116 3732 2124
rect 3772 2116 3780 2124
rect 3836 2116 3844 2124
rect 3916 2116 3924 2124
rect 3980 2116 3988 2124
rect 4012 2116 4020 2124
rect 4060 2116 4068 2124
rect 4092 2116 4100 2124
rect 4124 2116 4132 2124
rect 4284 2116 4292 2124
rect 4300 2116 4308 2124
rect 4364 2116 4372 2124
rect 4412 2116 4420 2124
rect 4428 2116 4436 2124
rect 4492 2116 4500 2124
rect 4524 2116 4532 2124
rect 4604 2116 4612 2124
rect 4636 2116 4644 2124
rect 4652 2116 4660 2124
rect 4716 2116 4724 2124
rect 4748 2116 4756 2124
rect 4764 2116 4772 2124
rect 5068 2116 5076 2124
rect 5180 2116 5188 2124
rect 3356 2096 3364 2104
rect 3644 2096 3652 2104
rect 3884 2096 3892 2104
rect 3948 2096 3956 2104
rect 4172 2096 4180 2104
rect 4780 2096 4788 2104
rect 5100 2096 5108 2104
rect 5212 2100 5220 2108
rect 252 2076 260 2084
rect 300 2076 308 2084
rect 444 2076 452 2084
rect 652 2076 660 2084
rect 716 2076 724 2084
rect 780 2076 788 2084
rect 1916 2076 1924 2084
rect 2028 2076 2036 2084
rect 4444 2076 4452 2084
rect 4492 2076 4500 2084
rect 5500 2076 5508 2084
rect 268 2056 276 2064
rect 3004 2054 3012 2062
rect 5212 2054 5220 2062
rect 28 2036 36 2044
rect 412 2036 420 2044
rect 460 2036 468 2044
rect 636 2036 644 2044
rect 732 2036 740 2044
rect 1196 2036 1204 2044
rect 1756 2036 1764 2044
rect 2012 2036 2020 2044
rect 2476 2036 2484 2044
rect 2732 2036 2740 2044
rect 2924 2036 2932 2044
rect 4012 2036 4020 2044
rect 4140 2036 4148 2044
rect 4684 2036 4692 2044
rect 4812 2036 4820 2044
rect 5100 2036 5108 2044
rect 1219 2006 1227 2014
rect 1229 2006 1237 2014
rect 1239 2006 1247 2014
rect 1249 2006 1257 2014
rect 1259 2006 1267 2014
rect 1269 2006 1277 2014
rect 4227 2006 4235 2014
rect 4237 2006 4245 2014
rect 4247 2006 4255 2014
rect 4257 2006 4265 2014
rect 4267 2006 4275 2014
rect 4277 2006 4285 2014
rect 428 1976 436 1984
rect 572 1976 580 1984
rect 988 1976 996 1984
rect 1468 1976 1476 1984
rect 1756 1976 1764 1984
rect 1836 1976 1844 1984
rect 2124 1976 2132 1984
rect 2236 1976 2244 1984
rect 3932 1976 3940 1984
rect 4076 1976 4084 1984
rect 4108 1976 4116 1984
rect 4204 1976 4212 1984
rect 4476 1976 4484 1984
rect 4652 1976 4660 1984
rect 4700 1976 4708 1984
rect 4988 1976 4996 1984
rect 5084 1976 5092 1984
rect 5148 1976 5156 1984
rect 5420 1976 5428 1984
rect 316 1956 324 1964
rect 732 1958 740 1966
rect 1228 1956 1236 1964
rect 2940 1958 2948 1966
rect 3228 1956 3236 1964
rect 3596 1956 3604 1964
rect 364 1936 372 1944
rect 412 1936 420 1944
rect 556 1936 564 1944
rect 2220 1936 2228 1944
rect 3916 1936 3924 1944
rect 4124 1936 4132 1944
rect 4156 1936 4164 1944
rect 4300 1936 4308 1944
rect 4460 1936 4468 1944
rect 4604 1936 4612 1944
rect 44 1916 52 1924
rect 60 1916 68 1924
rect 332 1916 340 1924
rect 444 1916 452 1924
rect 524 1916 532 1924
rect 588 1916 596 1924
rect 732 1912 740 1920
rect 1292 1912 1300 1920
rect 1468 1916 1476 1924
rect 2124 1916 2132 1924
rect 2332 1916 2340 1924
rect 108 1896 116 1904
rect 220 1896 228 1904
rect 252 1896 260 1904
rect 348 1896 356 1904
rect 428 1896 436 1904
rect 572 1896 580 1904
rect 620 1896 628 1904
rect 652 1896 660 1904
rect 908 1896 916 1904
rect 1228 1896 1236 1904
rect 1484 1896 1492 1904
rect 1916 1896 1924 1904
rect 2108 1896 2116 1904
rect 2188 1896 2196 1904
rect 2236 1896 2244 1904
rect 2348 1896 2356 1904
rect 2524 1916 2532 1924
rect 2940 1912 2948 1920
rect 3324 1916 3332 1924
rect 3452 1916 3460 1924
rect 3532 1912 3540 1920
rect 3804 1916 3812 1924
rect 3884 1916 3892 1924
rect 3948 1916 3956 1924
rect 4044 1916 4052 1924
rect 4092 1916 4100 1924
rect 4236 1916 4244 1924
rect 4332 1916 4340 1924
rect 4492 1916 4500 1924
rect 4604 1916 4612 1924
rect 4620 1916 4628 1924
rect 4988 1916 4996 1924
rect 2492 1896 2500 1904
rect 2540 1896 2548 1904
rect 2682 1896 2690 1904
rect 2972 1896 2980 1904
rect 3228 1896 3236 1904
rect 3420 1896 3428 1904
rect 3596 1896 3604 1904
rect 3790 1896 3798 1904
rect 3852 1896 3860 1904
rect 3900 1896 3908 1904
rect 4012 1896 4020 1904
rect 4108 1896 4116 1904
rect 4172 1896 4180 1904
rect 4348 1896 4356 1904
rect 4364 1896 4372 1904
rect 4412 1896 4420 1904
rect 4476 1896 4484 1904
rect 4508 1896 4516 1904
rect 4588 1896 4596 1904
rect 4652 1896 4660 1904
rect 4780 1896 4788 1904
rect 4972 1896 4980 1904
rect 5052 1896 5060 1904
rect 5084 1896 5092 1904
rect 5116 1896 5124 1904
rect 5132 1896 5140 1904
rect 5180 1896 5188 1904
rect 5276 1896 5284 1904
rect 5308 1896 5316 1904
rect 5420 1896 5428 1904
rect 5468 1916 5476 1924
rect 12 1876 20 1884
rect 92 1876 100 1884
rect 172 1880 180 1888
rect 284 1876 292 1884
rect 348 1876 356 1884
rect 492 1876 500 1884
rect 604 1876 612 1884
rect 796 1876 804 1884
rect 1228 1876 1236 1884
rect 1564 1876 1572 1884
rect 1820 1876 1828 1884
rect 2028 1876 2036 1884
rect 2300 1876 2308 1884
rect 2668 1876 2676 1884
rect 2876 1876 2884 1884
rect 3228 1876 3236 1884
rect 3452 1876 3460 1884
rect 3596 1876 3604 1884
rect 3868 1876 3876 1884
rect 3980 1876 3988 1884
rect 3996 1876 4004 1884
rect 4188 1876 4196 1884
rect 4588 1876 4596 1884
rect 4668 1876 4676 1884
rect 4892 1876 4900 1884
rect 5036 1876 5044 1884
rect 5100 1876 5108 1884
rect 5404 1876 5412 1884
rect 5500 1876 5508 1884
rect 140 1856 148 1864
rect 220 1856 228 1864
rect 268 1856 276 1864
rect 460 1856 468 1864
rect 828 1856 836 1864
rect 1196 1856 1204 1864
rect 1596 1856 1604 1864
rect 1996 1856 2004 1864
rect 2188 1856 2196 1864
rect 2284 1856 2292 1864
rect 2380 1856 2388 1864
rect 2444 1856 2452 1864
rect 2636 1856 2644 1864
rect 2844 1856 2852 1864
rect 3196 1856 3204 1864
rect 3372 1856 3380 1864
rect 3628 1856 3636 1864
rect 3804 1856 3812 1864
rect 3948 1856 3956 1864
rect 4060 1856 4068 1864
rect 4172 1856 4180 1864
rect 4332 1856 4340 1864
rect 4860 1856 4868 1864
rect 44 1836 52 1844
rect 76 1836 84 1844
rect 204 1836 212 1844
rect 476 1836 484 1844
rect 524 1836 532 1844
rect 1036 1836 1044 1844
rect 1788 1836 1796 1844
rect 2332 1836 2340 1844
rect 2396 1836 2404 1844
rect 3036 1836 3044 1844
rect 4044 1836 4052 1844
rect 4396 1836 4404 1844
rect 4540 1836 4548 1844
rect 5388 1836 5396 1844
rect 2723 1806 2731 1814
rect 2733 1806 2741 1814
rect 2743 1806 2751 1814
rect 2753 1806 2761 1814
rect 2763 1806 2771 1814
rect 2773 1806 2781 1814
rect 364 1776 372 1784
rect 492 1776 500 1784
rect 524 1776 532 1784
rect 572 1776 580 1784
rect 2540 1776 2548 1784
rect 2588 1776 2596 1784
rect 2716 1776 2724 1784
rect 3420 1776 3428 1784
rect 3628 1776 3636 1784
rect 4636 1776 4644 1784
rect 4748 1776 4756 1784
rect 4876 1776 4884 1784
rect 5116 1776 5124 1784
rect 5148 1776 5156 1784
rect 12 1756 20 1764
rect 76 1756 84 1764
rect 92 1756 100 1764
rect 124 1756 132 1764
rect 188 1756 196 1764
rect 220 1756 228 1764
rect 236 1756 244 1764
rect 428 1756 436 1764
rect 732 1756 740 1764
rect 1004 1756 1012 1764
rect 1340 1756 1348 1764
rect 1676 1756 1684 1764
rect 1932 1756 1940 1764
rect 1996 1756 2004 1764
rect 2188 1756 2196 1764
rect 2364 1756 2372 1764
rect 2444 1756 2452 1764
rect 2572 1756 2580 1764
rect 2700 1756 2708 1764
rect 2892 1756 2900 1764
rect 2908 1756 2916 1764
rect 3116 1756 3124 1764
rect 3340 1756 3348 1764
rect 3532 1756 3540 1764
rect 3564 1756 3572 1764
rect 3804 1756 3812 1764
rect 4092 1756 4100 1764
rect 4108 1756 4116 1764
rect 4348 1756 4356 1764
rect 4556 1756 4564 1764
rect 4652 1756 4660 1764
rect 4908 1756 4916 1764
rect 5020 1756 5028 1764
rect 5308 1756 5316 1764
rect 204 1736 212 1744
rect 380 1736 388 1744
rect 444 1736 452 1744
rect 460 1736 468 1744
rect 540 1736 548 1744
rect 764 1736 772 1744
rect 908 1736 916 1744
rect 1052 1736 1060 1744
rect 1068 1736 1076 1744
rect 1372 1736 1380 1744
rect 1644 1736 1652 1744
rect 1868 1736 1876 1744
rect 2220 1736 2228 1744
rect 2380 1736 2388 1744
rect 2460 1736 2468 1744
rect 2508 1736 2516 1744
rect 2556 1736 2564 1744
rect 2604 1736 2612 1744
rect 2652 1736 2660 1744
rect 2732 1736 2740 1744
rect 2828 1736 2836 1744
rect 2860 1736 2868 1744
rect 3148 1736 3156 1744
rect 3324 1736 3332 1744
rect 3484 1736 3492 1744
rect 3772 1736 3780 1744
rect 4380 1736 4388 1744
rect 4572 1736 4580 1744
rect 4604 1736 4612 1744
rect 4812 1736 4820 1744
rect 4988 1736 4996 1744
rect 5020 1736 5028 1744
rect 5052 1736 5060 1744
rect 5084 1736 5092 1744
rect 5228 1736 5236 1744
rect 5340 1736 5348 1744
rect 92 1716 100 1724
rect 124 1716 132 1724
rect 140 1716 148 1724
rect 284 1716 292 1724
rect 332 1716 340 1724
rect 396 1716 404 1724
rect 428 1716 436 1724
rect 860 1716 868 1724
rect 924 1716 932 1724
rect 972 1716 980 1724
rect 1004 1716 1012 1724
rect 1100 1716 1108 1724
rect 1260 1716 1268 1724
rect 1532 1716 1540 1724
rect 1756 1716 1764 1724
rect 1964 1716 1972 1724
rect 2108 1716 2116 1724
rect 2220 1716 2228 1724
rect 2412 1716 2420 1724
rect 2492 1716 2500 1724
rect 2620 1716 2628 1724
rect 2668 1716 2676 1724
rect 2812 1716 2820 1724
rect 2844 1716 2852 1724
rect 2924 1716 2932 1724
rect 3212 1716 3220 1724
rect 3244 1716 3252 1724
rect 3388 1716 3396 1724
rect 156 1696 164 1704
rect 300 1696 308 1704
rect 492 1696 500 1704
rect 828 1700 836 1708
rect 956 1696 964 1704
rect 1468 1696 1476 1704
rect 1548 1696 1556 1704
rect 1900 1696 1908 1704
rect 2316 1696 2324 1704
rect 2460 1696 2468 1704
rect 2524 1696 2532 1704
rect 2684 1696 2692 1704
rect 2876 1696 2884 1704
rect 3244 1696 3252 1704
rect 3292 1696 3300 1704
rect 3484 1716 3492 1724
rect 3500 1716 3508 1724
rect 3596 1716 3604 1724
rect 3884 1716 3892 1724
rect 4028 1716 4036 1724
rect 4060 1716 4068 1724
rect 4476 1716 4484 1724
rect 4524 1716 4532 1724
rect 4556 1716 4564 1724
rect 4620 1716 4628 1724
rect 4700 1716 4708 1724
rect 4764 1716 4772 1724
rect 4780 1716 4788 1724
rect 4844 1716 4852 1724
rect 4956 1716 4964 1724
rect 5068 1716 5076 1724
rect 3436 1696 3444 1704
rect 3628 1696 3636 1704
rect 3708 1700 3716 1708
rect 4028 1696 4036 1704
rect 4444 1700 4452 1708
rect 4716 1696 4724 1704
rect 4828 1696 4836 1704
rect 4972 1696 4980 1704
rect 5116 1696 5124 1704
rect 5404 1700 5412 1708
rect 300 1676 308 1684
rect 316 1676 324 1684
rect 2652 1676 2660 1684
rect 4012 1676 4020 1684
rect 4044 1676 4052 1684
rect 4684 1676 4692 1684
rect 4748 1676 4756 1684
rect 4796 1676 4804 1684
rect 4860 1676 4868 1684
rect 4892 1676 4900 1684
rect 4940 1676 4948 1684
rect 1260 1654 1268 1662
rect 4444 1654 4452 1662
rect 4668 1656 4676 1664
rect 5404 1654 5412 1662
rect 284 1636 292 1644
rect 828 1636 836 1644
rect 1180 1636 1188 1644
rect 1548 1636 1556 1644
rect 1836 1636 1844 1644
rect 2028 1636 2036 1644
rect 2316 1636 2324 1644
rect 3244 1636 3252 1644
rect 3308 1636 3316 1644
rect 3532 1636 3540 1644
rect 3708 1636 3716 1644
rect 3964 1636 3972 1644
rect 4028 1636 4036 1644
rect 4076 1636 4084 1644
rect 4540 1636 4548 1644
rect 4876 1636 4884 1644
rect 4956 1636 4964 1644
rect 5020 1636 5028 1644
rect 1219 1606 1227 1614
rect 1229 1606 1237 1614
rect 1239 1606 1247 1614
rect 1249 1606 1257 1614
rect 1259 1606 1267 1614
rect 1269 1606 1277 1614
rect 4227 1606 4235 1614
rect 4237 1606 4245 1614
rect 4247 1606 4255 1614
rect 4257 1606 4265 1614
rect 4267 1606 4275 1614
rect 4277 1606 4285 1614
rect 428 1576 436 1584
rect 1516 1576 1524 1584
rect 2588 1576 2596 1584
rect 2700 1576 2708 1584
rect 2860 1576 2868 1584
rect 3548 1576 3556 1584
rect 4620 1576 4628 1584
rect 4972 1576 4980 1584
rect 5100 1576 5108 1584
rect 5212 1576 5220 1584
rect 5436 1576 5444 1584
rect 972 1558 980 1566
rect 1212 1556 1220 1564
rect 2284 1558 2292 1566
rect 3148 1556 3156 1564
rect 76 1536 84 1544
rect 364 1536 372 1544
rect 1900 1536 1908 1544
rect 2716 1536 2724 1544
rect 3980 1536 3988 1544
rect 4044 1536 4052 1544
rect 4556 1536 4564 1544
rect 4572 1536 4580 1544
rect 4636 1536 4644 1544
rect 5116 1536 5124 1544
rect 60 1516 68 1524
rect 444 1516 452 1524
rect 44 1496 52 1504
rect 76 1496 84 1504
rect 188 1496 196 1504
rect 284 1496 292 1504
rect 316 1496 324 1504
rect 364 1496 372 1504
rect 508 1496 516 1504
rect 588 1496 596 1504
rect 652 1516 660 1524
rect 972 1512 980 1520
rect 1068 1516 1076 1524
rect 1180 1516 1188 1524
rect 1516 1516 1524 1524
rect 1884 1516 1892 1524
rect 1932 1516 1940 1524
rect 2204 1516 2212 1524
rect 2284 1512 2292 1520
rect 2556 1516 2564 1524
rect 2684 1516 2692 1524
rect 3212 1512 3220 1520
rect 3260 1516 3268 1524
rect 3292 1516 3300 1524
rect 3388 1516 3396 1524
rect 3452 1516 3460 1524
rect 3516 1516 3524 1524
rect 3628 1516 3636 1524
rect 3676 1516 3684 1524
rect 3884 1516 3892 1524
rect 3964 1516 3972 1524
rect 4012 1516 4020 1524
rect 4076 1516 4084 1524
rect 4092 1516 4100 1524
rect 4236 1516 4244 1524
rect 4604 1516 4612 1524
rect 796 1496 804 1504
rect 1004 1496 1012 1504
rect 1052 1496 1060 1504
rect 1148 1496 1156 1504
rect 1356 1496 1364 1504
rect 1516 1496 1524 1504
rect 1724 1496 1732 1504
rect 1852 1496 1860 1504
rect 1996 1496 2004 1504
rect 2044 1496 2052 1504
rect 2108 1496 2116 1504
rect 2188 1496 2196 1504
rect 2252 1496 2260 1504
rect 2668 1496 2676 1504
rect 2700 1496 2708 1504
rect 2908 1496 2916 1504
rect 2954 1496 2962 1504
rect 3148 1496 3156 1504
rect 3324 1496 3332 1504
rect 3404 1496 3412 1504
rect 3420 1496 3428 1504
rect 3468 1496 3476 1504
rect 3484 1496 3492 1504
rect 3580 1496 3588 1504
rect 3596 1496 3604 1504
rect 3612 1496 3620 1504
rect 3676 1496 3684 1504
rect 3692 1496 3700 1504
rect 3756 1496 3764 1504
rect 3788 1496 3796 1504
rect 3836 1496 3844 1504
rect 3852 1496 3860 1504
rect 3868 1496 3876 1504
rect 3932 1496 3940 1504
rect 3996 1496 4004 1504
rect 4060 1496 4068 1504
rect 4108 1496 4116 1504
rect 4124 1496 4132 1504
rect 4188 1496 4196 1504
rect 4204 1496 4212 1504
rect 4252 1496 4260 1504
rect 4444 1496 4452 1504
rect 4572 1496 4580 1504
rect 4620 1496 4628 1504
rect 4716 1496 4724 1504
rect 4812 1496 4820 1504
rect 4860 1496 4868 1504
rect 4876 1496 4884 1504
rect 4940 1496 4948 1504
rect 4972 1496 4980 1504
rect 5020 1496 5028 1504
rect 5068 1496 5076 1504
rect 5084 1496 5092 1504
rect 5164 1496 5172 1504
rect 5180 1496 5188 1504
rect 5244 1496 5252 1504
rect 5308 1494 5316 1502
rect 5452 1496 5460 1504
rect 12 1476 20 1484
rect 204 1476 212 1484
rect 412 1476 420 1484
rect 444 1476 452 1484
rect 572 1476 580 1484
rect 652 1476 660 1484
rect 908 1476 916 1484
rect 1084 1476 1092 1484
rect 1164 1476 1172 1484
rect 1340 1476 1348 1484
rect 1612 1476 1620 1484
rect 1932 1476 1940 1484
rect 2060 1476 2068 1484
rect 2076 1476 2084 1484
rect 2156 1476 2164 1484
rect 2348 1476 2356 1484
rect 2604 1476 2612 1484
rect 2620 1476 2628 1484
rect 2652 1476 2660 1484
rect 2796 1476 2804 1484
rect 2828 1480 2836 1488
rect 2876 1476 2884 1484
rect 3148 1476 3156 1484
rect 3292 1476 3300 1484
rect 3436 1476 3444 1484
rect 3500 1476 3508 1484
rect 3564 1476 3572 1484
rect 3644 1476 3652 1484
rect 3708 1476 3716 1484
rect 3740 1476 3748 1484
rect 3772 1476 3780 1484
rect 3948 1476 3956 1484
rect 4268 1476 4276 1484
rect 4364 1476 4372 1484
rect 4524 1476 4532 1484
rect 4700 1476 4708 1484
rect 4924 1476 4932 1484
rect 4988 1476 4996 1484
rect 5324 1476 5332 1484
rect 5516 1476 5524 1484
rect 252 1456 260 1464
rect 284 1456 292 1464
rect 332 1456 340 1464
rect 364 1456 372 1464
rect 396 1456 404 1464
rect 492 1456 500 1464
rect 876 1456 884 1464
rect 1196 1456 1204 1464
rect 1644 1456 1652 1464
rect 1948 1456 1956 1464
rect 2012 1456 2020 1464
rect 2076 1456 2084 1464
rect 2380 1456 2388 1464
rect 2620 1456 2628 1464
rect 3116 1456 3124 1464
rect 3372 1456 3380 1464
rect 3884 1456 3892 1464
rect 4156 1456 4164 1464
rect 4540 1456 4548 1464
rect 4684 1456 4692 1464
rect 4892 1456 4900 1464
rect 4908 1456 4916 1464
rect 5116 1456 5124 1464
rect 5148 1456 5156 1464
rect 76 1436 84 1444
rect 204 1436 212 1444
rect 492 1436 500 1444
rect 716 1436 724 1444
rect 1116 1436 1124 1444
rect 1468 1436 1476 1444
rect 1804 1436 1812 1444
rect 2540 1436 2548 1444
rect 3724 1436 3732 1444
rect 4044 1436 4052 1444
rect 4172 1436 4180 1444
rect 4700 1436 4708 1444
rect 4828 1436 4836 1444
rect 5036 1436 5044 1444
rect 2723 1406 2731 1414
rect 2733 1406 2741 1414
rect 2743 1406 2751 1414
rect 2753 1406 2761 1414
rect 2763 1406 2771 1414
rect 2773 1406 2781 1414
rect 508 1376 516 1384
rect 892 1376 900 1384
rect 1548 1376 1556 1384
rect 1724 1376 1732 1384
rect 1756 1376 1764 1384
rect 2508 1376 2516 1384
rect 2652 1376 2660 1384
rect 3964 1376 3972 1384
rect 4508 1376 4516 1384
rect 4972 1376 4980 1384
rect 44 1356 52 1364
rect 124 1356 132 1364
rect 668 1356 676 1364
rect 844 1356 852 1364
rect 972 1356 980 1364
rect 1148 1356 1156 1364
rect 1420 1356 1428 1364
rect 1660 1356 1668 1364
rect 1820 1356 1828 1364
rect 1996 1356 2004 1364
rect 2172 1356 2180 1364
rect 2428 1356 2436 1364
rect 2460 1356 2468 1364
rect 2524 1356 2532 1364
rect 2540 1356 2548 1364
rect 2732 1356 2740 1364
rect 2892 1356 2900 1364
rect 3148 1356 3156 1364
rect 3388 1356 3396 1364
rect 3564 1356 3572 1364
rect 3580 1356 3588 1364
rect 3612 1356 3620 1364
rect 3628 1356 3636 1364
rect 28 1336 36 1344
rect 60 1336 68 1344
rect 172 1336 180 1344
rect 204 1336 212 1344
rect 364 1336 372 1344
rect 412 1336 420 1344
rect 700 1336 708 1344
rect 908 1336 916 1344
rect 940 1336 948 1344
rect 1116 1336 1124 1344
rect 1436 1336 1444 1344
rect 1612 1336 1620 1344
rect 1676 1336 1684 1344
rect 2028 1336 2036 1344
rect 2188 1336 2196 1344
rect 2268 1336 2276 1344
rect 2284 1336 2292 1344
rect 2492 1336 2500 1344
rect 2524 1336 2532 1344
rect 92 1316 100 1324
rect 156 1316 164 1324
rect 188 1316 196 1324
rect 268 1316 276 1324
rect 332 1316 340 1324
rect 380 1316 388 1324
rect 460 1316 468 1324
rect 700 1316 708 1324
rect 796 1316 804 1324
rect 924 1316 932 1324
rect 972 1316 980 1324
rect 1004 1316 1012 1324
rect 1228 1316 1236 1324
rect 1452 1316 1460 1324
rect 1516 1316 1524 1324
rect 1596 1316 1604 1324
rect 1628 1316 1636 1324
rect 1692 1316 1700 1324
rect 1724 1316 1732 1324
rect 76 1296 84 1304
rect 220 1296 228 1304
rect 284 1296 292 1304
rect 348 1296 356 1304
rect 412 1296 420 1304
rect 476 1296 484 1304
rect 764 1300 772 1308
rect 860 1296 868 1304
rect 1052 1300 1060 1308
rect 1500 1296 1508 1304
rect 1564 1296 1572 1304
rect 1724 1296 1732 1304
rect 1834 1316 1842 1324
rect 2108 1316 2116 1324
rect 2268 1316 2276 1324
rect 2300 1316 2308 1324
rect 2316 1316 2324 1324
rect 2332 1316 2340 1324
rect 2380 1316 2388 1324
rect 2492 1316 2500 1324
rect 2572 1316 2580 1324
rect 2924 1336 2932 1344
rect 3068 1336 3076 1344
rect 3164 1336 3172 1344
rect 3212 1336 3220 1344
rect 3356 1336 3364 1344
rect 3612 1336 3620 1344
rect 3644 1336 3652 1344
rect 3708 1336 3716 1344
rect 3740 1336 3748 1344
rect 3788 1356 3796 1364
rect 3932 1356 3940 1364
rect 4124 1356 4132 1364
rect 4364 1356 4372 1364
rect 4460 1356 4468 1364
rect 4636 1356 4644 1364
rect 4812 1356 4820 1364
rect 5148 1356 5156 1364
rect 5324 1356 5332 1364
rect 3820 1336 3828 1344
rect 3852 1336 3860 1344
rect 4156 1336 4164 1344
rect 4428 1336 4436 1344
rect 4540 1336 4548 1344
rect 4780 1336 4788 1344
rect 5100 1336 5108 1344
rect 5356 1336 5364 1344
rect 2604 1316 2612 1324
rect 2812 1316 2820 1324
rect 3100 1316 3108 1324
rect 3196 1316 3204 1324
rect 3260 1316 3268 1324
rect 3660 1316 3668 1324
rect 3676 1316 3684 1324
rect 3692 1316 3700 1324
rect 3724 1316 3732 1324
rect 3820 1316 3828 1324
rect 3836 1316 3844 1324
rect 3900 1316 3908 1324
rect 4252 1316 4260 1324
rect 4348 1316 4356 1324
rect 4396 1316 4404 1324
rect 4412 1316 4420 1324
rect 4492 1316 4500 1324
rect 4556 1316 4564 1324
rect 4588 1316 4596 1324
rect 4700 1316 4708 1324
rect 5004 1316 5012 1324
rect 5020 1316 5028 1324
rect 5068 1316 5076 1324
rect 5436 1316 5444 1324
rect 2124 1296 2132 1304
rect 2220 1296 2228 1304
rect 2332 1296 2340 1304
rect 2636 1296 2644 1304
rect 3036 1296 3044 1304
rect 3068 1296 3076 1304
rect 3148 1296 3156 1304
rect 3292 1300 3300 1308
rect 4220 1300 4228 1308
rect 4476 1296 4484 1304
rect 4684 1296 4692 1304
rect 5132 1296 5140 1304
rect 5452 1296 5460 1304
rect 252 1276 260 1284
rect 316 1276 324 1284
rect 492 1276 500 1284
rect 2364 1276 2372 1284
rect 3884 1276 3892 1284
rect 5100 1276 5108 1284
rect 332 1256 340 1264
rect 1052 1254 1060 1262
rect 2812 1254 2820 1262
rect 4220 1254 4228 1262
rect 12 1236 20 1244
rect 268 1236 276 1244
rect 460 1236 468 1244
rect 764 1236 772 1244
rect 1308 1236 1316 1244
rect 1372 1236 1380 1244
rect 2124 1236 2132 1244
rect 2460 1236 2468 1244
rect 2508 1236 2516 1244
rect 3292 1236 3300 1244
rect 3772 1236 3780 1244
rect 3916 1236 3924 1244
rect 4572 1236 4580 1244
rect 4684 1236 4692 1244
rect 5052 1236 5060 1244
rect 5452 1236 5460 1244
rect 1219 1206 1227 1214
rect 1229 1206 1237 1214
rect 1239 1206 1247 1214
rect 1249 1206 1257 1214
rect 1259 1206 1267 1214
rect 1269 1206 1277 1214
rect 4227 1206 4235 1214
rect 4237 1206 4245 1214
rect 4247 1206 4255 1214
rect 4257 1206 4265 1214
rect 4267 1206 4275 1214
rect 4277 1206 4285 1214
rect 44 1176 52 1184
rect 92 1176 100 1184
rect 220 1176 228 1184
rect 300 1176 308 1184
rect 732 1176 740 1184
rect 876 1176 884 1184
rect 1164 1176 1172 1184
rect 1196 1176 1204 1184
rect 1596 1176 1604 1184
rect 1836 1176 1844 1184
rect 3420 1176 3428 1184
rect 3820 1176 3828 1184
rect 3900 1176 3908 1184
rect 4444 1176 4452 1184
rect 4812 1176 4820 1184
rect 5180 1176 5188 1184
rect 5468 1176 5476 1184
rect 156 1156 164 1164
rect 2940 1156 2948 1164
rect 60 1136 68 1144
rect 140 1136 148 1144
rect 204 1136 212 1144
rect 284 1136 292 1144
rect 2124 1136 2132 1144
rect 4428 1136 4436 1144
rect 44 1116 52 1124
rect 108 1116 116 1124
rect 172 1116 180 1124
rect 236 1116 244 1124
rect 252 1116 260 1124
rect 316 1116 324 1124
rect 732 1116 740 1124
rect 828 1116 836 1124
rect 876 1116 884 1124
rect 1308 1116 1316 1124
rect 1532 1116 1540 1124
rect 1676 1116 1684 1124
rect 1708 1116 1716 1124
rect 1788 1116 1796 1124
rect 1836 1116 1844 1124
rect 2220 1116 2228 1124
rect 2268 1116 2276 1124
rect 2476 1116 2484 1124
rect 2588 1116 2596 1124
rect 3004 1112 3012 1120
rect 3036 1116 3044 1124
rect 3132 1116 3140 1124
rect 44 1096 52 1104
rect 156 1096 164 1104
rect 220 1096 228 1104
rect 268 1096 276 1104
rect 364 1096 372 1104
rect 700 1096 708 1104
rect 796 1096 804 1104
rect 876 1096 884 1104
rect 1084 1096 1092 1104
rect 1276 1096 1284 1104
rect 1388 1096 1396 1104
rect 1436 1096 1444 1104
rect 1484 1096 1492 1104
rect 1500 1096 1508 1104
rect 1548 1096 1556 1104
rect 1644 1096 1652 1104
rect 1676 1096 1684 1104
rect 1708 1096 1716 1104
rect 1836 1096 1844 1104
rect 2204 1096 2212 1104
rect 2252 1096 2260 1104
rect 2364 1096 2372 1104
rect 2508 1096 2516 1104
rect 2524 1096 2532 1104
rect 2746 1096 2754 1104
rect 2940 1096 2948 1104
rect 3100 1096 3108 1104
rect 3420 1116 3428 1124
rect 4140 1116 4148 1124
rect 4172 1116 4180 1124
rect 4396 1116 4404 1124
rect 4524 1116 4532 1124
rect 4620 1116 4628 1124
rect 4716 1116 4724 1124
rect 4972 1116 4980 1124
rect 3180 1096 3188 1104
rect 3420 1096 3428 1104
rect 3756 1096 3764 1104
rect 3788 1096 3796 1104
rect 3852 1096 3860 1104
rect 3916 1096 3924 1104
rect 3932 1096 3940 1104
rect 4076 1096 4084 1104
rect 4124 1096 4132 1104
rect 4172 1096 4180 1104
rect 4188 1096 4196 1104
rect 4332 1096 4340 1104
rect 4380 1096 4388 1104
rect 4412 1096 4420 1104
rect 4460 1096 4468 1104
rect 4556 1096 4564 1104
rect 4588 1096 4596 1104
rect 4636 1096 4644 1104
rect 4668 1096 4676 1104
rect 4716 1096 4724 1104
rect 4764 1096 4772 1104
rect 4828 1096 4836 1104
rect 4844 1096 4852 1104
rect 4860 1096 4868 1104
rect 4908 1096 4916 1104
rect 5004 1096 5012 1104
rect 5052 1116 5060 1124
rect 5100 1116 5108 1124
rect 5468 1116 5476 1124
rect 5132 1096 5140 1104
rect 5436 1096 5444 1104
rect 5452 1096 5460 1104
rect 76 1076 84 1084
rect 332 1076 340 1084
rect 364 1076 372 1084
rect 412 1076 420 1084
rect 636 1076 644 1084
rect 780 1076 788 1084
rect 972 1076 980 1084
rect 1372 1076 1380 1084
rect 1484 1076 1492 1084
rect 1516 1076 1524 1084
rect 1548 1076 1556 1084
rect 1756 1076 1764 1084
rect 1932 1076 1940 1084
rect 2156 1076 2164 1084
rect 2252 1076 2260 1084
rect 2332 1076 2340 1084
rect 2428 1076 2436 1084
rect 2460 1076 2468 1084
rect 2524 1076 2532 1084
rect 2540 1076 2548 1084
rect 2620 1076 2628 1084
rect 2940 1076 2948 1084
rect 3084 1076 3092 1084
rect 3164 1076 3172 1084
rect 3244 1076 3252 1084
rect 3372 1076 3380 1084
rect 3516 1076 3524 1084
rect 3740 1076 3748 1084
rect 3772 1076 3780 1084
rect 3836 1076 3844 1084
rect 3900 1076 3908 1084
rect 3996 1076 4004 1084
rect 4060 1076 4068 1084
rect 4124 1076 4132 1084
rect 4188 1076 4196 1084
rect 4316 1076 4324 1084
rect 4380 1076 4388 1084
rect 4476 1076 4484 1084
rect 4492 1076 4500 1084
rect 4556 1076 4564 1084
rect 4572 1076 4580 1084
rect 4668 1076 4676 1084
rect 4732 1076 4740 1084
rect 4780 1076 4788 1084
rect 4812 1076 4820 1084
rect 4908 1076 4916 1084
rect 4924 1076 4932 1084
rect 4988 1076 4996 1084
rect 5084 1076 5092 1084
rect 5116 1076 5124 1084
rect 5148 1076 5156 1084
rect 5372 1076 5380 1084
rect 604 1056 612 1064
rect 1004 1056 1012 1064
rect 1292 1056 1300 1064
rect 1324 1056 1332 1064
rect 1340 1056 1348 1064
rect 1404 1056 1412 1064
rect 1436 1056 1444 1064
rect 1468 1056 1476 1064
rect 1596 1056 1604 1064
rect 1612 1056 1620 1064
rect 1740 1056 1748 1064
rect 1772 1056 1780 1064
rect 1964 1056 1972 1064
rect 2140 1056 2148 1064
rect 2332 1056 2340 1064
rect 2364 1056 2372 1064
rect 2396 1056 2404 1064
rect 2412 1056 2420 1064
rect 2668 1056 2676 1064
rect 2908 1056 2916 1064
rect 3212 1056 3220 1064
rect 3548 1056 3556 1064
rect 3836 1056 3844 1064
rect 3932 1056 3940 1064
rect 3964 1056 3972 1064
rect 3980 1056 3988 1064
rect 4044 1056 4052 1064
rect 4236 1056 4244 1064
rect 4332 1056 4340 1064
rect 4636 1056 4644 1064
rect 5340 1056 5348 1064
rect 92 1036 100 1044
rect 396 1036 404 1044
rect 444 1036 452 1044
rect 828 1036 836 1044
rect 1356 1036 1364 1044
rect 2476 1036 2484 1044
rect 2636 1036 2644 1044
rect 3708 1036 3716 1044
rect 4028 1036 4036 1044
rect 4076 1036 4084 1044
rect 4220 1036 4228 1044
rect 4652 1036 4660 1044
rect 4700 1036 4708 1044
rect 4972 1036 4980 1044
rect 5036 1036 5044 1044
rect 2723 1006 2731 1014
rect 2733 1006 2741 1014
rect 2743 1006 2751 1014
rect 2753 1006 2761 1014
rect 2763 1006 2771 1014
rect 2773 1006 2781 1014
rect 140 976 148 984
rect 380 976 388 984
rect 812 976 820 984
rect 1404 976 1412 984
rect 1740 976 1748 984
rect 1836 976 1844 984
rect 2508 976 2516 984
rect 2588 976 2596 984
rect 4092 976 4100 984
rect 4172 976 4180 984
rect 4316 976 4324 984
rect 4540 976 4548 984
rect 4684 976 4692 984
rect 4748 976 4756 984
rect 4828 976 4836 984
rect 5180 976 5188 984
rect 92 956 100 964
rect 620 956 628 964
rect 876 956 884 964
rect 1148 956 1156 964
rect 1372 956 1380 964
rect 1420 956 1428 964
rect 1436 956 1444 964
rect 1852 956 1860 964
rect 1932 956 1940 964
rect 1964 956 1972 964
rect 2124 956 2132 964
rect 2188 956 2196 964
rect 2268 956 2276 964
rect 2284 956 2292 964
rect 2316 956 2324 964
rect 2492 956 2500 964
rect 2604 956 2612 964
rect 2860 956 2868 964
rect 3036 956 3044 964
rect 3068 956 3076 964
rect 3244 956 3252 964
rect 3708 956 3716 964
rect 4156 956 4164 964
rect 4300 956 4308 964
rect 4332 956 4340 964
rect 4988 956 4996 964
rect 5340 956 5348 964
rect 12 936 20 944
rect 236 936 244 944
rect 300 936 308 944
rect 396 936 404 944
rect 428 936 436 944
rect 588 936 596 944
rect 876 936 884 944
rect 908 936 916 944
rect 956 936 964 944
rect 1116 936 1124 944
rect 1452 936 1460 944
rect 1548 936 1556 944
rect 1644 936 1652 944
rect 1932 936 1940 944
rect 2092 936 2100 944
rect 2236 936 2244 944
rect 2316 936 2324 944
rect 2348 936 2356 944
rect 2380 936 2388 944
rect 2444 936 2452 944
rect 2892 936 2900 944
rect 3276 936 3284 944
rect 3420 936 3428 944
rect 3452 936 3460 944
rect 3532 936 3540 944
rect 3676 936 3684 944
rect 3932 936 3940 944
rect 3980 936 3988 944
rect 3996 936 4004 944
rect 4044 936 4052 944
rect 4364 936 4372 944
rect 4460 936 4468 944
rect 4668 936 4676 944
rect 4716 936 4724 944
rect 5020 936 5028 944
rect 5372 936 5380 944
rect 140 916 148 924
rect 204 916 212 924
rect 236 916 244 924
rect 300 916 308 924
rect 412 916 420 924
rect 700 916 708 924
rect 844 916 852 924
rect 908 916 916 924
rect 972 916 980 924
rect 1036 916 1044 924
rect 1500 916 1508 924
rect 1532 916 1540 924
rect 1612 918 1620 926
rect 1756 916 1764 924
rect 1804 916 1812 924
rect 1884 916 1892 924
rect 44 896 52 904
rect 156 896 164 904
rect 220 896 228 904
rect 284 896 292 904
rect 332 896 340 904
rect 380 896 388 904
rect 444 896 452 904
rect 476 896 484 904
rect 812 896 820 904
rect 1052 900 1060 908
rect 1500 896 1508 904
rect 1532 896 1540 904
rect 2076 916 2084 924
rect 1996 896 2004 904
rect 2044 896 2052 904
rect 2124 896 2132 904
rect 2220 916 2228 924
rect 2364 916 2372 924
rect 2460 916 2468 924
rect 2476 916 2484 924
rect 2572 916 2580 924
rect 2780 916 2788 924
rect 3004 916 3012 924
rect 3164 916 3172 924
rect 3436 916 3444 924
rect 2268 896 2276 904
rect 2428 896 2436 904
rect 2988 896 2996 904
rect 3372 896 3380 904
rect 3516 916 3524 924
rect 3676 916 3684 924
rect 3788 916 3796 924
rect 3900 916 3908 924
rect 3484 896 3492 904
rect 3612 900 3620 908
rect 3900 896 3908 904
rect 3932 896 3940 904
rect 4028 896 4036 904
rect 4076 896 4084 904
rect 4124 916 4132 924
rect 4220 916 4228 924
rect 4380 916 4388 924
rect 4412 916 4420 924
rect 4492 916 4500 924
rect 4556 916 4564 924
rect 4620 916 4628 924
rect 4636 916 4644 924
rect 4652 916 4660 924
rect 4716 916 4724 924
rect 4732 916 4740 924
rect 4796 916 4804 924
rect 5116 916 5124 924
rect 5260 916 5268 924
rect 5452 916 5460 924
rect 4396 896 4404 904
rect 4492 896 4500 904
rect 5084 900 5092 908
rect 5436 900 5444 908
rect 124 876 132 884
rect 188 876 196 884
rect 796 876 804 884
rect 2236 876 2244 884
rect 3884 876 3892 884
rect 4412 876 4420 884
rect 700 854 708 862
rect 1052 854 1060 862
rect 3164 854 3172 862
rect 5084 854 5092 862
rect 76 836 84 844
rect 108 836 116 844
rect 204 836 212 844
rect 1788 836 1796 844
rect 1932 836 1940 844
rect 2316 836 2324 844
rect 2988 836 2996 844
rect 3052 836 3060 844
rect 3612 836 3620 844
rect 3916 836 3924 844
rect 3964 836 3972 844
rect 4012 836 4020 844
rect 4188 836 4196 844
rect 4332 836 4340 844
rect 4444 836 4452 844
rect 4476 836 4484 844
rect 4540 836 4548 844
rect 4604 836 4612 844
rect 5436 836 5444 844
rect 1219 806 1227 814
rect 1229 806 1237 814
rect 1239 806 1247 814
rect 1249 806 1257 814
rect 1259 806 1267 814
rect 1269 806 1277 814
rect 4227 806 4235 814
rect 4237 806 4245 814
rect 4247 806 4255 814
rect 4257 806 4265 814
rect 4267 806 4275 814
rect 4277 806 4285 814
rect 28 776 36 784
rect 156 776 164 784
rect 236 776 244 784
rect 268 776 276 784
rect 652 776 660 784
rect 828 776 836 784
rect 876 776 884 784
rect 1212 776 1220 784
rect 1340 776 1348 784
rect 1756 776 1764 784
rect 2044 776 2052 784
rect 2092 776 2100 784
rect 4108 776 4116 784
rect 4172 776 4180 784
rect 4460 776 4468 784
rect 4572 776 4580 784
rect 5020 776 5028 784
rect 5452 776 5460 784
rect 1532 756 1540 764
rect 2348 758 2356 766
rect 2940 756 2948 764
rect 3340 756 3348 764
rect 3644 758 3652 766
rect 812 736 820 744
rect 860 736 868 744
rect 1676 736 1684 744
rect 364 716 372 724
rect 396 716 404 724
rect 44 696 52 704
rect 92 696 100 704
rect 124 696 132 704
rect 220 696 228 704
rect 268 696 276 704
rect 316 696 324 704
rect 460 696 468 704
rect 492 696 500 704
rect 540 696 548 704
rect 588 716 596 724
rect 1212 716 1220 724
rect 1628 716 1636 724
rect 1756 716 1764 724
rect 2348 712 2356 720
rect 764 696 772 704
rect 796 696 804 704
rect 876 696 884 704
rect 1196 696 1204 704
rect 1532 696 1540 704
rect 1708 696 1716 704
rect 1772 696 1780 704
rect 1964 696 1972 704
rect 2172 696 2180 704
rect 2396 696 2404 704
rect 2460 696 2468 704
rect 2524 696 2532 704
rect 2572 716 2580 724
rect 3036 716 3044 724
rect 2604 696 2612 704
rect 2732 696 2740 704
rect 2940 696 2948 704
rect 3100 696 3108 704
rect 3148 716 3156 724
rect 3644 712 3652 720
rect 3772 716 3780 724
rect 3916 716 3924 724
rect 3948 716 3956 724
rect 4460 716 4468 724
rect 4508 716 4516 724
rect 4668 716 4676 724
rect 4908 716 4916 724
rect 4972 716 4980 724
rect 4988 716 4996 724
rect 5052 716 5060 724
rect 5084 716 5092 724
rect 5452 716 5460 724
rect 3180 696 3188 704
rect 3212 696 3220 704
rect 3276 696 3284 704
rect 3308 696 3316 704
rect 3676 696 3684 704
rect 3740 696 3748 704
rect 3756 696 3764 704
rect 3804 696 3812 704
rect 3852 696 3860 704
rect 3884 696 3892 704
rect 4012 696 4020 704
rect 4460 696 4468 704
rect 4556 696 4564 704
rect 4668 696 4676 704
rect 4764 696 4772 704
rect 4780 696 4788 704
rect 4844 696 4852 704
rect 4876 696 4884 704
rect 4924 696 4932 704
rect 4940 696 4948 704
rect 5020 696 5028 704
rect 5420 696 5428 704
rect 140 676 148 684
rect 300 676 308 684
rect 396 676 404 684
rect 444 676 452 684
rect 508 676 516 684
rect 524 676 532 684
rect 556 676 564 684
rect 620 676 628 684
rect 764 676 772 684
rect 1116 676 1124 684
rect 1532 676 1540 684
rect 1852 676 1860 684
rect 2284 676 2292 684
rect 2620 676 2628 684
rect 2940 676 2948 684
rect 3084 676 3092 684
rect 3116 676 3124 684
rect 3196 676 3204 684
rect 3260 676 3268 684
rect 3580 676 3588 684
rect 3724 676 3732 684
rect 3788 676 3796 684
rect 3868 676 3876 684
rect 3932 676 3940 684
rect 3996 676 4004 684
rect 4364 676 4372 684
rect 4588 676 4596 684
rect 4652 676 4660 684
rect 4748 676 4756 684
rect 4876 676 4884 684
rect 4908 676 4916 684
rect 5036 676 5044 684
rect 5100 676 5108 684
rect 5148 676 5156 684
rect 5162 676 5170 684
rect 5356 676 5364 684
rect 12 656 20 664
rect 28 656 36 664
rect 60 656 68 664
rect 92 656 100 664
rect 172 656 180 664
rect 188 656 196 664
rect 252 656 260 664
rect 300 656 308 664
rect 348 656 356 664
rect 428 656 436 664
rect 1084 656 1092 664
rect 1500 656 1508 664
rect 1884 656 1892 664
rect 2252 656 2260 664
rect 2428 656 2436 664
rect 2476 656 2484 664
rect 2636 656 2644 664
rect 2668 656 2676 664
rect 2908 656 2916 664
rect 3244 656 3252 664
rect 3548 656 3556 664
rect 3948 656 3956 664
rect 3980 656 3988 664
rect 4044 656 4052 664
rect 4060 656 4068 664
rect 4332 656 4340 664
rect 4588 656 4596 664
rect 4604 656 4612 664
rect 4684 656 4692 664
rect 4716 656 4724 664
rect 4828 656 4836 664
rect 5324 656 5332 664
rect 364 636 372 644
rect 492 636 500 644
rect 924 636 932 644
rect 2556 636 2564 644
rect 3276 636 3284 644
rect 3804 636 3812 644
rect 3916 636 3924 644
rect 4028 636 4036 644
rect 4508 636 4516 644
rect 4972 636 4980 644
rect 5052 636 5060 644
rect 5116 636 5124 644
rect 2723 606 2731 614
rect 2733 606 2741 614
rect 2743 606 2751 614
rect 2753 606 2761 614
rect 2763 606 2771 614
rect 2773 606 2781 614
rect 76 576 84 584
rect 156 576 164 584
rect 348 576 356 584
rect 380 576 388 584
rect 876 576 884 584
rect 1340 576 1348 584
rect 1596 576 1604 584
rect 1692 576 1700 584
rect 3132 576 3140 584
rect 3676 576 3684 584
rect 4060 576 4068 584
rect 4428 576 4436 584
rect 5148 576 5156 584
rect 12 556 20 564
rect 92 556 100 564
rect 396 556 404 564
rect 572 556 580 564
rect 748 556 756 564
rect 1068 556 1076 564
rect 1324 556 1332 564
rect 1356 556 1364 564
rect 1388 556 1396 564
rect 1548 556 1556 564
rect 1660 556 1668 564
rect 1708 556 1716 564
rect 1932 556 1940 564
rect 2268 556 2276 564
rect 2348 556 2356 564
rect 2524 556 2532 564
rect 2972 556 2980 564
rect 3164 556 3172 564
rect 3356 556 3364 564
rect 3548 556 3556 564
rect 3580 556 3588 564
rect 3596 556 3604 564
rect 3900 556 3908 564
rect 4204 556 4212 564
rect 4588 556 4596 564
rect 5308 556 5316 564
rect 44 536 52 544
rect 108 536 116 544
rect 124 536 132 544
rect 172 536 180 544
rect 236 536 244 544
rect 252 536 260 544
rect 316 536 324 544
rect 332 536 340 544
rect 540 536 548 544
rect 764 536 772 544
rect 1036 536 1044 544
rect 1484 536 1492 544
rect 1628 536 1636 544
rect 1740 536 1748 544
rect 1900 536 1908 544
rect 2124 536 2132 544
rect 2236 536 2244 544
rect 2556 536 2564 544
rect 2940 536 2948 544
rect 3180 536 3188 544
rect 3324 536 3332 544
rect 3724 536 3732 544
rect 3868 536 3876 544
rect 4092 536 4100 544
rect 4300 536 4308 544
rect 4380 536 4388 544
rect 4620 536 4628 544
rect 4764 536 4772 544
rect 188 516 196 524
rect 220 516 228 524
rect 268 516 276 524
rect 300 516 308 524
rect 460 516 468 524
rect 1148 516 1156 524
rect 1230 516 1238 524
rect 1356 516 1364 524
rect 1484 516 1492 524
rect 44 496 52 504
rect 156 496 164 504
rect 476 500 484 508
rect 940 496 948 504
rect 1452 496 1460 504
rect 1580 516 1588 524
rect 1628 516 1636 524
rect 1660 516 1668 524
rect 2012 516 2020 524
rect 2140 516 2148 524
rect 2156 516 2164 524
rect 1596 496 1604 504
rect 1804 496 1812 504
rect 2220 516 2228 524
rect 2300 516 2308 524
rect 2362 516 2370 524
rect 2444 516 2452 524
rect 2700 516 2708 524
rect 3052 516 3060 524
rect 3212 516 3220 524
rect 3436 516 3444 524
rect 3548 516 3556 524
rect 3580 516 3588 524
rect 3644 516 3652 524
rect 2188 496 2196 504
rect 2332 496 2340 504
rect 2620 500 2628 508
rect 2844 496 2852 504
rect 3260 500 3268 508
rect 3772 516 3780 524
rect 4108 516 4116 524
rect 4156 516 4164 524
rect 4172 516 4180 524
rect 4252 516 4260 524
rect 4348 516 4356 524
rect 4364 516 4372 524
rect 4508 516 4516 524
rect 4732 516 4740 524
rect 4828 516 4836 524
rect 4844 516 4852 524
rect 4876 516 4884 524
rect 4892 516 4900 524
rect 4924 516 4932 524
rect 4972 516 4980 524
rect 5004 536 5012 544
rect 5036 536 5044 544
rect 5068 536 5076 544
rect 5116 536 5124 544
rect 5340 536 5348 544
rect 5084 516 5092 524
rect 5340 516 5348 524
rect 5420 516 5428 524
rect 3692 496 3700 504
rect 3804 500 3812 508
rect 4684 500 4692 508
rect 4796 496 4804 504
rect 5052 496 5060 504
rect 5132 496 5140 504
rect 5404 500 5412 508
rect 2108 476 2116 484
rect 2268 476 2276 484
rect 4188 476 4196 484
rect 1148 454 1156 462
rect 2012 454 2020 462
rect 2444 454 2452 462
rect 3052 454 3060 462
rect 3260 454 3268 462
rect 3804 454 3812 462
rect 4684 454 4692 462
rect 5404 454 5412 462
rect 204 436 212 444
rect 268 436 276 444
rect 476 436 484 444
rect 1420 436 1428 444
rect 2796 436 2804 444
rect 4780 436 4788 444
rect 1219 406 1227 414
rect 1229 406 1237 414
rect 1239 406 1247 414
rect 1249 406 1257 414
rect 1259 406 1267 414
rect 1269 406 1277 414
rect 4227 406 4235 414
rect 4237 406 4245 414
rect 4247 406 4255 414
rect 4257 406 4265 414
rect 4267 406 4275 414
rect 4277 406 4285 414
rect 28 376 36 384
rect 316 376 324 384
rect 380 376 388 384
rect 668 376 676 384
rect 1340 376 1348 384
rect 1692 376 1700 384
rect 2252 376 2260 384
rect 3756 376 3764 384
rect 4044 376 4052 384
rect 4140 376 4148 384
rect 4204 376 4212 384
rect 4492 376 4500 384
rect 4828 376 4836 384
rect 5196 376 5204 384
rect 5308 376 5316 384
rect 5468 376 5476 384
rect 972 358 980 366
rect 1532 356 1540 364
rect 1884 356 1892 364
rect 2508 356 2516 364
rect 3084 356 3092 364
rect 3500 358 3508 366
rect 5084 358 5092 366
rect 2140 336 2148 344
rect 316 316 324 324
rect 668 316 676 324
rect 972 312 980 320
rect 1628 316 1636 324
rect 1948 312 1956 320
rect 316 296 324 304
rect 460 296 468 304
rect 668 296 676 304
rect 748 296 756 304
rect 940 296 948 304
rect 1148 296 1156 304
rect 1532 296 1540 304
rect 1884 296 1892 304
rect 2076 316 2084 324
rect 2188 316 2196 324
rect 2220 316 2228 324
rect 2300 316 2308 324
rect 2620 316 2628 324
rect 2108 296 2116 304
rect 2140 296 2148 304
rect 2220 296 2228 304
rect 2508 296 2516 304
rect 2700 296 2708 304
rect 2812 316 2820 324
rect 3148 312 3156 320
rect 3500 312 3508 320
rect 3756 316 3764 324
rect 4204 316 4212 324
rect 4796 316 4804 324
rect 5084 312 5092 320
rect 2876 296 2884 304
rect 3084 296 3092 304
rect 3242 296 3250 304
rect 3436 296 3444 304
rect 3772 296 3780 304
rect 3964 296 3972 304
rect 4204 296 4212 304
rect 4588 296 4596 304
rect 4652 294 4660 302
rect 4764 296 4772 304
rect 4908 296 4916 304
rect 5100 296 5108 304
rect 5180 296 5188 304
rect 5228 296 5236 304
rect 5244 296 5252 304
rect 5276 296 5284 304
rect 5324 296 5332 304
rect 220 276 228 284
rect 572 276 580 284
rect 764 276 772 284
rect 1036 276 1044 284
rect 1532 276 1540 284
rect 1884 276 1892 284
rect 2028 276 2036 284
rect 2044 276 2052 284
rect 2124 276 2132 284
rect 2172 276 2180 284
rect 2236 276 2244 284
rect 2508 276 2516 284
rect 2716 276 2724 284
rect 2860 276 2868 284
rect 3084 276 3092 284
rect 3436 276 3444 284
rect 3708 276 3716 284
rect 3852 276 3860 284
rect 4300 276 4308 284
rect 4684 276 4692 284
rect 5020 276 5028 284
rect 5356 276 5364 284
rect 188 256 196 264
rect 540 256 548 264
rect 1068 256 1076 264
rect 1500 256 1508 264
rect 1852 256 1860 264
rect 2140 256 2148 264
rect 2476 256 2484 264
rect 2652 256 2660 264
rect 3052 256 3060 264
rect 3404 256 3412 264
rect 3884 256 3892 264
rect 4076 256 4084 264
rect 4332 256 4340 264
rect 4588 256 4596 264
rect 4716 256 4724 264
rect 4988 256 4996 264
rect 716 236 724 244
rect 876 236 884 244
rect 1228 236 1236 244
rect 1756 236 1764 244
rect 2316 236 2324 244
rect 2668 236 2676 244
rect 2892 236 2900 244
rect 3596 236 3604 244
rect 4796 236 4804 244
rect 2723 206 2731 214
rect 2733 206 2741 214
rect 2743 206 2751 214
rect 2753 206 2761 214
rect 2763 206 2771 214
rect 2773 206 2781 214
rect 28 176 36 184
rect 1212 176 1220 184
rect 2140 176 2148 184
rect 2348 176 2356 184
rect 2876 176 2884 184
rect 3356 176 3364 184
rect 4284 176 4292 184
rect 4988 176 4996 184
rect 5036 176 5044 184
rect 188 156 196 164
rect 524 156 532 164
rect 1004 156 1012 164
rect 1196 156 1204 164
rect 1548 156 1556 164
rect 1980 156 1988 164
rect 2652 156 2660 164
rect 2668 156 2676 164
rect 3068 156 3076 164
rect 3548 156 3556 164
rect 4124 156 4132 164
rect 4828 156 4836 164
rect 5020 156 5028 164
rect 5212 156 5220 164
rect 220 136 228 144
rect 492 136 500 144
rect 780 136 788 144
rect 972 136 980 144
rect 1356 136 1364 144
rect 1580 136 1588 144
rect 1948 136 1956 144
rect 2172 136 2180 144
rect 2236 136 2244 144
rect 2268 136 2276 144
rect 2332 136 2340 144
rect 2380 136 2388 144
rect 2444 136 2452 144
rect 2556 136 2564 144
rect 2620 136 2628 144
rect 2636 136 2644 144
rect 2684 136 2692 144
rect 2700 136 2708 144
rect 2780 136 2788 144
rect 2796 136 2804 144
rect 3100 136 3108 144
rect 3244 136 3252 144
rect 3308 136 3316 144
rect 3580 136 3588 144
rect 3868 136 3876 144
rect 4092 136 4100 144
rect 4796 136 4804 144
rect 5180 136 5188 144
rect 316 116 324 124
rect 604 116 612 124
rect 686 116 694 124
rect 700 116 708 124
rect 748 116 756 124
rect 796 116 804 124
rect 828 116 836 124
rect 908 116 916 124
rect 1166 116 1174 124
rect 1660 116 1668 124
rect 1756 116 1764 124
rect 2060 116 2068 124
rect 2220 116 2228 124
rect 2252 116 2260 124
rect 2396 116 2404 124
rect 2460 116 2468 124
rect 316 96 324 104
rect 428 100 436 108
rect 876 96 884 104
rect 1308 96 1316 104
rect 1644 100 1652 108
rect 1852 96 1860 104
rect 2252 96 2260 104
rect 2316 96 2324 104
rect 2364 96 2372 104
rect 2428 96 2436 104
rect 2492 96 2500 104
rect 2540 116 2548 124
rect 2556 116 2564 124
rect 2620 116 2628 124
rect 2716 116 2724 124
rect 2812 116 2820 124
rect 2906 116 2914 124
rect 2988 116 2996 124
rect 3260 116 3268 124
rect 3292 116 3300 124
rect 3324 116 3332 124
rect 3676 116 3684 124
rect 3900 118 3908 126
rect 3996 116 4004 124
rect 4204 116 4212 124
rect 4428 118 4436 126
rect 4492 116 4500 124
rect 4620 116 4628 124
rect 4732 116 4740 124
rect 4908 116 4916 124
rect 5100 116 5108 124
rect 5452 116 5460 124
rect 2572 96 2580 104
rect 2652 96 2660 104
rect 2748 96 2756 104
rect 2876 96 2884 104
rect 3212 96 3220 104
rect 3388 96 3396 104
rect 3644 100 3652 108
rect 3996 96 4004 104
rect 4700 96 4708 104
rect 5084 96 5092 104
rect 2284 76 2292 84
rect 2396 76 2404 84
rect 2540 76 2548 84
rect 5516 76 5524 84
rect 2060 54 2068 62
rect 2988 54 2996 62
rect 3644 54 3652 62
rect 316 36 324 44
rect 428 36 436 44
rect 876 36 884 44
rect 1644 36 1652 44
rect 1724 36 1732 44
rect 1804 36 1812 44
rect 3724 36 3732 44
rect 3996 36 4004 44
rect 4604 36 4612 44
rect 4652 36 4660 44
rect 4700 36 4708 44
rect 5084 36 5092 44
rect 5436 36 5444 44
rect 1219 6 1227 14
rect 1229 6 1237 14
rect 1239 6 1247 14
rect 1249 6 1257 14
rect 1259 6 1267 14
rect 1269 6 1277 14
rect 4227 6 4235 14
rect 4237 6 4245 14
rect 4247 6 4255 14
rect 4257 6 4265 14
rect 4267 6 4275 14
rect 4277 6 4285 14
<< metal2 >>
rect 2061 3824 2067 3863
rect 3405 3824 3411 3863
rect 2746 3814 2758 3816
rect 2731 3806 2733 3814
rect 2741 3806 2743 3814
rect 2751 3806 2753 3814
rect 2761 3806 2763 3814
rect 2771 3806 2773 3814
rect 2746 3804 2758 3806
rect 3437 3804 3443 3863
rect 13 3364 19 3676
rect 189 3464 195 3756
rect 285 3504 291 3716
rect 317 3644 323 3696
rect 429 3644 435 3700
rect 493 3643 499 3736
rect 493 3637 515 3643
rect 317 3524 323 3576
rect 189 3404 195 3456
rect 221 3364 227 3396
rect 13 3124 19 3356
rect 253 3304 259 3336
rect 317 3324 323 3496
rect 381 3464 387 3576
rect 429 3464 435 3516
rect 445 3504 451 3576
rect 397 3344 403 3436
rect 29 3184 35 3236
rect 13 3104 19 3116
rect 45 3064 51 3276
rect 349 3244 355 3296
rect 301 3184 307 3216
rect 173 3144 179 3176
rect 253 3124 259 3176
rect 276 3117 291 3123
rect 13 2564 19 3056
rect 29 2784 35 2896
rect 45 2883 51 2916
rect 77 2883 83 3096
rect 221 3084 227 3116
rect 221 3064 227 3076
rect 189 2984 195 3036
rect 109 2924 115 2956
rect 141 2924 147 2956
rect 237 2924 243 3096
rect 285 2984 291 3117
rect 301 3084 307 3096
rect 317 3084 323 3176
rect 333 3044 339 3056
rect 333 2964 339 2976
rect 365 2964 371 3096
rect 381 3064 387 3136
rect 397 3043 403 3336
rect 413 3324 419 3436
rect 445 3384 451 3476
rect 477 3464 483 3516
rect 493 3464 499 3576
rect 461 3344 467 3436
rect 509 3424 515 3637
rect 541 3484 547 3516
rect 525 3404 531 3456
rect 573 3384 579 3516
rect 605 3504 611 3716
rect 733 3584 739 3676
rect 653 3520 659 3558
rect 493 3344 499 3356
rect 621 3337 636 3343
rect 525 3324 531 3336
rect 429 3284 435 3296
rect 445 3184 451 3296
rect 477 3264 483 3316
rect 573 3304 579 3316
rect 589 3304 595 3316
rect 589 3283 595 3296
rect 573 3277 595 3283
rect 541 3164 547 3276
rect 573 3184 579 3277
rect 605 3164 611 3276
rect 381 3037 403 3043
rect 141 2904 147 2916
rect 221 2904 227 2916
rect 45 2877 83 2883
rect 45 2564 51 2836
rect 45 2243 51 2296
rect 36 2237 51 2243
rect 45 2144 51 2237
rect 61 2224 67 2877
rect 189 2664 195 2816
rect 237 2784 243 2836
rect 221 2684 227 2736
rect 285 2724 291 2896
rect 301 2704 307 2756
rect 317 2724 323 2776
rect 93 2544 99 2556
rect 141 2544 147 2556
rect 125 2504 131 2516
rect 189 2464 195 2656
rect 237 2564 243 2576
rect 205 2524 211 2536
rect 61 2164 67 2216
rect 77 2164 83 2436
rect 189 2284 195 2436
rect 221 2284 227 2316
rect 285 2304 291 2696
rect 301 2584 307 2676
rect 317 2544 323 2556
rect 221 2223 227 2256
rect 301 2244 307 2436
rect 317 2324 323 2376
rect 205 2217 227 2223
rect 61 2124 67 2156
rect 173 2144 179 2156
rect 93 2124 99 2136
rect 125 2084 131 2136
rect 13 1764 19 1876
rect 29 1524 35 2036
rect 45 1904 51 1916
rect 109 1904 115 1916
rect 45 1764 51 1836
rect 61 1703 67 1896
rect 93 1864 99 1876
rect 77 1764 83 1836
rect 109 1764 115 1896
rect 125 1764 131 2076
rect 109 1717 124 1723
rect 61 1697 83 1703
rect 45 1504 51 1576
rect 77 1544 83 1697
rect 13 1484 19 1496
rect 77 1384 83 1436
rect 29 1344 35 1376
rect 45 1324 51 1356
rect 77 1304 83 1356
rect 109 1303 115 1717
rect 157 1723 163 2136
rect 205 2103 211 2217
rect 221 2144 227 2196
rect 269 2124 275 2156
rect 285 2104 291 2196
rect 301 2144 307 2156
rect 196 2097 211 2103
rect 269 2064 275 2096
rect 301 2084 307 2136
rect 317 2124 323 2196
rect 333 2004 339 2936
rect 365 2924 371 2956
rect 381 2924 387 3037
rect 397 2984 403 3016
rect 413 2964 419 3096
rect 429 3084 435 3116
rect 445 3104 451 3116
rect 477 3104 483 3156
rect 445 3084 451 3096
rect 349 2683 355 2876
rect 365 2724 371 2836
rect 349 2677 364 2683
rect 365 2544 371 2656
rect 365 2504 371 2536
rect 381 2524 387 2676
rect 365 2463 371 2496
rect 381 2484 387 2516
rect 349 2457 371 2463
rect 349 2124 355 2457
rect 381 2364 387 2476
rect 397 2464 403 2836
rect 413 2624 419 2696
rect 429 2684 435 2996
rect 445 2864 451 3076
rect 493 3004 499 3076
rect 509 3064 515 3076
rect 541 3044 547 3116
rect 557 3104 563 3116
rect 573 3104 579 3136
rect 621 3104 627 3337
rect 637 3184 643 3296
rect 653 3124 659 3276
rect 685 3184 691 3416
rect 653 3104 659 3116
rect 669 3104 675 3116
rect 573 3004 579 3036
rect 477 2764 483 2916
rect 557 2824 563 2956
rect 589 2944 595 3096
rect 621 3024 627 3076
rect 653 3044 659 3096
rect 669 3064 675 3076
rect 653 2862 659 2900
rect 669 2784 675 3016
rect 701 2944 707 3296
rect 717 3224 723 3476
rect 749 3444 755 3456
rect 893 3444 899 3756
rect 989 3662 995 3700
rect 925 3504 931 3656
rect 733 3344 739 3376
rect 925 3364 931 3496
rect 973 3464 979 3576
rect 1005 3504 1011 3716
rect 1309 3643 1315 3756
rect 1341 3744 1347 3756
rect 1613 3724 1619 3736
rect 1293 3637 1315 3643
rect 1242 3614 1254 3616
rect 1227 3606 1229 3614
rect 1237 3606 1239 3614
rect 1247 3606 1249 3614
rect 1257 3606 1259 3614
rect 1267 3606 1269 3614
rect 1242 3604 1254 3606
rect 1053 3520 1059 3558
rect 797 3344 803 3356
rect 893 3304 899 3336
rect 861 3284 867 3296
rect 941 3284 947 3456
rect 957 3384 963 3436
rect 973 3344 979 3456
rect 1149 3424 1155 3456
rect 1117 3364 1123 3416
rect 1149 3304 1155 3336
rect 1229 3324 1235 3496
rect 1293 3424 1299 3637
rect 1405 3504 1411 3716
rect 1437 3644 1443 3696
rect 1437 3524 1443 3576
rect 1533 3504 1539 3716
rect 1549 3644 1555 3700
rect 717 3024 723 3096
rect 733 3084 739 3136
rect 877 3064 883 3236
rect 925 3104 931 3256
rect 957 3124 963 3236
rect 749 3044 755 3056
rect 429 2584 435 2676
rect 445 2664 451 2716
rect 477 2684 483 2716
rect 797 2704 803 3056
rect 909 2964 915 3076
rect 925 3064 931 3076
rect 493 2684 499 2696
rect 637 2684 643 2696
rect 525 2644 531 2656
rect 461 2564 467 2636
rect 397 2384 403 2436
rect 413 2384 419 2456
rect 365 2304 371 2316
rect 381 2304 387 2336
rect 381 2164 387 2296
rect 397 2284 403 2336
rect 429 2284 435 2536
rect 461 2484 467 2496
rect 477 2464 483 2496
rect 493 2424 499 2516
rect 509 2484 515 2496
rect 557 2443 563 2656
rect 573 2584 579 2636
rect 573 2464 579 2496
rect 557 2437 579 2443
rect 397 2144 403 2236
rect 429 2224 435 2276
rect 445 2124 451 2296
rect 461 2124 467 2416
rect 493 2284 499 2396
rect 525 2364 531 2436
rect 509 2304 515 2356
rect 381 2104 387 2116
rect 381 2044 387 2096
rect 148 1717 163 1723
rect 141 1524 147 1716
rect 173 1504 179 1876
rect 205 1804 211 1836
rect 253 1803 259 1896
rect 269 1864 275 1876
rect 285 1824 291 1876
rect 237 1797 259 1803
rect 237 1784 243 1797
rect 237 1764 243 1776
rect 189 1723 195 1756
rect 285 1724 291 1796
rect 189 1717 211 1723
rect 189 1504 195 1516
rect 205 1484 211 1717
rect 301 1704 307 1736
rect 317 1684 323 1936
rect 333 1863 339 1916
rect 349 1904 355 1916
rect 333 1857 355 1863
rect 205 1464 211 1476
rect 253 1464 259 1536
rect 205 1423 211 1436
rect 285 1424 291 1456
rect 205 1417 227 1423
rect 125 1364 131 1416
rect 157 1324 163 1356
rect 205 1344 211 1396
rect 173 1324 179 1336
rect 189 1324 195 1336
rect 221 1304 227 1417
rect 285 1304 291 1316
rect 93 1297 115 1303
rect 13 944 19 1236
rect 45 1184 51 1216
rect 93 1184 99 1297
rect 221 1284 227 1296
rect 221 1184 227 1256
rect 301 1243 307 1676
rect 349 1644 355 1857
rect 365 1784 371 1936
rect 365 1744 371 1776
rect 381 1744 387 1756
rect 397 1724 403 2116
rect 477 2104 483 2116
rect 429 2077 444 2083
rect 429 2064 435 2077
rect 413 1944 419 2036
rect 429 1984 435 2016
rect 445 1924 451 2056
rect 461 2044 467 2096
rect 413 1897 428 1903
rect 381 1717 396 1723
rect 365 1504 371 1516
rect 317 1464 323 1496
rect 333 1384 339 1456
rect 365 1364 371 1456
rect 365 1344 371 1356
rect 333 1324 339 1336
rect 381 1324 387 1717
rect 413 1664 419 1897
rect 461 1864 467 2036
rect 493 2003 499 2276
rect 557 2204 563 2236
rect 573 2184 579 2437
rect 589 2304 595 2456
rect 605 2344 611 2676
rect 621 2624 627 2636
rect 685 2524 691 2656
rect 701 2544 707 2636
rect 733 2544 739 2576
rect 749 2564 755 2656
rect 765 2564 771 2656
rect 829 2563 835 2696
rect 861 2684 867 2696
rect 820 2557 835 2563
rect 669 2503 675 2516
rect 669 2497 684 2503
rect 621 2324 627 2456
rect 653 2444 659 2476
rect 653 2304 659 2436
rect 701 2304 707 2376
rect 717 2344 723 2516
rect 733 2404 739 2536
rect 749 2403 755 2536
rect 749 2397 771 2403
rect 605 2284 611 2296
rect 653 2284 659 2296
rect 733 2284 739 2336
rect 749 2304 755 2376
rect 509 2024 515 2156
rect 525 2104 531 2136
rect 637 2124 643 2136
rect 477 1997 499 2003
rect 477 1864 483 1997
rect 541 1964 547 2116
rect 621 2084 627 2096
rect 637 2064 643 2116
rect 653 2084 659 2176
rect 637 2024 643 2036
rect 525 1924 531 1936
rect 493 1884 499 1896
rect 445 1744 451 1856
rect 429 1724 435 1736
rect 429 1584 435 1676
rect 445 1624 451 1736
rect 461 1724 467 1736
rect 365 1317 380 1323
rect 349 1304 355 1316
rect 333 1264 339 1276
rect 285 1237 307 1243
rect 205 1144 211 1156
rect 61 1124 67 1136
rect 29 1097 44 1103
rect 13 904 19 936
rect 29 784 35 1097
rect 45 1084 51 1096
rect 45 884 51 896
rect 13 564 19 656
rect 45 564 51 696
rect 61 684 67 1116
rect 93 964 99 1036
rect 141 984 147 1096
rect 141 924 147 956
rect 157 944 163 1096
rect 77 744 83 836
rect 61 664 67 676
rect 77 657 92 663
rect 77 584 83 657
rect 109 584 115 836
rect 141 684 147 916
rect 173 904 179 1116
rect 189 884 195 1136
rect 269 1124 275 1236
rect 285 1144 291 1237
rect 301 1184 307 1216
rect 237 1003 243 1116
rect 365 1104 371 1317
rect 237 997 259 1003
rect 237 944 243 956
rect 237 904 243 916
rect 205 844 211 876
rect 157 784 163 816
rect 157 657 172 663
rect 157 584 163 657
rect 205 564 211 836
rect 237 784 243 896
rect 253 884 259 997
rect 269 924 275 1096
rect 333 1064 339 1076
rect 269 784 275 916
rect 285 904 291 976
rect 301 884 307 916
rect 317 704 323 1016
rect 333 904 339 976
rect 365 724 371 1076
rect 381 984 387 1296
rect 413 1284 419 1296
rect 397 964 403 1036
rect 429 944 435 1556
rect 445 1524 451 1536
rect 445 1304 451 1476
rect 477 1343 483 1836
rect 493 1784 499 1856
rect 557 1824 563 1936
rect 573 1864 579 1896
rect 605 1884 611 2016
rect 621 1904 627 1996
rect 525 1784 531 1816
rect 541 1744 547 1796
rect 493 1464 499 1596
rect 509 1504 515 1536
rect 461 1337 483 1343
rect 461 1324 467 1337
rect 493 1284 499 1436
rect 509 1384 515 1456
rect 445 1024 451 1036
rect 461 984 467 1236
rect 525 1084 531 1516
rect 573 1484 579 1616
rect 589 1504 595 1636
rect 605 1544 611 1876
rect 621 1484 627 1896
rect 637 1564 643 1996
rect 669 1924 675 2236
rect 685 2104 691 2176
rect 765 2124 771 2397
rect 797 2304 803 2516
rect 829 2284 835 2316
rect 845 2304 851 2336
rect 861 2264 867 2296
rect 797 2244 803 2256
rect 701 2004 707 2116
rect 717 2084 723 2096
rect 749 2044 755 2096
rect 781 2084 787 2176
rect 813 2104 819 2236
rect 861 2184 867 2236
rect 733 2004 739 2036
rect 829 1984 835 2136
rect 877 2124 883 2336
rect 893 2304 899 2636
rect 909 2604 915 2956
rect 941 2944 947 3116
rect 989 3104 995 3116
rect 1037 3084 1043 3296
rect 1005 2844 1011 2900
rect 1021 2844 1027 3076
rect 1069 2963 1075 3216
rect 1085 3064 1091 3116
rect 1117 3064 1123 3276
rect 1213 3262 1219 3300
rect 1242 3214 1254 3216
rect 1227 3206 1229 3214
rect 1237 3206 1239 3214
rect 1247 3206 1249 3214
rect 1257 3206 1259 3214
rect 1267 3206 1269 3214
rect 1242 3204 1254 3206
rect 1085 2984 1091 3056
rect 1069 2957 1084 2963
rect 1181 2944 1187 3056
rect 1197 3004 1203 3076
rect 1197 2964 1203 2976
rect 1229 2924 1235 3056
rect 1261 2924 1267 3036
rect 1293 2944 1299 3116
rect 1309 3044 1315 3436
rect 1405 3324 1411 3496
rect 1517 3364 1523 3416
rect 1533 3404 1539 3476
rect 1565 3424 1571 3456
rect 1645 3424 1651 3756
rect 1965 3744 1971 3776
rect 1725 3704 1731 3716
rect 1405 3184 1411 3296
rect 1421 3244 1427 3300
rect 1485 3184 1491 3336
rect 1517 3224 1523 3356
rect 1597 3324 1603 3336
rect 1565 3184 1571 3216
rect 1677 3204 1683 3236
rect 1341 3004 1347 3136
rect 1405 3104 1411 3136
rect 1357 3044 1363 3056
rect 1357 2963 1363 3036
rect 1357 2957 1372 2963
rect 1437 2944 1443 3116
rect 1597 3104 1603 3196
rect 1565 2964 1571 3036
rect 1597 2944 1603 3096
rect 1613 3064 1619 3076
rect 1629 3057 1644 3063
rect 1533 2924 1539 2936
rect 1613 2923 1619 3056
rect 1629 2984 1635 3057
rect 1661 2984 1667 3116
rect 1677 3104 1683 3176
rect 1709 3104 1715 3476
rect 1725 3184 1731 3436
rect 1757 3384 1763 3716
rect 1869 3704 1875 3716
rect 1773 3404 1779 3436
rect 1821 3364 1827 3676
rect 1901 3644 1907 3700
rect 1997 3624 2003 3756
rect 2285 3724 2291 3736
rect 2349 3724 2355 3736
rect 2269 3704 2275 3716
rect 2333 3704 2339 3716
rect 2397 3703 2403 3736
rect 2461 3724 2467 3736
rect 2445 3704 2451 3716
rect 2397 3697 2419 3703
rect 1933 3464 1939 3616
rect 2029 3520 2035 3558
rect 2157 3524 2163 3696
rect 2189 3644 2195 3696
rect 2365 3684 2371 3696
rect 2397 3664 2403 3676
rect 2413 3664 2419 3697
rect 2509 3684 2515 3696
rect 2461 3584 2467 3636
rect 2525 3584 2531 3656
rect 2541 3584 2547 3636
rect 2381 3520 2387 3558
rect 1933 3424 1939 3456
rect 1965 3424 1971 3476
rect 1917 3364 1923 3396
rect 1997 3384 2003 3416
rect 2093 3384 2099 3496
rect 2132 3437 2147 3443
rect 1757 3104 1763 3136
rect 1693 2964 1699 3016
rect 1604 2917 1619 2923
rect 1661 2917 1676 2923
rect 973 2720 979 2758
rect 1037 2704 1043 2916
rect 1229 2904 1235 2916
rect 1140 2897 1155 2903
rect 1085 2844 1091 2896
rect 1149 2724 1155 2897
rect 1242 2814 1254 2816
rect 1227 2806 1229 2814
rect 1237 2806 1239 2814
rect 1247 2806 1249 2814
rect 1257 2806 1259 2814
rect 1267 2806 1269 2814
rect 1242 2804 1254 2806
rect 1325 2704 1331 2896
rect 1357 2844 1363 2896
rect 1341 2784 1347 2836
rect 1453 2764 1459 2896
rect 1501 2744 1507 2836
rect 1037 2644 1043 2676
rect 1069 2604 1075 2656
rect 973 2564 979 2596
rect 1005 2524 1011 2536
rect 1069 2462 1075 2500
rect 1101 2484 1107 2516
rect 1149 2484 1155 2696
rect 925 2144 931 2296
rect 1005 2284 1011 2356
rect 1021 2304 1027 2376
rect 973 2244 979 2256
rect 957 2203 963 2236
rect 941 2197 963 2203
rect 941 2144 947 2197
rect 957 2157 972 2163
rect 877 2104 883 2116
rect 957 1964 963 2157
rect 989 2004 995 2236
rect 1021 2104 1027 2276
rect 1037 2144 1043 2396
rect 1197 2383 1203 2596
rect 1229 2584 1235 2676
rect 1325 2564 1331 2676
rect 1341 2664 1347 2676
rect 1229 2504 1235 2536
rect 1325 2524 1331 2556
rect 1341 2543 1347 2656
rect 1373 2584 1379 2616
rect 1389 2544 1395 2676
rect 1405 2624 1411 2716
rect 1421 2584 1427 2636
rect 1341 2537 1356 2543
rect 1242 2414 1254 2416
rect 1227 2406 1229 2414
rect 1237 2406 1239 2414
rect 1247 2406 1249 2414
rect 1257 2406 1259 2414
rect 1267 2406 1269 2414
rect 1242 2404 1254 2406
rect 1197 2377 1219 2383
rect 1213 2264 1219 2377
rect 1309 2320 1315 2358
rect 1341 2304 1347 2476
rect 1357 2464 1363 2536
rect 1389 2284 1395 2536
rect 1412 2517 1427 2523
rect 1245 2244 1251 2276
rect 1133 2184 1139 2236
rect 733 1920 739 1958
rect 909 1904 915 1916
rect 653 1884 659 1896
rect 829 1784 835 1856
rect 733 1764 739 1776
rect 909 1764 915 1896
rect 573 1204 579 1476
rect 589 1304 595 1476
rect 733 1464 739 1756
rect 765 1744 771 1756
rect 861 1724 867 1756
rect 829 1644 835 1700
rect 909 1624 915 1736
rect 925 1724 931 1856
rect 989 1763 995 1956
rect 989 1757 1004 1763
rect 957 1684 963 1696
rect 973 1520 979 1558
rect 669 1364 675 1456
rect 717 1424 723 1436
rect 669 1204 675 1356
rect 605 1064 611 1196
rect 701 1104 707 1316
rect 765 1244 771 1300
rect 733 1124 739 1176
rect 781 1084 787 1356
rect 797 1324 803 1496
rect 893 1384 899 1416
rect 973 1364 979 1436
rect 989 1424 995 1757
rect 1005 1724 1011 1736
rect 1021 1524 1027 2096
rect 1053 2084 1059 2116
rect 1197 2044 1203 2096
rect 1242 2014 1254 2016
rect 1227 2006 1229 2014
rect 1237 2006 1239 2014
rect 1247 2006 1249 2014
rect 1257 2006 1259 2014
rect 1267 2006 1269 2014
rect 1242 2004 1254 2006
rect 1229 1904 1235 1956
rect 1293 1924 1299 2116
rect 1325 2043 1331 2156
rect 1405 2124 1411 2476
rect 1325 2037 1347 2043
rect 1037 1564 1043 1836
rect 1197 1784 1203 1856
rect 1341 1784 1347 2037
rect 1421 1964 1427 2517
rect 1453 2324 1459 2716
rect 1485 2684 1491 2696
rect 1517 2684 1523 2896
rect 1629 2844 1635 2896
rect 1613 2704 1619 2736
rect 1629 2684 1635 2836
rect 1661 2724 1667 2917
rect 1677 2824 1683 2896
rect 1661 2704 1667 2716
rect 1517 2644 1523 2656
rect 1581 2564 1587 2656
rect 1661 2604 1667 2636
rect 1677 2624 1683 2676
rect 1613 2544 1619 2556
rect 1693 2524 1699 2876
rect 1709 2804 1715 3076
rect 1757 3064 1763 3096
rect 1773 2984 1779 3116
rect 1805 3104 1811 3316
rect 1821 3224 1827 3356
rect 1869 3324 1875 3336
rect 1885 3284 1891 3296
rect 1821 3124 1827 3176
rect 1805 3064 1811 3096
rect 1869 3064 1875 3236
rect 1917 3184 1923 3356
rect 1949 3184 1955 3376
rect 2141 3364 2147 3437
rect 1789 3024 1795 3056
rect 1725 2844 1731 2916
rect 1741 2904 1747 2916
rect 1757 2763 1763 2936
rect 1741 2757 1763 2763
rect 1741 2744 1747 2757
rect 1725 2724 1731 2736
rect 1789 2724 1795 2816
rect 1805 2724 1811 2936
rect 1837 2903 1843 3036
rect 1853 2904 1859 3016
rect 1869 2944 1875 3056
rect 1901 2924 1907 3096
rect 1917 3064 1923 3116
rect 1965 3103 1971 3316
rect 2125 3304 2131 3336
rect 1997 3164 2003 3296
rect 1956 3097 1971 3103
rect 1981 3077 1996 3083
rect 1965 2963 1971 3076
rect 1981 2964 1987 3077
rect 2013 3063 2019 3116
rect 2029 3104 2035 3236
rect 2109 3223 2115 3236
rect 2093 3217 2115 3223
rect 2061 3124 2067 3216
rect 2093 3144 2099 3217
rect 2093 3104 2099 3136
rect 2109 3084 2115 3176
rect 2125 3084 2131 3216
rect 2141 3184 2147 3356
rect 2205 3324 2211 3496
rect 2285 3364 2291 3456
rect 2317 3444 2323 3476
rect 2477 3364 2483 3536
rect 2493 3504 2499 3556
rect 2541 3544 2547 3556
rect 2557 3524 2563 3656
rect 2685 3524 2691 3576
rect 2701 3524 2707 3756
rect 2733 3744 2739 3756
rect 2989 3724 2995 3736
rect 2813 3544 2819 3716
rect 2973 3704 2979 3716
rect 2829 3644 2835 3696
rect 2925 3644 2931 3676
rect 2989 3624 2995 3716
rect 3021 3544 3027 3596
rect 3037 3584 3043 3696
rect 3053 3644 3059 3656
rect 3037 3524 3043 3556
rect 3053 3524 3059 3636
rect 3069 3624 3075 3736
rect 3277 3724 3283 3776
rect 3421 3764 3427 3776
rect 3085 3664 3091 3696
rect 3101 3564 3107 3676
rect 3117 3584 3123 3656
rect 2557 3504 2563 3516
rect 2573 3484 2579 3516
rect 2653 3384 2659 3436
rect 2189 3124 2195 3136
rect 2205 3123 2211 3236
rect 2205 3117 2220 3123
rect 2004 3057 2019 3063
rect 2029 3024 2035 3036
rect 1949 2957 1971 2963
rect 1908 2917 1916 2923
rect 1828 2897 1843 2903
rect 1821 2884 1827 2896
rect 1469 2384 1475 2456
rect 1501 2344 1507 2496
rect 1517 2462 1523 2500
rect 1581 2484 1587 2516
rect 1453 2264 1459 2276
rect 1517 2264 1523 2416
rect 1469 2204 1475 2236
rect 1517 2164 1523 2256
rect 1549 2124 1555 2156
rect 1565 2144 1571 2316
rect 1581 2304 1587 2316
rect 1613 2304 1619 2336
rect 1629 2304 1635 2316
rect 1597 2284 1603 2296
rect 1597 2224 1603 2276
rect 1517 2104 1523 2116
rect 1597 2104 1603 2136
rect 1613 2124 1619 2136
rect 1629 2124 1635 2216
rect 1645 2144 1651 2316
rect 1693 2304 1699 2516
rect 1709 2344 1715 2716
rect 1741 2644 1747 2696
rect 1757 2384 1763 2676
rect 1773 2584 1779 2696
rect 1789 2664 1795 2716
rect 1805 2663 1811 2716
rect 1821 2684 1827 2696
rect 1837 2663 1843 2716
rect 1805 2657 1843 2663
rect 1821 2584 1827 2657
rect 1821 2384 1827 2476
rect 1805 2324 1811 2336
rect 1709 2284 1715 2316
rect 1693 2244 1699 2276
rect 1725 2244 1731 2280
rect 1677 2144 1683 2196
rect 1693 2144 1699 2156
rect 1741 2144 1747 2276
rect 1757 2184 1763 2236
rect 1773 2164 1779 2276
rect 1789 2264 1795 2316
rect 1469 1924 1475 1976
rect 1485 1904 1491 1916
rect 1341 1764 1347 1776
rect 1069 1724 1075 1736
rect 1101 1564 1107 1716
rect 1261 1662 1267 1716
rect 1188 1637 1203 1643
rect 1197 1584 1203 1637
rect 1242 1614 1254 1616
rect 1227 1606 1229 1614
rect 1237 1606 1239 1614
rect 1247 1606 1249 1614
rect 1257 1606 1259 1614
rect 1267 1606 1269 1614
rect 1242 1604 1254 1606
rect 797 1084 803 1096
rect 637 1064 643 1076
rect 605 1023 611 1056
rect 605 1017 627 1023
rect 397 924 403 936
rect 413 904 419 916
rect 445 904 451 976
rect 381 884 387 896
rect 461 704 467 956
rect 253 644 259 656
rect 13 544 19 556
rect 29 384 35 536
rect 93 204 99 556
rect 125 544 131 556
rect 221 524 227 576
rect 253 504 259 536
rect 285 523 291 696
rect 317 684 323 696
rect 477 683 483 896
rect 493 704 499 976
rect 621 964 627 1017
rect 813 984 819 1036
rect 509 684 515 936
rect 621 824 627 956
rect 701 862 707 916
rect 797 884 803 956
rect 829 924 835 1036
rect 845 924 851 1076
rect 820 897 835 903
rect 653 784 659 816
rect 525 684 531 736
rect 797 704 803 876
rect 829 784 835 897
rect 845 744 851 916
rect 861 744 867 1216
rect 877 1124 883 1176
rect 909 1124 915 1336
rect 925 1324 931 1356
rect 941 1224 947 1336
rect 1005 1324 1011 1496
rect 1053 1424 1059 1496
rect 1085 1484 1091 1556
rect 1149 1504 1155 1536
rect 1165 1444 1171 1476
rect 1181 1464 1187 1516
rect 1197 1504 1203 1576
rect 1197 1464 1203 1496
rect 1341 1484 1347 1756
rect 1021 1184 1027 1396
rect 1117 1364 1123 1436
rect 1341 1364 1347 1476
rect 1117 1324 1123 1336
rect 1053 1262 1059 1300
rect 973 1044 979 1076
rect 1085 1004 1091 1096
rect 1149 1064 1155 1356
rect 1437 1344 1443 1436
rect 1229 1324 1235 1336
rect 1453 1324 1459 1556
rect 1437 1317 1452 1323
rect 1293 1237 1308 1243
rect 1165 1184 1171 1236
rect 1197 1184 1203 1216
rect 1242 1214 1254 1216
rect 1227 1206 1229 1214
rect 1237 1206 1239 1214
rect 1247 1206 1249 1214
rect 1257 1206 1259 1214
rect 1267 1206 1269 1214
rect 1242 1204 1254 1206
rect 1165 1104 1171 1176
rect 1293 1064 1299 1237
rect 1341 1064 1347 1116
rect 1373 1084 1379 1236
rect 1437 1104 1443 1317
rect 1501 1304 1507 1996
rect 1533 1704 1539 1716
rect 1549 1644 1555 1696
rect 1565 1623 1571 1876
rect 1677 1764 1683 1856
rect 1741 1824 1747 2116
rect 1757 2004 1763 2036
rect 1773 1983 1779 2156
rect 1789 2144 1795 2216
rect 1837 2164 1843 2657
rect 1853 2564 1859 2796
rect 1885 2704 1891 2776
rect 1933 2744 1939 2836
rect 1901 2724 1907 2736
rect 1949 2723 1955 2957
rect 1981 2944 1987 2956
rect 1965 2924 1971 2936
rect 1997 2924 2003 3016
rect 2013 2984 2019 2996
rect 2020 2937 2035 2943
rect 2029 2924 2035 2937
rect 1972 2917 1987 2923
rect 1981 2784 1987 2917
rect 1949 2717 1964 2723
rect 1949 2684 1955 2696
rect 1892 2677 1907 2683
rect 1885 2584 1891 2636
rect 1901 2584 1907 2677
rect 1860 2537 1875 2543
rect 1853 2304 1859 2396
rect 1869 2284 1875 2537
rect 1885 2344 1891 2496
rect 1917 2343 1923 2676
rect 1933 2584 1939 2656
rect 2013 2603 2019 2896
rect 2029 2724 2035 2916
rect 2061 2764 2067 2916
rect 2093 2704 2099 2716
rect 2125 2703 2131 2956
rect 2157 2943 2163 3116
rect 2221 3104 2227 3116
rect 2269 3084 2275 3176
rect 2173 2944 2179 3036
rect 2189 2964 2195 3036
rect 2205 2984 2211 3056
rect 2285 2963 2291 3036
rect 2301 2984 2307 3156
rect 2333 3124 2339 3196
rect 2365 3164 2371 3356
rect 2461 3262 2467 3300
rect 2445 3184 2451 3216
rect 2381 3084 2387 3176
rect 2381 2984 2387 3056
rect 2269 2957 2291 2963
rect 2148 2937 2163 2943
rect 2125 2697 2140 2703
rect 1997 2597 2019 2603
rect 1933 2504 1939 2576
rect 1997 2564 2003 2597
rect 1981 2557 1996 2563
rect 1949 2384 1955 2556
rect 1981 2524 1987 2557
rect 2013 2544 2019 2576
rect 2045 2344 2051 2656
rect 2093 2564 2099 2696
rect 2109 2664 2115 2696
rect 2157 2684 2163 2937
rect 2205 2924 2211 2936
rect 2269 2924 2275 2957
rect 2285 2924 2291 2936
rect 2349 2924 2355 2956
rect 2429 2944 2435 2976
rect 2365 2924 2371 2936
rect 2253 2804 2259 2916
rect 2333 2904 2339 2916
rect 2205 2664 2211 2716
rect 2317 2704 2323 2876
rect 2349 2724 2355 2736
rect 2365 2723 2371 2916
rect 2397 2903 2403 2936
rect 2445 2924 2451 3096
rect 2477 3064 2483 3116
rect 2541 3104 2547 3336
rect 2397 2897 2419 2903
rect 2365 2717 2387 2723
rect 2317 2684 2323 2696
rect 2381 2684 2387 2717
rect 2413 2684 2419 2897
rect 2445 2884 2451 2916
rect 2429 2704 2435 2736
rect 2141 2584 2147 2656
rect 2237 2544 2243 2556
rect 2349 2544 2355 2636
rect 1901 2337 1923 2343
rect 1901 2324 1907 2337
rect 1949 2304 1955 2336
rect 1869 2244 1875 2276
rect 1965 2224 1971 2276
rect 1853 2124 1859 2216
rect 1885 2144 1891 2156
rect 1805 1984 1811 2116
rect 1949 2104 1955 2156
rect 1997 2144 2003 2196
rect 1997 2104 2003 2136
rect 2013 2063 2019 2156
rect 2061 2123 2067 2236
rect 2093 2184 2099 2316
rect 2125 2284 2131 2416
rect 2237 2383 2243 2536
rect 2221 2377 2243 2383
rect 2125 2144 2131 2276
rect 2221 2264 2227 2377
rect 2333 2304 2339 2516
rect 2413 2504 2419 2676
rect 2445 2664 2451 2676
rect 2429 2584 2435 2656
rect 2365 2444 2371 2496
rect 2413 2424 2419 2496
rect 2349 2324 2355 2376
rect 2253 2264 2259 2276
rect 2445 2264 2451 2656
rect 2461 2624 2467 2976
rect 2493 2964 2499 3096
rect 2557 2984 2563 3336
rect 2669 3164 2675 3516
rect 3037 3504 3043 3516
rect 2669 3064 2675 3156
rect 2701 3104 2707 3496
rect 2781 3464 2787 3476
rect 2813 3444 2819 3456
rect 3069 3444 3075 3496
rect 2746 3414 2758 3416
rect 2731 3406 2733 3414
rect 2741 3406 2743 3414
rect 2751 3406 2753 3414
rect 2761 3406 2763 3414
rect 2771 3406 2773 3414
rect 2746 3404 2758 3406
rect 2909 3384 2915 3436
rect 2909 3364 2915 3376
rect 2781 3244 2787 3296
rect 2797 3124 2803 3176
rect 2813 3104 2819 3316
rect 2877 3184 2883 3336
rect 3069 3264 3075 3436
rect 3069 3204 3075 3236
rect 2589 2964 2595 3036
rect 2669 2964 2675 3056
rect 2701 2984 2707 3076
rect 2746 3014 2758 3016
rect 2731 3006 2733 3014
rect 2741 3006 2743 3014
rect 2751 3006 2753 3014
rect 2761 3006 2763 3014
rect 2771 3006 2773 3014
rect 2746 3004 2758 3006
rect 2477 2664 2483 2896
rect 2509 2704 2515 2836
rect 2541 2824 2547 2936
rect 2573 2784 2579 2956
rect 2813 2804 2819 3096
rect 3085 3064 3091 3376
rect 3101 3324 3107 3456
rect 3117 3324 3123 3536
rect 3149 3524 3155 3716
rect 3197 3584 3203 3716
rect 3213 3544 3219 3656
rect 3261 3584 3267 3696
rect 3277 3664 3283 3696
rect 3293 3684 3299 3696
rect 3245 3544 3251 3576
rect 3213 3504 3219 3516
rect 3229 3484 3235 3536
rect 3181 3464 3187 3476
rect 3261 3444 3267 3496
rect 3277 3404 3283 3516
rect 3309 3504 3315 3756
rect 3357 3744 3363 3756
rect 3373 3704 3379 3716
rect 3325 3684 3331 3696
rect 3469 3584 3475 3736
rect 3373 3524 3379 3536
rect 3293 3444 3299 3456
rect 3325 3443 3331 3476
rect 3341 3464 3347 3496
rect 3373 3484 3379 3496
rect 3389 3484 3395 3496
rect 3405 3464 3411 3516
rect 3325 3437 3347 3443
rect 3261 3364 3267 3376
rect 3149 3224 3155 3316
rect 3165 3262 3171 3300
rect 3117 3104 3123 3156
rect 3181 3120 3187 3216
rect 3229 3124 3235 3336
rect 3325 3144 3331 3196
rect 2925 2984 2931 3036
rect 2957 2944 2963 2956
rect 3053 2924 3059 3016
rect 3021 2862 3027 2900
rect 2557 2704 2563 2716
rect 2893 2704 2899 2756
rect 2957 2720 2963 2796
rect 2493 2664 2499 2696
rect 2541 2684 2547 2696
rect 2381 2257 2396 2263
rect 2205 2144 2211 2216
rect 2221 2164 2227 2256
rect 2381 2204 2387 2257
rect 2061 2117 2076 2123
rect 1997 2057 2019 2063
rect 1764 1977 1779 1983
rect 1645 1744 1651 1756
rect 1677 1724 1683 1756
rect 1757 1724 1763 1896
rect 1789 1744 1795 1836
rect 1549 1617 1571 1623
rect 1517 1524 1523 1576
rect 1517 1344 1523 1496
rect 1549 1384 1555 1617
rect 1645 1464 1651 1716
rect 1757 1623 1763 1716
rect 1741 1617 1763 1623
rect 1741 1503 1747 1617
rect 1732 1497 1747 1503
rect 1613 1344 1619 1436
rect 1517 1283 1523 1316
rect 1501 1277 1523 1283
rect 1501 1104 1507 1277
rect 1597 1184 1603 1276
rect 1645 1224 1651 1456
rect 1725 1384 1731 1456
rect 1661 1344 1667 1356
rect 1725 1324 1731 1336
rect 1693 1304 1699 1316
rect 1709 1297 1724 1303
rect 877 784 883 936
rect 957 924 963 936
rect 1037 924 1043 996
rect 1149 964 1155 1056
rect 1053 862 1059 900
rect 1242 814 1254 816
rect 1227 806 1229 814
rect 1237 806 1239 814
rect 1247 806 1249 814
rect 1257 806 1259 814
rect 1267 806 1269 814
rect 1242 804 1254 806
rect 749 697 764 703
rect 749 684 755 697
rect 461 677 483 683
rect 301 624 307 656
rect 317 563 323 676
rect 397 664 403 676
rect 429 664 435 676
rect 349 584 355 616
rect 381 584 387 636
rect 397 564 403 656
rect 445 644 451 676
rect 317 557 339 563
rect 301 524 307 556
rect 333 544 339 557
rect 276 517 291 523
rect 205 384 211 436
rect 269 404 275 436
rect 221 284 227 396
rect 397 383 403 556
rect 461 524 467 677
rect 493 604 499 636
rect 557 603 563 676
rect 541 597 563 603
rect 541 544 547 597
rect 749 564 755 676
rect 388 377 403 383
rect 317 324 323 376
rect 461 304 467 516
rect 477 444 483 500
rect 573 444 579 556
rect 765 544 771 676
rect 29 184 35 196
rect 189 164 195 256
rect 317 124 323 296
rect 541 264 547 436
rect 669 324 675 376
rect 541 223 547 256
rect 669 224 675 296
rect 765 284 771 536
rect 525 217 547 223
rect 525 164 531 217
rect 605 124 611 216
rect 701 124 707 136
rect 317 44 323 96
rect 429 44 435 100
rect 717 -17 723 236
rect 781 144 787 696
rect 797 304 803 696
rect 813 584 819 736
rect 1213 724 1219 776
rect 877 584 883 656
rect 925 244 931 636
rect 1037 544 1043 556
rect 941 304 947 496
rect 973 320 979 358
rect 877 164 883 236
rect 941 224 947 296
rect 829 124 835 136
rect 909 124 915 216
rect 1005 164 1011 216
rect 1037 204 1043 276
rect 1069 264 1075 556
rect 1149 462 1155 516
rect 1197 304 1203 696
rect 1309 544 1315 696
rect 1325 604 1331 1056
rect 1357 944 1363 1036
rect 1389 1004 1395 1096
rect 1405 984 1411 1036
rect 1437 1024 1443 1056
rect 1437 964 1443 1016
rect 1453 944 1459 1076
rect 1501 1024 1507 1096
rect 1453 804 1459 936
rect 1517 903 1523 1076
rect 1533 984 1539 1116
rect 1597 1064 1603 1156
rect 1645 1104 1651 1136
rect 1709 1124 1715 1297
rect 1741 1084 1747 1497
rect 1757 1384 1763 1496
rect 1789 1304 1795 1736
rect 1821 1423 1827 1876
rect 1997 1864 2003 2057
rect 2141 2044 2147 2116
rect 2157 2104 2163 2136
rect 2013 1983 2019 2036
rect 2013 1977 2035 1983
rect 2029 1884 2035 1977
rect 2125 1924 2131 1976
rect 2189 1944 2195 2136
rect 2237 1984 2243 2156
rect 2269 2144 2275 2196
rect 2333 2124 2339 2156
rect 2109 1724 2115 1896
rect 2189 1864 2195 1876
rect 2221 1864 2227 1936
rect 2237 1844 2243 1896
rect 2269 1824 2275 2116
rect 2285 2084 2291 2116
rect 2285 1944 2291 2056
rect 2317 1924 2323 2096
rect 2333 1924 2339 2076
rect 2285 1864 2291 1916
rect 2333 1883 2339 1916
rect 2381 1884 2387 2196
rect 2445 2144 2451 2256
rect 2404 2117 2419 2123
rect 2413 2104 2419 2117
rect 2397 2084 2403 2096
rect 2333 1877 2355 1883
rect 2189 1724 2195 1756
rect 1965 1704 1971 1716
rect 1837 1524 1843 1636
rect 1901 1544 1907 1696
rect 1805 1417 1827 1423
rect 1805 1164 1811 1417
rect 1837 1403 1843 1516
rect 1933 1504 1939 1516
rect 1997 1504 2003 1696
rect 1821 1397 1843 1403
rect 1821 1364 1827 1397
rect 1853 1323 1859 1496
rect 2013 1464 2019 1516
rect 2029 1464 2035 1636
rect 2189 1504 2195 1636
rect 2205 1524 2211 1616
rect 2077 1484 2083 1496
rect 2109 1464 2115 1496
rect 1844 1317 1859 1323
rect 1789 1124 1795 1136
rect 1837 1124 1843 1176
rect 1837 1084 1843 1096
rect 1613 1044 1619 1056
rect 1757 1044 1763 1076
rect 1837 984 1843 1076
rect 1853 964 1859 1276
rect 1997 1224 2003 1356
rect 2173 1324 2179 1356
rect 1965 1064 1971 1216
rect 1965 1023 1971 1056
rect 1965 1017 1987 1023
rect 1508 897 1523 903
rect 1549 884 1555 936
rect 1613 904 1619 918
rect 1341 784 1347 796
rect 1533 704 1539 756
rect 1325 564 1331 596
rect 1341 584 1347 676
rect 1389 564 1395 576
rect 1444 557 1475 563
rect 1242 414 1254 416
rect 1227 406 1229 414
rect 1237 406 1239 414
rect 1247 406 1249 414
rect 1257 406 1259 414
rect 1267 406 1269 414
rect 1242 404 1254 406
rect 1069 224 1075 256
rect 1197 164 1203 236
rect 1213 184 1219 196
rect 749 -17 755 116
rect 1309 104 1315 536
rect 1373 523 1379 556
rect 1364 517 1379 523
rect 1469 523 1475 557
rect 1485 544 1491 616
rect 1597 584 1603 676
rect 1645 664 1651 936
rect 1677 724 1683 736
rect 1709 704 1715 916
rect 1853 864 1859 956
rect 1885 924 1891 996
rect 1940 957 1964 963
rect 1757 724 1763 776
rect 1773 704 1779 716
rect 1709 564 1715 576
rect 1549 524 1555 556
rect 1469 517 1484 523
rect 1453 504 1459 516
rect 1597 504 1603 556
rect 1661 524 1667 556
rect 1341 384 1347 496
rect 1357 244 1363 336
rect 1357 144 1363 236
rect 1421 144 1427 436
rect 1661 424 1667 516
rect 1773 504 1779 696
rect 1533 304 1539 356
rect 1629 324 1635 396
rect 1629 304 1635 316
rect 1501 224 1507 256
rect 1533 244 1539 276
rect 1549 164 1555 216
rect 1661 124 1667 396
rect 1693 384 1699 416
rect 1789 404 1795 836
rect 1933 804 1939 836
rect 1853 684 1859 796
rect 1981 664 1987 1017
rect 2077 964 2083 1056
rect 2045 904 2051 936
rect 2077 924 2083 956
rect 2093 944 2099 976
rect 2045 884 2051 896
rect 2045 784 2051 876
rect 2093 784 2099 936
rect 2109 704 2115 1316
rect 2205 1304 2211 1516
rect 2221 1504 2227 1716
rect 2301 1684 2307 1856
rect 2333 1804 2339 1836
rect 2317 1644 2323 1696
rect 2349 1664 2355 1877
rect 2381 1864 2387 1876
rect 2365 1644 2371 1756
rect 2381 1644 2387 1716
rect 2285 1520 2291 1558
rect 2381 1464 2387 1636
rect 2397 1584 2403 1836
rect 2429 1624 2435 2076
rect 2461 1903 2467 2116
rect 2477 2064 2483 2436
rect 2493 2344 2499 2656
rect 2557 2644 2563 2696
rect 2589 2664 2595 2696
rect 2605 2664 2611 2676
rect 2525 2604 2531 2636
rect 2746 2614 2758 2616
rect 2731 2606 2733 2614
rect 2741 2606 2743 2614
rect 2751 2606 2753 2614
rect 2761 2606 2763 2614
rect 2771 2606 2773 2614
rect 2746 2604 2758 2606
rect 2861 2604 2867 2656
rect 2861 2564 2867 2596
rect 2893 2584 2899 2656
rect 3053 2624 3059 2916
rect 3069 2724 3075 2796
rect 3085 2664 3091 3056
rect 3117 2944 3123 3076
rect 3181 3024 3187 3112
rect 3261 3104 3267 3136
rect 3229 3024 3235 3096
rect 3229 2944 3235 3016
rect 3277 2984 3283 3076
rect 3309 3064 3315 3076
rect 3309 2964 3315 2976
rect 3229 2924 3235 2936
rect 3101 2604 3107 2916
rect 3293 2884 3299 2896
rect 3165 2704 3171 2756
rect 3165 2604 3171 2676
rect 3053 2564 3059 2596
rect 2557 2462 2563 2516
rect 2637 2424 2643 2556
rect 2669 2424 2675 2536
rect 2573 2264 2579 2416
rect 2669 2320 2675 2358
rect 2765 2324 2771 2496
rect 2973 2462 2979 2516
rect 3053 2384 3059 2556
rect 3085 2404 3091 2536
rect 3181 2504 3187 2616
rect 3229 2584 3235 2596
rect 2765 2304 2771 2316
rect 3021 2264 3027 2376
rect 3053 2304 3059 2356
rect 3053 2264 3059 2276
rect 2573 2204 2579 2256
rect 2746 2214 2758 2216
rect 2731 2206 2733 2214
rect 2741 2206 2743 2214
rect 2751 2206 2753 2214
rect 2761 2206 2763 2214
rect 2771 2206 2773 2214
rect 2746 2204 2758 2206
rect 2477 1924 2483 2036
rect 2461 1897 2483 1903
rect 2445 1784 2451 1856
rect 2477 1743 2483 1897
rect 2493 1864 2499 1896
rect 2509 1744 2515 2176
rect 2557 2064 2563 2176
rect 2637 2164 2643 2196
rect 2669 2104 2675 2136
rect 2525 1904 2531 1916
rect 2541 1784 2547 1896
rect 2557 1744 2563 2056
rect 2733 2044 2739 2100
rect 2589 1784 2595 2016
rect 2845 1864 2851 2216
rect 2861 2164 2867 2236
rect 3021 2224 3027 2256
rect 2893 2184 2899 2196
rect 3085 2164 3091 2216
rect 2861 2144 2867 2156
rect 3181 2124 3187 2496
rect 3213 2384 3219 2556
rect 3277 2544 3283 2616
rect 3229 2504 3235 2536
rect 3293 2504 3299 2516
rect 3245 2284 3251 2316
rect 3293 2303 3299 2496
rect 3309 2364 3315 2876
rect 3325 2704 3331 3136
rect 3341 3103 3347 3437
rect 3421 3404 3427 3496
rect 3453 3424 3459 3456
rect 3373 3144 3379 3396
rect 3485 3384 3491 3816
rect 3421 3184 3427 3376
rect 3437 3324 3443 3336
rect 3341 3097 3356 3103
rect 3373 3084 3379 3136
rect 3437 3004 3443 3276
rect 3469 3184 3475 3236
rect 3469 3104 3475 3176
rect 3485 3144 3491 3336
rect 3453 2984 3459 3096
rect 3469 3044 3475 3076
rect 3469 2924 3475 2936
rect 3357 2904 3363 2916
rect 3437 2864 3443 2916
rect 3373 2584 3379 2596
rect 3389 2544 3395 2716
rect 3405 2624 3411 2636
rect 3421 2604 3427 2676
rect 3405 2564 3411 2576
rect 3325 2304 3331 2316
rect 3293 2297 3315 2303
rect 3229 2224 3235 2276
rect 3005 2062 3011 2116
rect 3181 2108 3187 2116
rect 2941 1920 2947 1958
rect 2573 1744 2579 1756
rect 2605 1744 2611 1796
rect 2477 1737 2499 1743
rect 2493 1724 2499 1737
rect 2461 1624 2467 1696
rect 2493 1424 2499 1716
rect 2509 1704 2515 1736
rect 2621 1724 2627 1856
rect 2525 1704 2531 1716
rect 2525 1663 2531 1696
rect 2509 1657 2531 1663
rect 2285 1344 2291 1396
rect 2333 1324 2339 1416
rect 2509 1384 2515 1657
rect 2557 1524 2563 1536
rect 2541 1364 2547 1436
rect 2381 1324 2387 1336
rect 2541 1324 2547 1356
rect 2125 1244 2131 1296
rect 2141 1164 2147 1196
rect 2125 1124 2131 1136
rect 2141 1064 2147 1156
rect 2221 1124 2227 1176
rect 2269 1124 2275 1316
rect 2221 1004 2227 1116
rect 2253 1064 2259 1076
rect 2253 984 2259 1056
rect 2189 964 2195 976
rect 2317 964 2323 1316
rect 2493 1304 2499 1316
rect 2365 1104 2371 1276
rect 2461 1144 2467 1236
rect 2340 1077 2355 1083
rect 2349 1024 2355 1077
rect 2397 1064 2403 1116
rect 2493 1084 2499 1296
rect 2509 1184 2515 1236
rect 2525 1104 2531 1136
rect 2557 1104 2563 1516
rect 2573 1364 2579 1696
rect 2589 1584 2595 1656
rect 2605 1484 2611 1496
rect 2605 1344 2611 1476
rect 2637 1464 2643 1856
rect 2669 1724 2675 1756
rect 2685 1704 2691 1836
rect 2701 1764 2707 1816
rect 2746 1814 2758 1816
rect 2731 1806 2733 1814
rect 2741 1806 2743 1814
rect 2751 1806 2753 1814
rect 2761 1806 2763 1814
rect 2771 1806 2773 1814
rect 2746 1804 2758 1806
rect 2813 1757 2867 1763
rect 2813 1724 2819 1757
rect 2861 1744 2867 1757
rect 2893 1744 2899 1756
rect 2685 1524 2691 1696
rect 2701 1584 2707 1716
rect 2925 1704 2931 1716
rect 2861 1584 2867 1676
rect 2669 1484 2675 1496
rect 2797 1484 2803 1536
rect 2909 1504 2915 1576
rect 2957 1504 2963 1956
rect 2973 1824 2979 1896
rect 3197 1864 3203 2216
rect 3261 2204 3267 2276
rect 3293 2264 3299 2276
rect 3309 2124 3315 2297
rect 3341 2284 3347 2536
rect 3453 2524 3459 2896
rect 3469 2724 3475 2916
rect 3501 2864 3507 3796
rect 3517 3664 3523 3696
rect 3645 3644 3651 3756
rect 3869 3724 3875 3736
rect 3725 3662 3731 3716
rect 3613 3584 3619 3616
rect 3693 3584 3699 3616
rect 3725 3524 3731 3576
rect 3517 3384 3523 3436
rect 3533 3344 3539 3496
rect 3565 3404 3571 3516
rect 3725 3504 3731 3516
rect 3549 3344 3555 3396
rect 3549 3324 3555 3336
rect 3517 3064 3523 3296
rect 3533 3224 3539 3316
rect 3533 3084 3539 3116
rect 3565 3084 3571 3256
rect 3581 3124 3587 3296
rect 3613 3284 3619 3496
rect 3629 3384 3635 3476
rect 3645 3464 3651 3476
rect 3661 3444 3667 3496
rect 3645 3403 3651 3416
rect 3677 3403 3683 3436
rect 3693 3423 3699 3496
rect 3709 3444 3715 3476
rect 3693 3417 3731 3423
rect 3645 3397 3683 3403
rect 3645 3344 3651 3356
rect 3725 3343 3731 3417
rect 3741 3364 3747 3496
rect 3757 3364 3763 3496
rect 3725 3337 3740 3343
rect 3757 3324 3763 3356
rect 3597 3184 3603 3276
rect 3661 3224 3667 3296
rect 3709 3244 3715 3316
rect 3757 3284 3763 3296
rect 3613 3124 3619 3136
rect 3517 2944 3523 3056
rect 3597 2984 3603 3096
rect 3645 3064 3651 3216
rect 3693 3184 3699 3216
rect 3757 3204 3763 3276
rect 3613 2964 3619 3036
rect 3629 2984 3635 3036
rect 3709 2984 3715 3136
rect 3757 3124 3763 3136
rect 3725 3044 3731 3076
rect 3773 3064 3779 3476
rect 3789 3464 3795 3536
rect 3805 3344 3811 3636
rect 3821 3484 3827 3576
rect 3869 3564 3875 3716
rect 3885 3684 3891 3696
rect 3901 3624 3907 3676
rect 3981 3644 3987 3696
rect 3997 3664 4003 3716
rect 4077 3684 4083 3736
rect 4109 3644 4115 3756
rect 3885 3584 3891 3596
rect 3837 3504 3843 3536
rect 3869 3484 3875 3556
rect 3917 3484 3923 3616
rect 3933 3504 3939 3596
rect 3949 3563 3955 3616
rect 3981 3583 3987 3596
rect 4061 3584 4067 3596
rect 3972 3577 3987 3583
rect 3949 3557 3987 3563
rect 3949 3463 3955 3496
rect 3965 3484 3971 3516
rect 3981 3504 3987 3557
rect 3997 3557 4083 3563
rect 3997 3544 4003 3557
rect 4077 3544 4083 3557
rect 4013 3504 4019 3536
rect 3949 3457 3971 3463
rect 3885 3384 3891 3456
rect 3965 3444 3971 3457
rect 3949 3384 3955 3436
rect 3997 3384 4003 3456
rect 4013 3444 4019 3496
rect 4029 3484 4035 3516
rect 4061 3504 4067 3536
rect 3917 3324 3923 3356
rect 3981 3344 3987 3356
rect 3789 3104 3795 3256
rect 3821 3084 3827 3316
rect 3933 3244 3939 3336
rect 3869 3144 3875 3236
rect 3981 3144 3987 3296
rect 3997 3184 4003 3276
rect 4029 3204 4035 3336
rect 4045 3264 4051 3496
rect 4077 3464 4083 3516
rect 4093 3464 4099 3556
rect 4125 3544 4131 3616
rect 4250 3614 4262 3616
rect 4235 3606 4237 3614
rect 4245 3606 4247 3614
rect 4255 3606 4257 3614
rect 4265 3606 4267 3614
rect 4275 3606 4277 3614
rect 4250 3604 4262 3606
rect 4461 3584 4467 3736
rect 4205 3524 4211 3536
rect 4413 3524 4419 3576
rect 4541 3544 4547 3756
rect 4573 3584 4579 3736
rect 4205 3464 4211 3496
rect 4093 3344 4099 3436
rect 4221 3364 4227 3496
rect 4237 3364 4243 3456
rect 4173 3344 4179 3356
rect 4077 3284 4083 3316
rect 4093 3263 4099 3296
rect 4084 3257 4099 3263
rect 4077 3184 4083 3216
rect 3837 3104 3843 3116
rect 3869 3104 3875 3136
rect 4077 3124 4083 3136
rect 4093 3124 4099 3196
rect 3924 3117 3980 3123
rect 4100 3117 4115 3123
rect 3789 2984 3795 3076
rect 3901 3004 3907 3056
rect 3965 2984 3971 3076
rect 3997 3064 4003 3096
rect 4077 3084 4083 3096
rect 4061 2984 4067 3076
rect 3469 2564 3475 2636
rect 3485 2584 3491 2616
rect 3357 2344 3363 2516
rect 3469 2497 3484 2503
rect 3357 2304 3363 2336
rect 3396 2317 3411 2323
rect 3373 2304 3379 2316
rect 3389 2304 3395 2316
rect 3341 1964 3347 2156
rect 3389 2124 3395 2196
rect 3357 2104 3363 2116
rect 3229 1904 3235 1956
rect 3037 1764 3043 1836
rect 3229 1784 3235 1876
rect 3325 1824 3331 1916
rect 3357 1864 3363 2096
rect 3373 1904 3379 1936
rect 3373 1864 3379 1896
rect 3037 1524 3043 1756
rect 3117 1644 3123 1756
rect 3149 1744 3155 1776
rect 3245 1724 3251 1816
rect 3325 1744 3331 1796
rect 3149 1504 3155 1556
rect 3213 1520 3219 1716
rect 3245 1644 3251 1696
rect 2813 1483 2819 1496
rect 2813 1480 2828 1483
rect 2813 1477 2835 1480
rect 2653 1384 2659 1476
rect 2509 1084 2515 1096
rect 2525 1084 2531 1096
rect 2125 944 2131 956
rect 2189 944 2195 956
rect 2221 924 2227 956
rect 2285 944 2291 956
rect 2349 944 2355 956
rect 2253 923 2259 936
rect 2365 924 2371 936
rect 2237 917 2259 923
rect 2221 904 2227 916
rect 2237 884 2243 917
rect 2381 884 2387 936
rect 2413 924 2419 1056
rect 2429 964 2435 1076
rect 2429 904 2435 956
rect 2445 944 2451 1056
rect 2541 1044 2547 1076
rect 2573 1064 2579 1316
rect 2605 1304 2611 1316
rect 2637 1304 2643 1316
rect 2669 1204 2675 1456
rect 2746 1414 2758 1416
rect 2731 1406 2733 1414
rect 2741 1406 2743 1414
rect 2751 1406 2753 1414
rect 2761 1406 2763 1414
rect 2771 1406 2773 1414
rect 2746 1404 2758 1406
rect 2589 1104 2595 1116
rect 2461 924 2467 996
rect 2477 943 2483 1036
rect 2509 984 2515 1016
rect 2589 984 2595 1096
rect 2621 1004 2627 1076
rect 2669 1064 2675 1196
rect 2749 1104 2755 1276
rect 2813 1262 2819 1316
rect 2893 1243 2899 1356
rect 3101 1324 3107 1416
rect 2893 1237 2915 1243
rect 2909 1064 2915 1237
rect 2941 1104 2947 1156
rect 3037 1124 3043 1296
rect 2477 937 2499 943
rect 2317 804 2323 836
rect 2285 684 2291 796
rect 2349 720 2355 758
rect 1901 524 1907 536
rect 1805 404 1811 496
rect 1933 424 1939 556
rect 2013 462 2019 516
rect 1853 264 1859 416
rect 1885 304 1891 356
rect 1949 320 1955 396
rect 2029 284 2035 536
rect 2125 503 2131 536
rect 2141 524 2147 596
rect 2189 504 2195 596
rect 2125 497 2147 503
rect 2109 304 2115 476
rect 2141 344 2147 497
rect 2125 284 2131 296
rect 1757 124 1763 236
rect 1853 224 1859 256
rect 2029 224 2035 276
rect 2125 243 2131 276
rect 2141 264 2147 296
rect 2237 284 2243 536
rect 2269 524 2275 556
rect 2301 524 2307 596
rect 2253 384 2259 496
rect 2269 324 2275 476
rect 2301 324 2307 516
rect 2397 504 2403 696
rect 2461 684 2467 696
rect 2477 664 2483 736
rect 2429 584 2435 656
rect 2493 604 2499 937
rect 2525 704 2531 716
rect 2605 704 2611 816
rect 2621 684 2627 976
rect 2637 944 2643 1036
rect 2746 1014 2758 1016
rect 2731 1006 2733 1014
rect 2741 1006 2743 1014
rect 2751 1006 2753 1014
rect 2761 1006 2763 1014
rect 2771 1006 2773 1014
rect 2746 1004 2758 1006
rect 2909 1004 2915 1056
rect 2861 964 2867 996
rect 2621 664 2627 676
rect 2637 664 2643 856
rect 2781 703 2787 916
rect 2861 804 2867 956
rect 3005 924 3011 1112
rect 3037 964 3043 1036
rect 3085 984 3091 1076
rect 2989 844 2995 896
rect 2781 697 2803 703
rect 2445 462 2451 516
rect 2525 424 2531 556
rect 2557 544 2563 556
rect 2701 524 2707 676
rect 2746 614 2758 616
rect 2731 606 2733 614
rect 2741 606 2743 614
rect 2751 606 2753 614
rect 2761 606 2763 614
rect 2771 606 2773 614
rect 2746 604 2758 606
rect 2797 504 2803 697
rect 2125 237 2147 243
rect 1981 164 1987 216
rect 2141 184 2147 237
rect 2173 144 2179 276
rect 2237 264 2243 276
rect 2269 144 2275 256
rect 1661 104 1667 116
rect 877 44 883 96
rect 1645 44 1651 100
rect 2061 62 2067 116
rect 2221 104 2227 116
rect 2301 104 2307 316
rect 2477 264 2483 416
rect 2509 304 2515 356
rect 2621 324 2627 496
rect 2797 284 2803 436
rect 2813 304 2819 316
rect 2509 244 2515 276
rect 2317 184 2323 236
rect 2333 144 2339 216
rect 2349 184 2355 236
rect 2381 144 2387 176
rect 2397 124 2403 156
rect 2445 144 2451 216
rect 2461 124 2467 176
rect 2621 144 2627 196
rect 2653 184 2659 256
rect 2669 204 2675 236
rect 2701 224 2707 276
rect 2717 244 2723 276
rect 2669 164 2675 176
rect 2429 104 2435 116
rect 2541 104 2547 116
rect 2573 104 2579 136
rect 2653 124 2659 156
rect 2701 144 2707 216
rect 2746 214 2758 216
rect 2731 206 2733 214
rect 2741 206 2743 214
rect 2751 206 2753 214
rect 2761 206 2763 214
rect 2771 206 2773 214
rect 2746 204 2758 206
rect 2628 117 2643 123
rect 2308 97 2316 103
rect 2637 103 2643 117
rect 2781 104 2787 136
rect 2813 124 2819 296
rect 2637 97 2652 103
rect 2253 84 2259 96
rect 2365 84 2371 96
rect 1242 14 1254 16
rect 1227 6 1229 14
rect 1237 6 1239 14
rect 1247 6 1249 14
rect 1257 6 1259 14
rect 1267 6 1269 14
rect 1242 4 1254 6
rect 1725 -17 1731 36
rect 1805 -17 1811 36
rect 2829 -17 2835 676
rect 2909 664 2915 796
rect 3053 764 3059 836
rect 3101 824 3107 1096
rect 3117 1064 3123 1456
rect 3149 1304 3155 1316
rect 3165 1304 3171 1336
rect 2941 704 2947 756
rect 2941 664 2947 676
rect 2909 604 2915 656
rect 3037 644 3043 716
rect 3085 704 3091 796
rect 3133 744 3139 1036
rect 3149 924 3155 1296
rect 3181 1124 3187 1396
rect 3197 1324 3203 1356
rect 3213 1344 3219 1436
rect 3261 1324 3267 1516
rect 3309 1464 3315 1636
rect 3341 1544 3347 1756
rect 3389 1724 3395 1856
rect 3405 1703 3411 2317
rect 3421 2264 3427 2296
rect 3453 2184 3459 2476
rect 3421 2164 3427 2176
rect 3421 2004 3427 2136
rect 3469 2104 3475 2497
rect 3485 2043 3491 2296
rect 3501 2264 3507 2856
rect 3549 2764 3555 2956
rect 3693 2924 3699 2956
rect 3565 2884 3571 2916
rect 3725 2884 3731 2936
rect 3757 2924 3763 2956
rect 3549 2704 3555 2712
rect 3613 2704 3619 2756
rect 3549 2524 3555 2696
rect 3613 2624 3619 2676
rect 3629 2544 3635 2556
rect 3549 2504 3555 2516
rect 3565 2462 3571 2500
rect 3629 2443 3635 2516
rect 3613 2437 3635 2443
rect 3565 2384 3571 2416
rect 3613 2384 3619 2437
rect 3485 2037 3507 2043
rect 3460 1917 3475 1923
rect 3421 1864 3427 1896
rect 3437 1704 3443 1856
rect 3389 1697 3411 1703
rect 3373 1504 3379 1556
rect 3389 1524 3395 1697
rect 3325 1424 3331 1496
rect 3373 1464 3379 1496
rect 3389 1424 3395 1516
rect 3405 1504 3411 1516
rect 3421 1504 3427 1696
rect 3437 1523 3443 1696
rect 3437 1517 3452 1523
rect 3437 1484 3443 1496
rect 3437 1444 3443 1476
rect 3453 1404 3459 1516
rect 3469 1504 3475 1917
rect 3485 1764 3491 1996
rect 3485 1744 3491 1756
rect 3501 1724 3507 2037
rect 3485 1704 3491 1716
rect 3501 1684 3507 1716
rect 3517 1584 3523 2356
rect 3549 2184 3555 2276
rect 3613 2144 3619 2356
rect 3645 2304 3651 2376
rect 3661 2364 3667 2556
rect 3757 2324 3763 2596
rect 3789 2384 3795 2976
rect 3837 2964 3843 2976
rect 3805 2864 3811 2916
rect 3821 2884 3827 2936
rect 3917 2884 3923 2936
rect 3933 2864 3939 2936
rect 3949 2924 3955 2936
rect 3981 2904 3987 2976
rect 4093 2964 4099 2996
rect 4109 2984 4115 3117
rect 4125 3084 4131 3236
rect 4141 3104 4147 3316
rect 4173 3064 4179 3336
rect 4189 3064 4195 3356
rect 4285 3264 4291 3376
rect 4349 3324 4355 3516
rect 4365 3384 4371 3476
rect 4397 3324 4403 3436
rect 4308 3317 4323 3323
rect 4250 3214 4262 3216
rect 4235 3206 4237 3214
rect 4245 3206 4247 3214
rect 4255 3206 4257 3214
rect 4265 3206 4267 3214
rect 4275 3206 4277 3214
rect 4250 3204 4262 3206
rect 4301 3104 4307 3116
rect 4029 2884 4035 2936
rect 3805 2584 3811 2636
rect 3661 2304 3667 2316
rect 3677 2304 3683 2316
rect 3661 2144 3667 2296
rect 3693 2204 3699 2296
rect 3709 2284 3715 2316
rect 3725 2264 3731 2276
rect 3709 2144 3715 2176
rect 3741 2144 3747 2236
rect 3581 2104 3587 2118
rect 3613 1983 3619 2136
rect 3645 2084 3651 2096
rect 3693 2044 3699 2136
rect 3757 2084 3763 2316
rect 3789 2164 3795 2236
rect 3613 1977 3635 1983
rect 3533 1824 3539 1912
rect 3597 1904 3603 1956
rect 3629 1864 3635 1977
rect 3533 1504 3539 1636
rect 3549 1584 3555 1776
rect 3565 1744 3571 1756
rect 3565 1604 3571 1736
rect 3597 1724 3603 1856
rect 3629 1844 3635 1856
rect 3709 1784 3715 2076
rect 3773 1924 3779 2116
rect 3789 1984 3795 2136
rect 3821 2104 3827 2136
rect 3837 2124 3843 2476
rect 3853 2244 3859 2436
rect 3869 2304 3875 2696
rect 3885 2564 3891 2856
rect 3901 2720 3907 2758
rect 4093 2704 4099 2956
rect 4141 2924 4147 3056
rect 4173 2744 4179 3056
rect 4189 2964 4195 3056
rect 4285 2864 4291 3056
rect 4301 2984 4307 3056
rect 4317 3044 4323 3317
rect 4381 3244 4387 3296
rect 4413 3284 4419 3296
rect 4317 2924 4323 3036
rect 4349 2924 4355 3156
rect 4397 3084 4403 3236
rect 4397 3044 4403 3056
rect 4413 2924 4419 3216
rect 4429 3184 4435 3456
rect 4477 3404 4483 3476
rect 4484 3397 4499 3403
rect 4445 3304 4451 3356
rect 4493 3344 4499 3397
rect 4509 3384 4515 3516
rect 4525 3484 4531 3516
rect 4541 3464 4547 3476
rect 4557 3424 4563 3496
rect 4605 3444 4611 3476
rect 4573 3364 4579 3416
rect 4637 3324 4643 3716
rect 4669 3644 4675 3696
rect 4781 3662 4787 3700
rect 4653 3364 4659 3496
rect 4733 3464 4739 3496
rect 4701 3404 4707 3456
rect 4733 3424 4739 3456
rect 4749 3364 4755 3536
rect 4765 3524 4771 3556
rect 4829 3524 4835 3536
rect 4781 3484 4787 3496
rect 4797 3464 4803 3496
rect 4845 3464 4851 3496
rect 4877 3484 4883 3596
rect 4925 3544 4931 3556
rect 4973 3504 4979 3516
rect 4877 3464 4883 3476
rect 4461 3304 4467 3316
rect 4525 3284 4531 3316
rect 4621 3244 4627 3296
rect 4250 2814 4262 2816
rect 4235 2806 4237 2814
rect 4245 2806 4247 2814
rect 4255 2806 4257 2814
rect 4265 2806 4267 2814
rect 4275 2806 4277 2814
rect 4250 2804 4262 2806
rect 4173 2664 4179 2736
rect 4221 2664 4227 2756
rect 3949 2264 3955 2556
rect 4045 2320 4051 2358
rect 3901 2144 3907 2216
rect 3965 2144 3971 2156
rect 3933 2097 3948 2103
rect 3805 2064 3811 2076
rect 3805 1924 3811 2056
rect 3885 2024 3891 2096
rect 3933 1984 3939 2097
rect 3997 2044 4003 2176
rect 4029 2144 4035 2216
rect 4093 2143 4099 2536
rect 4157 2444 4163 2500
rect 4189 2324 4195 2436
rect 4205 2384 4211 2636
rect 4221 2504 4227 2656
rect 4301 2544 4307 2556
rect 4317 2544 4323 2916
rect 4429 2904 4435 3176
rect 4445 3124 4451 3176
rect 4653 3104 4659 3316
rect 4445 3064 4451 3096
rect 4653 3004 4659 3096
rect 4749 3064 4755 3356
rect 4781 3184 4787 3216
rect 4845 3204 4851 3456
rect 4861 3304 4867 3436
rect 4461 2844 4467 2936
rect 4605 2924 4611 2996
rect 4685 2964 4691 3056
rect 4717 2924 4723 2936
rect 4781 2862 4787 2900
rect 4333 2584 4339 2676
rect 4250 2414 4262 2416
rect 4235 2406 4237 2414
rect 4245 2406 4247 2414
rect 4255 2406 4257 2414
rect 4265 2406 4267 2414
rect 4275 2406 4277 2414
rect 4250 2404 4262 2406
rect 4301 2343 4307 2356
rect 4269 2337 4307 2343
rect 4109 2164 4115 2236
rect 4125 2184 4131 2236
rect 4141 2224 4147 2236
rect 4109 2144 4115 2156
rect 4084 2137 4099 2143
rect 4013 2124 4019 2136
rect 4045 2103 4051 2136
rect 4125 2124 4131 2176
rect 4157 2164 4163 2316
rect 4173 2264 4179 2296
rect 4221 2203 4227 2336
rect 4269 2324 4275 2337
rect 4205 2197 4227 2203
rect 4157 2124 4163 2136
rect 4068 2117 4083 2123
rect 4045 2097 4067 2103
rect 3885 1904 3891 1916
rect 3901 1904 3907 1936
rect 3853 1864 3859 1896
rect 3613 1697 3628 1703
rect 3613 1504 3619 1697
rect 3677 1524 3683 1776
rect 3805 1764 3811 1836
rect 3709 1644 3715 1700
rect 3693 1504 3699 1536
rect 3485 1484 3491 1496
rect 3501 1484 3507 1496
rect 3565 1484 3571 1496
rect 3485 1364 3491 1476
rect 3581 1364 3587 1496
rect 3357 1324 3363 1336
rect 3181 1104 3187 1116
rect 3197 1004 3203 1316
rect 3293 1244 3299 1300
rect 3213 1064 3219 1096
rect 3245 1064 3251 1076
rect 3245 964 3251 1056
rect 3085 684 3091 696
rect 3117 664 3123 676
rect 2941 544 2947 636
rect 2973 564 2979 596
rect 3133 584 3139 736
rect 3149 724 3155 916
rect 3165 862 3171 916
rect 3149 704 3155 716
rect 3165 564 3171 816
rect 3213 704 3219 776
rect 3261 764 3267 836
rect 3213 684 3219 696
rect 3197 664 3203 676
rect 3053 462 3059 516
rect 3085 304 3091 356
rect 3149 320 3155 496
rect 2877 184 2883 276
rect 2893 184 2899 236
rect 3053 203 3059 256
rect 3053 197 3068 203
rect 3069 164 3075 196
rect 2989 62 2995 116
rect 3101 84 3107 136
rect 717 -23 739 -17
rect 749 -23 771 -17
rect 1725 -23 1747 -17
rect 1789 -23 1811 -17
rect 2813 -23 2835 -17
rect 3165 -23 3171 556
rect 3213 524 3219 636
rect 3213 104 3219 516
rect 3229 -17 3235 696
rect 3261 684 3267 756
rect 3309 704 3315 716
rect 3357 704 3363 1296
rect 3373 1084 3379 1236
rect 3373 1023 3379 1076
rect 3389 1064 3395 1356
rect 3581 1204 3587 1356
rect 3597 1304 3603 1496
rect 3709 1484 3715 1516
rect 3757 1504 3763 1556
rect 3773 1484 3779 1736
rect 3885 1724 3891 1816
rect 3917 1784 3923 1936
rect 3949 1924 3955 1936
rect 3981 1884 3987 1896
rect 3997 1884 4003 2036
rect 4013 1944 4019 2036
rect 4013 1904 4019 1916
rect 4013 1884 4019 1896
rect 3981 1684 3987 1876
rect 4013 1684 4019 1776
rect 4029 1724 4035 2076
rect 4061 2063 4067 2097
rect 4077 2084 4083 2117
rect 4061 2057 4083 2063
rect 4045 1924 4051 2056
rect 4077 1984 4083 2057
rect 4109 2004 4115 2076
rect 4109 1984 4115 1996
rect 4125 1944 4131 2096
rect 4173 2064 4179 2096
rect 4045 1844 4051 1896
rect 4045 1744 4051 1836
rect 4077 1763 4083 1936
rect 4141 1924 4147 2036
rect 4205 1984 4211 2197
rect 4237 2144 4243 2236
rect 4285 2124 4291 2136
rect 4285 2104 4291 2116
rect 4250 2014 4262 2016
rect 4235 2006 4237 2014
rect 4245 2006 4247 2014
rect 4255 2006 4257 2014
rect 4265 2006 4267 2014
rect 4275 2006 4277 2014
rect 4250 2004 4262 2006
rect 4189 1944 4195 1976
rect 4093 1883 4099 1916
rect 4109 1904 4115 1916
rect 4093 1877 4108 1883
rect 4109 1804 4115 1876
rect 4173 1864 4179 1896
rect 4189 1884 4195 1936
rect 4109 1764 4115 1796
rect 4077 1757 4092 1763
rect 4029 1684 4035 1696
rect 4029 1663 4035 1676
rect 4013 1657 4035 1663
rect 3965 1624 3971 1636
rect 3789 1504 3795 1556
rect 3709 1364 3715 1416
rect 3725 1364 3731 1436
rect 3741 1404 3747 1476
rect 3709 1344 3715 1356
rect 3741 1344 3747 1396
rect 3421 1124 3427 1176
rect 3645 1164 3651 1336
rect 3661 1324 3667 1336
rect 3693 1104 3699 1316
rect 3373 1017 3395 1023
rect 3373 904 3379 996
rect 3277 684 3283 696
rect 3245 564 3251 656
rect 3277 604 3283 636
rect 3325 544 3331 576
rect 3357 564 3363 636
rect 3373 624 3379 896
rect 3389 664 3395 1017
rect 3421 1004 3427 1096
rect 3549 964 3555 1056
rect 3725 1044 3731 1316
rect 3757 1104 3763 1336
rect 3773 1184 3779 1236
rect 3789 1224 3795 1356
rect 3709 1004 3715 1036
rect 3741 1024 3747 1076
rect 3421 844 3427 936
rect 3485 904 3491 916
rect 3533 824 3539 936
rect 3549 664 3555 956
rect 3677 944 3683 976
rect 3613 844 3619 900
rect 3581 684 3587 736
rect 3645 720 3651 758
rect 3677 704 3683 916
rect 3789 844 3795 916
rect 3549 644 3555 656
rect 3677 624 3683 696
rect 3437 524 3443 616
rect 3581 524 3587 536
rect 3597 524 3603 556
rect 3693 524 3699 696
rect 3725 684 3731 756
rect 3757 704 3763 736
rect 3773 724 3779 736
rect 3789 684 3795 796
rect 3805 704 3811 1576
rect 3821 1344 3827 1516
rect 3853 1483 3859 1496
rect 3853 1477 3868 1483
rect 3837 1324 3843 1456
rect 3821 1184 3827 1216
rect 3853 1143 3859 1336
rect 3837 1137 3859 1143
rect 3837 1084 3843 1137
rect 3853 1104 3859 1116
rect 3837 1004 3843 1056
rect 3853 724 3859 1036
rect 3869 904 3875 1476
rect 3901 1463 3907 1616
rect 3949 1484 3955 1536
rect 3997 1504 4003 1636
rect 4013 1524 4019 1657
rect 4013 1504 4019 1516
rect 3892 1457 3907 1463
rect 3901 1324 3907 1457
rect 3933 1364 3939 1456
rect 3965 1384 3971 1436
rect 3940 1357 3955 1363
rect 3901 1184 3907 1196
rect 3917 1123 3923 1236
rect 3901 1117 3923 1123
rect 3901 1084 3907 1117
rect 3933 1104 3939 1156
rect 3901 964 3907 1076
rect 3917 1064 3923 1096
rect 3933 1004 3939 1056
rect 3949 1044 3955 1357
rect 3981 1064 3987 1296
rect 3933 944 3939 996
rect 3853 704 3859 716
rect 3885 704 3891 876
rect 3917 744 3923 836
rect 3949 724 3955 1016
rect 3965 944 3971 1056
rect 4013 943 4019 1436
rect 4029 1244 4035 1636
rect 4045 1544 4051 1676
rect 4061 1504 4067 1596
rect 4077 1524 4083 1536
rect 4077 1504 4083 1516
rect 4109 1504 4115 1716
rect 4125 1504 4131 1856
rect 4173 1564 4179 1856
rect 4205 1523 4211 1976
rect 4301 1944 4307 2116
rect 4317 1864 4323 2276
rect 4333 2264 4339 2416
rect 4381 2404 4387 2716
rect 4413 2424 4419 2696
rect 4445 2624 4451 2716
rect 4461 2664 4467 2836
rect 4541 2784 4547 2856
rect 4797 2704 4803 2916
rect 4477 2604 4483 2636
rect 4509 2564 4515 2656
rect 4413 2384 4419 2396
rect 4349 2284 4355 2296
rect 4333 2224 4339 2256
rect 4381 2244 4387 2256
rect 4333 2184 4339 2216
rect 4349 2144 4355 2176
rect 4381 2164 4387 2236
rect 4413 2164 4419 2296
rect 4445 2283 4451 2376
rect 4445 2277 4460 2283
rect 4445 2164 4451 2277
rect 4493 2184 4499 2316
rect 4509 2284 4515 2456
rect 4541 2304 4547 2536
rect 4621 2524 4627 2696
rect 4733 2684 4739 2696
rect 4605 2462 4611 2500
rect 4653 2384 4659 2616
rect 4669 2483 4675 2616
rect 4685 2504 4691 2556
rect 4717 2524 4723 2536
rect 4733 2524 4739 2576
rect 4701 2504 4707 2516
rect 4749 2504 4755 2516
rect 4669 2477 4691 2483
rect 4557 2324 4563 2376
rect 4653 2304 4659 2316
rect 4596 2297 4611 2303
rect 4365 2124 4371 2156
rect 4349 1904 4355 2116
rect 4365 1944 4371 2116
rect 4413 2044 4419 2116
rect 4365 1904 4371 1916
rect 4413 1904 4419 2036
rect 4429 2004 4435 2116
rect 4461 2084 4467 2156
rect 4477 2144 4483 2156
rect 4493 2104 4499 2116
rect 4477 1984 4483 2096
rect 4333 1864 4339 1876
rect 4317 1804 4323 1856
rect 4381 1837 4396 1843
rect 4349 1764 4355 1836
rect 4250 1614 4262 1616
rect 4235 1606 4237 1614
rect 4245 1606 4247 1614
rect 4255 1606 4257 1614
rect 4265 1606 4267 1614
rect 4275 1606 4277 1614
rect 4250 1604 4262 1606
rect 4205 1517 4227 1523
rect 4125 1464 4131 1496
rect 4045 1124 4051 1436
rect 4141 1423 4147 1516
rect 4189 1484 4195 1496
rect 4157 1444 4163 1456
rect 4205 1444 4211 1496
rect 4141 1417 4163 1423
rect 4157 1344 4163 1417
rect 4221 1344 4227 1517
rect 4269 1364 4275 1476
rect 4077 1104 4083 1216
rect 4125 1104 4131 1336
rect 4221 1262 4227 1300
rect 4253 1264 4259 1316
rect 4250 1214 4262 1216
rect 4235 1206 4237 1214
rect 4245 1206 4247 1214
rect 4255 1206 4257 1214
rect 4265 1206 4267 1214
rect 4275 1206 4277 1214
rect 4250 1204 4262 1206
rect 4157 1103 4163 1156
rect 4205 1124 4211 1196
rect 4180 1117 4195 1123
rect 4189 1104 4195 1117
rect 4317 1104 4323 1196
rect 4333 1104 4339 1556
rect 4349 1543 4355 1756
rect 4381 1744 4387 1837
rect 4461 1784 4467 1936
rect 4477 1884 4483 1896
rect 4477 1724 4483 1816
rect 4493 1804 4499 1916
rect 4509 1904 4515 2256
rect 4525 2224 4531 2296
rect 4557 2144 4563 2296
rect 4605 2284 4611 2297
rect 4525 2124 4531 2136
rect 4445 1662 4451 1700
rect 4349 1537 4371 1543
rect 4365 1484 4371 1537
rect 4141 1097 4163 1103
rect 4029 944 4035 1036
rect 4077 944 4083 1036
rect 4125 1003 4131 1076
rect 4109 997 4131 1003
rect 4109 964 4115 997
rect 4004 937 4019 943
rect 3965 904 3971 936
rect 4029 864 4035 896
rect 3965 724 3971 836
rect 4013 704 4019 836
rect 3805 684 3811 696
rect 4045 664 4051 896
rect 4109 784 4115 956
rect 4125 904 4131 916
rect 3261 462 3267 500
rect 3437 304 3443 516
rect 3693 504 3699 516
rect 3501 320 3507 358
rect 3709 284 3715 656
rect 3949 644 3955 656
rect 3805 624 3811 636
rect 3725 544 3731 556
rect 3773 524 3779 616
rect 3917 604 3923 636
rect 3757 324 3763 376
rect 3773 304 3779 516
rect 3805 462 3811 500
rect 3901 443 3907 556
rect 3885 437 3907 443
rect 3357 184 3363 216
rect 3405 204 3411 256
rect 3437 224 3443 276
rect 3597 204 3603 236
rect 3549 164 3555 196
rect 3581 124 3587 136
rect 3677 124 3683 216
rect 3261 44 3267 116
rect 3325 104 3331 116
rect 3645 62 3651 100
rect 3709 44 3715 276
rect 3773 224 3779 296
rect 3885 264 3891 437
rect 3885 203 3891 256
rect 3876 197 3891 203
rect 3869 164 3875 196
rect 3869 144 3875 156
rect 3901 126 3907 216
rect 3965 124 3971 296
rect 3981 224 3987 656
rect 4029 284 4035 636
rect 4045 384 4051 636
rect 4061 584 4067 656
rect 4077 264 4083 336
rect 4093 144 4099 536
rect 4109 524 4115 536
rect 4125 524 4131 896
rect 4141 384 4147 1097
rect 4173 1077 4188 1083
rect 4173 984 4179 1077
rect 4237 1064 4243 1076
rect 4317 1044 4323 1076
rect 4333 1064 4339 1076
rect 4221 1024 4227 1036
rect 4317 984 4323 1036
rect 4157 964 4163 976
rect 4349 963 4355 1316
rect 4365 1304 4371 1356
rect 4413 1324 4419 1376
rect 4429 1344 4435 1396
rect 4381 1317 4396 1323
rect 4381 1104 4387 1317
rect 4445 1184 4451 1496
rect 4461 1364 4467 1516
rect 4509 1504 4515 1896
rect 4525 1724 4531 2116
rect 4541 1824 4547 1836
rect 4573 1823 4579 2256
rect 4589 2144 4595 2276
rect 4685 2223 4691 2477
rect 4781 2444 4787 2556
rect 4781 2304 4787 2316
rect 4797 2304 4803 2676
rect 4813 2664 4819 3036
rect 4877 2984 4883 3436
rect 4973 3383 4979 3496
rect 4957 3377 4979 3383
rect 4909 3044 4915 3236
rect 4957 3184 4963 3377
rect 4957 3104 4963 3176
rect 4925 3024 4931 3076
rect 4973 3064 4979 3296
rect 4989 3224 4995 3496
rect 5021 3444 5027 3736
rect 5037 3604 5043 3636
rect 5053 3584 5059 3696
rect 5085 3584 5091 3736
rect 5293 3724 5299 3756
rect 5140 3637 5155 3643
rect 5037 3384 5043 3496
rect 5085 3464 5091 3516
rect 5069 3444 5075 3456
rect 5069 3364 5075 3376
rect 5037 3344 5043 3356
rect 5021 3304 5027 3316
rect 5037 3284 5043 3336
rect 4989 3184 4995 3196
rect 5037 3064 5043 3096
rect 4829 2724 4835 2776
rect 4861 2724 4867 2956
rect 4925 2944 4931 2956
rect 4941 2924 4947 2976
rect 4733 2284 4739 2296
rect 4701 2244 4707 2256
rect 4749 2244 4755 2256
rect 4685 2217 4707 2223
rect 4605 2024 4611 2116
rect 4653 1984 4659 1996
rect 4685 1984 4691 2036
rect 4701 1984 4707 2217
rect 4733 2144 4739 2236
rect 4781 2124 4787 2296
rect 4797 2264 4803 2276
rect 4813 2184 4819 2636
rect 4829 2524 4835 2696
rect 4909 2664 4915 2916
rect 4973 2784 4979 3056
rect 5053 3024 5059 3236
rect 5069 3064 5075 3276
rect 5117 3204 5123 3476
rect 5149 3384 5155 3637
rect 5165 3424 5171 3436
rect 5149 3344 5155 3376
rect 5165 3364 5171 3416
rect 5229 3384 5235 3536
rect 5325 3464 5331 3716
rect 5389 3644 5395 3700
rect 5421 3504 5427 3716
rect 5453 3524 5459 3576
rect 5245 3364 5251 3416
rect 5165 3324 5171 3336
rect 5133 3284 5139 3296
rect 5149 3124 5155 3316
rect 5117 3083 5123 3096
rect 5101 3077 5123 3083
rect 5005 2984 5011 2996
rect 4989 2944 4995 2956
rect 5021 2944 5027 2976
rect 5037 2944 5043 2956
rect 5069 2924 5075 3036
rect 5101 2984 5107 3077
rect 5117 2944 5123 3016
rect 5133 2964 5139 3076
rect 5069 2897 5084 2903
rect 5069 2884 5075 2897
rect 5149 2684 5155 3036
rect 5165 2944 5171 3056
rect 5181 2964 5187 3316
rect 5213 3304 5219 3316
rect 5197 3104 5203 3296
rect 5213 3084 5219 3296
rect 5245 3184 5251 3316
rect 5325 3083 5331 3456
rect 5357 3423 5363 3476
rect 5341 3417 5363 3423
rect 5341 3384 5347 3417
rect 5357 3103 5363 3336
rect 5373 3324 5379 3376
rect 5453 3284 5459 3296
rect 5405 3124 5411 3276
rect 5357 3097 5372 3103
rect 5309 3077 5331 3083
rect 5261 3064 5267 3076
rect 5245 3004 5251 3056
rect 5309 2964 5315 3077
rect 5373 3044 5379 3096
rect 4909 2644 4915 2656
rect 5053 2644 5059 2656
rect 4957 2564 4963 2636
rect 4861 2462 4867 2500
rect 4829 2263 4835 2436
rect 4861 2284 4867 2356
rect 4829 2257 4844 2263
rect 4749 2104 4755 2116
rect 4589 1904 4595 1956
rect 4557 1817 4579 1823
rect 4557 1764 4563 1817
rect 4573 1744 4579 1796
rect 4605 1764 4611 1916
rect 4621 1884 4627 1916
rect 4637 1784 4643 1936
rect 4669 1884 4675 1896
rect 4749 1884 4755 2096
rect 4749 1784 4755 1876
rect 4765 1804 4771 2116
rect 4781 2064 4787 2096
rect 4893 2064 4899 2316
rect 4941 2284 4947 2336
rect 4909 2224 4915 2236
rect 4941 2204 4947 2276
rect 4957 2264 4963 2556
rect 5149 2544 5155 2556
rect 5165 2444 5171 2936
rect 5181 2724 5187 2776
rect 5197 2704 5203 2916
rect 5309 2824 5315 2956
rect 5341 2944 5347 3036
rect 5405 2862 5411 2900
rect 5277 2684 5283 2816
rect 5309 2702 5315 2796
rect 5277 2644 5283 2676
rect 4957 2203 4963 2256
rect 5053 2223 5059 2296
rect 5165 2284 5171 2296
rect 5229 2264 5235 2636
rect 5277 2544 5283 2636
rect 5357 2524 5363 2676
rect 5437 2603 5443 3036
rect 5437 2597 5459 2603
rect 5261 2324 5267 2376
rect 5309 2264 5315 2436
rect 5325 2303 5331 2496
rect 5357 2304 5363 2316
rect 5325 2297 5347 2303
rect 5341 2284 5347 2297
rect 5373 2284 5379 2316
rect 5405 2284 5411 2316
rect 5421 2304 5427 2518
rect 5373 2264 5379 2276
rect 5053 2217 5075 2223
rect 4957 2197 4979 2203
rect 4973 2164 4979 2197
rect 4813 2004 4819 2036
rect 4781 1824 4787 1896
rect 4893 1884 4899 1976
rect 4973 1904 4979 2116
rect 4989 1924 4995 1976
rect 5005 1924 5011 2136
rect 5069 2124 5075 2217
rect 5085 1984 5091 2216
rect 5133 2164 5139 2256
rect 5325 2204 5331 2236
rect 5101 2044 5107 2096
rect 5149 1984 5155 2176
rect 5181 2024 5187 2116
rect 5213 2062 5219 2100
rect 5053 1884 5059 1896
rect 4861 1844 4867 1856
rect 4877 1784 4883 1816
rect 4909 1764 4915 1796
rect 4605 1744 4611 1756
rect 4525 1604 4531 1716
rect 4525 1504 4531 1596
rect 4541 1524 4547 1636
rect 4557 1544 4563 1716
rect 4573 1704 4579 1736
rect 4621 1644 4627 1716
rect 4605 1637 4620 1643
rect 4573 1504 4579 1536
rect 4509 1384 4515 1436
rect 4541 1344 4547 1416
rect 4557 1324 4563 1496
rect 4589 1324 4595 1556
rect 4605 1524 4611 1637
rect 4621 1584 4627 1596
rect 4637 1584 4643 1736
rect 4653 1724 4659 1756
rect 4685 1684 4691 1756
rect 4701 1724 4707 1756
rect 4813 1724 4819 1736
rect 4717 1704 4723 1716
rect 4685 1664 4691 1676
rect 4621 1504 4627 1516
rect 4685 1464 4691 1636
rect 4701 1524 4707 1696
rect 4749 1664 4755 1676
rect 4765 1664 4771 1716
rect 4845 1684 4851 1716
rect 4861 1684 4867 1756
rect 4797 1524 4803 1676
rect 4909 1664 4915 1756
rect 4989 1744 4995 1876
rect 4957 1704 4963 1716
rect 4973 1704 4979 1716
rect 4973 1684 4979 1696
rect 4701 1484 4707 1516
rect 4717 1504 4723 1516
rect 4813 1504 4819 1576
rect 4877 1564 4883 1636
rect 4957 1604 4963 1636
rect 4877 1544 4883 1556
rect 4941 1504 4947 1536
rect 4957 1503 4963 1596
rect 4973 1584 4979 1656
rect 4957 1497 4972 1503
rect 4861 1464 4867 1496
rect 4637 1364 4643 1416
rect 4701 1344 4707 1436
rect 4829 1424 4835 1436
rect 4781 1344 4787 1416
rect 4493 1304 4499 1316
rect 4477 1284 4483 1296
rect 4541 1264 4547 1276
rect 4429 1144 4435 1176
rect 4381 964 4387 1076
rect 4413 1024 4419 1096
rect 4461 1044 4467 1096
rect 4477 1084 4483 1096
rect 4340 957 4355 963
rect 4157 924 4163 956
rect 4301 864 4307 956
rect 4461 944 4467 996
rect 4525 964 4531 1116
rect 4541 984 4547 1256
rect 4685 1244 4691 1296
rect 4701 1284 4707 1316
rect 4557 1104 4563 1196
rect 4573 1104 4579 1236
rect 4589 1084 4595 1096
rect 4365 864 4371 936
rect 4381 924 4387 936
rect 4413 924 4419 936
rect 4557 924 4563 976
rect 4397 884 4403 896
rect 4173 784 4179 856
rect 4413 844 4419 876
rect 4250 814 4262 816
rect 4235 806 4237 814
rect 4245 806 4247 814
rect 4255 806 4257 814
rect 4265 806 4267 814
rect 4275 806 4277 814
rect 4250 804 4262 806
rect 4189 524 4195 556
rect 4253 544 4259 716
rect 4365 684 4371 816
rect 4253 524 4259 536
rect 4157 484 4163 516
rect 4250 414 4262 416
rect 4235 406 4237 414
rect 4245 406 4247 414
rect 4255 406 4257 414
rect 4265 406 4267 414
rect 4275 406 4277 414
rect 4250 404 4262 406
rect 4205 324 4211 376
rect 4205 124 4211 296
rect 4301 284 4307 476
rect 4333 264 4339 656
rect 4429 584 4435 856
rect 4461 724 4467 776
rect 4477 744 4483 836
rect 4509 724 4515 736
rect 4541 704 4547 836
rect 4557 704 4563 896
rect 4573 784 4579 1076
rect 4589 944 4595 976
rect 4605 923 4611 1136
rect 4621 1124 4627 1236
rect 4813 1184 4819 1296
rect 4621 1063 4627 1096
rect 4621 1057 4636 1063
rect 4653 964 4659 1036
rect 4669 1004 4675 1076
rect 4717 1064 4723 1096
rect 4733 1084 4739 1116
rect 4845 1104 4851 1136
rect 4685 984 4691 1016
rect 4653 924 4659 936
rect 4605 917 4620 923
rect 4605 704 4611 836
rect 4349 537 4380 543
rect 4349 524 4355 537
rect 4365 504 4371 516
rect 4285 184 4291 216
rect 4333 164 4339 256
rect 4429 126 4435 516
rect 4477 484 4483 636
rect 4493 524 4499 656
rect 4541 624 4547 696
rect 4557 644 4563 696
rect 4653 684 4659 916
rect 4669 784 4675 936
rect 4685 723 4691 956
rect 4701 724 4707 1036
rect 4717 944 4723 1056
rect 4781 984 4787 1076
rect 4797 944 4803 1096
rect 4861 1084 4867 1096
rect 4813 1064 4819 1076
rect 4829 984 4835 1076
rect 4797 924 4803 936
rect 4877 924 4883 1136
rect 4893 1064 4899 1396
rect 4909 1104 4915 1456
rect 4925 1164 4931 1476
rect 4957 1124 4963 1497
rect 4989 1484 4995 1536
rect 5005 1523 5011 1856
rect 5037 1664 5043 1876
rect 5085 1824 5091 1896
rect 5069 1724 5075 1736
rect 5005 1517 5027 1523
rect 5021 1504 5027 1517
rect 4973 1384 4979 1456
rect 5005 1324 5011 1496
rect 5037 1424 5043 1436
rect 4973 1124 4979 1296
rect 5005 1144 5011 1316
rect 4909 1064 4915 1076
rect 5005 1064 5011 1096
rect 4973 1004 4979 1036
rect 5021 984 5027 1316
rect 5053 1264 5059 1716
rect 5085 1644 5091 1736
rect 5101 1724 5107 1876
rect 5117 1784 5123 1816
rect 5133 1744 5139 1896
rect 5149 1784 5155 1876
rect 5101 1584 5107 1656
rect 5117 1624 5123 1696
rect 5165 1544 5171 1916
rect 5181 1884 5187 1896
rect 5069 1504 5075 1536
rect 5085 1504 5091 1516
rect 5101 1484 5107 1516
rect 5181 1484 5187 1496
rect 5117 1464 5123 1476
rect 5101 1457 5116 1463
rect 5101 1344 5107 1457
rect 5149 1364 5155 1456
rect 5053 1144 5059 1236
rect 5101 1124 5107 1276
rect 5133 1104 5139 1136
rect 5149 1084 5155 1196
rect 5181 1184 5187 1476
rect 5197 1304 5203 1916
rect 5213 1584 5219 1836
rect 5229 1744 5235 2016
rect 5309 1904 5315 2156
rect 5277 1824 5283 1896
rect 5309 1764 5315 1896
rect 5405 1884 5411 2116
rect 5421 1984 5427 2136
rect 5389 1804 5395 1836
rect 5405 1743 5411 1876
rect 5421 1844 5427 1896
rect 5405 1737 5427 1743
rect 5037 1004 5043 1036
rect 5085 984 5091 1076
rect 5117 1064 5123 1076
rect 4717 744 4723 916
rect 4733 904 4739 916
rect 4676 717 4691 723
rect 4781 704 4787 896
rect 4845 744 4851 776
rect 4845 704 4851 736
rect 4877 704 4883 916
rect 5021 784 5027 936
rect 5085 862 5091 900
rect 5149 764 5155 1076
rect 4989 724 4995 756
rect 4973 704 4979 716
rect 4884 697 4899 703
rect 4509 524 4515 616
rect 4605 604 4611 656
rect 4669 604 4675 696
rect 4685 624 4691 656
rect 4717 584 4723 656
rect 4765 564 4771 696
rect 4493 384 4499 516
rect 4589 304 4595 556
rect 4621 544 4627 556
rect 4685 462 4691 500
rect 4653 302 4659 416
rect 4685 264 4691 276
rect 3901 117 3907 118
rect 4493 124 4499 256
rect 4589 124 4595 256
rect 4717 244 4723 256
rect 4733 124 4739 516
rect 4781 464 4787 696
rect 4829 664 4835 676
rect 4797 504 4803 636
rect 4877 604 4883 676
rect 4877 524 4883 596
rect 4893 524 4899 697
rect 4909 684 4915 696
rect 4941 584 4947 696
rect 5021 684 5027 696
rect 5037 684 5043 756
rect 4925 524 4931 556
rect 4973 544 4979 636
rect 5005 544 5011 576
rect 5037 544 5043 656
rect 4765 304 4771 336
rect 4781 323 4787 436
rect 4797 344 4803 496
rect 4877 384 4883 516
rect 4973 444 4979 516
rect 4781 317 4796 323
rect 4797 144 4803 236
rect 4829 164 4835 256
rect 4909 124 4915 296
rect 5021 284 5027 536
rect 5053 504 5059 636
rect 5069 584 5075 756
rect 5101 684 5107 736
rect 5069 544 5075 576
rect 5117 563 5123 636
rect 5149 584 5155 676
rect 5149 564 5155 576
rect 5117 557 5139 563
rect 5085 320 5091 358
rect 5101 304 5107 516
rect 5133 504 5139 557
rect 5181 304 5187 316
rect 4989 184 4995 236
rect 5021 164 5027 236
rect 5037 184 5043 216
rect 5101 124 5107 296
rect 5181 144 5187 276
rect 5213 264 5219 496
rect 5229 304 5235 1716
rect 5309 1502 5315 1503
rect 5245 1464 5251 1496
rect 5309 1444 5315 1494
rect 5325 1364 5331 1476
rect 5341 1404 5347 1736
rect 5405 1662 5411 1700
rect 5325 1243 5331 1356
rect 5357 1344 5363 1416
rect 5325 1237 5347 1243
rect 5341 1064 5347 1237
rect 5421 1204 5427 1737
rect 5437 1584 5443 2436
rect 5453 2304 5459 2597
rect 5469 2584 5475 3636
rect 5485 3444 5491 3756
rect 5485 2444 5491 3316
rect 5517 2684 5523 2696
rect 5517 2384 5523 2396
rect 5469 2264 5475 2296
rect 5501 1904 5507 2076
rect 5501 1884 5507 1896
rect 5453 1504 5459 1516
rect 5517 1484 5523 1496
rect 5437 1104 5443 1316
rect 5453 1244 5459 1296
rect 5469 1124 5475 1176
rect 5373 1064 5379 1076
rect 5341 964 5347 1056
rect 5341 843 5347 956
rect 5373 944 5379 996
rect 5453 924 5459 1096
rect 5437 844 5443 900
rect 5325 837 5347 843
rect 5325 664 5331 837
rect 5453 824 5459 916
rect 5421 704 5427 816
rect 5453 724 5459 776
rect 5357 664 5363 676
rect 5325 623 5331 656
rect 5309 617 5331 623
rect 5309 564 5315 617
rect 5309 504 5315 556
rect 5421 524 5427 696
rect 5405 462 5411 500
rect 5469 384 5475 496
rect 5277 304 5283 336
rect 5325 304 5331 316
rect 5213 164 5219 256
rect 4429 117 4435 118
rect 3997 44 4003 96
rect 4701 44 4707 96
rect 5085 44 5091 96
rect 5357 44 5363 276
rect 5517 84 5523 96
rect 3213 -23 3235 -17
rect 3261 -23 3267 16
rect 3293 -23 3299 36
rect 3517 -23 3523 16
rect 3725 -17 3731 36
rect 4250 14 4262 16
rect 4235 6 4237 14
rect 4245 6 4247 14
rect 4255 6 4257 14
rect 4265 6 4267 14
rect 4275 6 4277 14
rect 4250 4 4262 6
rect 4605 -17 4611 36
rect 4653 -17 4659 36
rect 3725 -23 3747 -17
rect 4589 -23 4611 -17
rect 4637 -23 4659 -17
rect 4701 -23 4707 16
rect 5165 -23 5171 36
rect 5437 -17 5443 36
rect 5421 -23 5443 -17
<< m3contact >>
rect 2060 3816 2068 3824
rect 3404 3816 3412 3824
rect 2723 3806 2731 3814
rect 2733 3806 2741 3814
rect 2743 3806 2751 3814
rect 2753 3806 2761 3814
rect 2763 3806 2771 3814
rect 2773 3806 2781 3814
rect 3484 3816 3492 3824
rect 3436 3796 3444 3804
rect 1964 3776 1972 3784
rect 2188 3776 2196 3784
rect 3276 3776 3284 3784
rect 188 3756 196 3764
rect 524 3756 532 3764
rect 892 3756 900 3764
rect 1340 3756 1348 3764
rect 220 3736 228 3744
rect 316 3716 324 3724
rect 380 3716 388 3724
rect 380 3576 388 3584
rect 444 3576 452 3584
rect 492 3576 500 3584
rect 220 3476 228 3484
rect 28 3436 36 3444
rect 188 3396 196 3404
rect 220 3396 228 3404
rect 428 3516 436 3524
rect 476 3516 484 3524
rect 444 3476 452 3484
rect 396 3436 404 3444
rect 252 3296 260 3304
rect 28 3176 36 3184
rect 12 3116 20 3124
rect 300 3216 308 3224
rect 172 3176 180 3184
rect 252 3176 260 3184
rect 316 3176 324 3184
rect 92 3136 100 3144
rect 124 3136 132 3144
rect 236 3136 244 3144
rect 60 3116 68 3124
rect 76 3096 84 3104
rect 188 3096 196 3104
rect 44 3056 52 3064
rect 28 2896 36 2904
rect 60 2896 68 2904
rect 236 3096 244 3104
rect 140 3056 148 3064
rect 220 3056 228 3064
rect 108 3036 116 3044
rect 188 2976 196 2984
rect 124 2956 132 2964
rect 188 2956 196 2964
rect 204 2956 212 2964
rect 380 3136 388 3144
rect 300 3076 308 3084
rect 348 3056 356 3064
rect 332 3036 340 3044
rect 332 2976 340 2984
rect 540 3516 548 3524
rect 508 3416 516 3424
rect 524 3396 532 3404
rect 732 3676 740 3684
rect 684 3636 692 3644
rect 732 3576 740 3584
rect 828 3496 836 3504
rect 684 3416 692 3424
rect 572 3376 580 3384
rect 492 3356 500 3364
rect 460 3336 468 3344
rect 524 3336 532 3344
rect 412 3316 420 3324
rect 572 3316 580 3324
rect 444 3296 452 3304
rect 428 3276 436 3284
rect 508 3296 516 3304
rect 588 3296 596 3304
rect 476 3256 484 3264
rect 524 3256 532 3264
rect 476 3156 484 3164
rect 524 3156 532 3164
rect 540 3156 548 3164
rect 604 3156 612 3164
rect 412 3136 420 3144
rect 428 3116 436 3124
rect 444 3116 452 3124
rect 364 2956 372 2964
rect 332 2936 340 2944
rect 108 2916 116 2924
rect 220 2916 228 2924
rect 140 2896 148 2904
rect 12 2556 20 2564
rect 44 2516 52 2524
rect 44 2296 52 2304
rect 188 2876 196 2884
rect 252 2876 260 2884
rect 188 2816 196 2824
rect 236 2776 244 2784
rect 220 2736 228 2744
rect 300 2756 308 2764
rect 284 2716 292 2724
rect 92 2556 100 2564
rect 140 2556 148 2564
rect 76 2516 84 2524
rect 124 2516 132 2524
rect 156 2516 164 2524
rect 108 2476 116 2484
rect 236 2576 244 2584
rect 204 2536 212 2544
rect 252 2536 260 2544
rect 236 2516 244 2524
rect 268 2516 276 2524
rect 188 2456 196 2464
rect 60 2216 68 2224
rect 220 2316 228 2324
rect 300 2676 308 2684
rect 316 2556 324 2564
rect 316 2516 324 2524
rect 188 2276 196 2284
rect 188 2256 196 2264
rect 220 2256 228 2264
rect 300 2236 308 2244
rect 156 2176 164 2184
rect 76 2156 84 2164
rect 172 2156 180 2164
rect 92 2136 100 2144
rect 156 2136 164 2144
rect 188 2136 196 2144
rect 124 2076 132 2084
rect 12 1876 20 1884
rect 60 1916 68 1924
rect 108 1916 116 1924
rect 44 1896 52 1904
rect 60 1896 68 1904
rect 44 1756 52 1764
rect 92 1856 100 1864
rect 140 1856 148 1864
rect 92 1756 100 1764
rect 108 1756 116 1764
rect 92 1716 100 1724
rect 44 1576 52 1584
rect 28 1516 36 1524
rect 76 1536 84 1544
rect 60 1516 68 1524
rect 12 1496 20 1504
rect 76 1496 84 1504
rect 28 1376 36 1384
rect 76 1376 84 1384
rect 76 1356 84 1364
rect 60 1336 68 1344
rect 44 1316 52 1324
rect 92 1316 100 1324
rect 172 2116 180 2124
rect 220 2196 228 2204
rect 284 2196 292 2204
rect 316 2196 324 2204
rect 268 2156 276 2164
rect 300 2156 308 2164
rect 268 2096 276 2104
rect 252 2076 260 2084
rect 396 3016 404 3024
rect 572 3136 580 3144
rect 444 3076 452 3084
rect 492 3076 500 3084
rect 428 2996 436 3004
rect 412 2956 420 2964
rect 380 2916 388 2924
rect 348 2876 356 2884
rect 380 2736 388 2744
rect 364 2716 372 2724
rect 380 2696 388 2704
rect 380 2676 388 2684
rect 364 2656 372 2664
rect 364 2536 372 2544
rect 348 2516 356 2524
rect 380 2476 388 2484
rect 508 3056 516 3064
rect 636 3316 644 3324
rect 668 3316 676 3324
rect 652 3276 660 3284
rect 700 3296 708 3304
rect 668 3116 676 3124
rect 556 3096 564 3104
rect 588 3096 596 3104
rect 620 3096 628 3104
rect 652 3096 660 3104
rect 540 3036 548 3044
rect 492 2996 500 3004
rect 572 2996 580 3004
rect 556 2956 564 2964
rect 444 2856 452 2864
rect 668 3056 676 3064
rect 652 3036 660 3044
rect 620 3016 628 3024
rect 668 3016 676 3024
rect 556 2816 564 2824
rect 924 3736 932 3744
rect 924 3656 932 3664
rect 972 3576 980 3584
rect 748 3436 756 3444
rect 892 3436 900 3444
rect 732 3376 740 3384
rect 1148 3656 1156 3664
rect 1612 3716 1620 3724
rect 1219 3606 1227 3614
rect 1229 3606 1237 3614
rect 1239 3606 1247 3614
rect 1249 3606 1257 3614
rect 1259 3606 1267 3614
rect 1269 3606 1277 3614
rect 1004 3496 1012 3504
rect 1228 3496 1236 3504
rect 1116 3476 1124 3484
rect 748 3356 756 3364
rect 796 3336 804 3344
rect 892 3336 900 3344
rect 828 3316 836 3324
rect 876 3316 884 3324
rect 908 3316 916 3324
rect 748 3296 756 3304
rect 860 3296 868 3304
rect 956 3376 964 3384
rect 1116 3416 1124 3424
rect 1148 3416 1156 3424
rect 972 3336 980 3344
rect 1404 3496 1412 3504
rect 1436 3496 1444 3504
rect 1292 3416 1300 3424
rect 1036 3296 1044 3304
rect 1148 3296 1156 3304
rect 940 3276 948 3284
rect 924 3256 932 3264
rect 716 3216 724 3224
rect 732 3136 740 3144
rect 732 3076 740 3084
rect 780 3076 788 3084
rect 956 3116 964 3124
rect 764 3056 772 3064
rect 796 3056 804 3064
rect 876 3056 884 3064
rect 748 3036 756 3044
rect 716 3016 724 3024
rect 700 2936 708 2944
rect 684 2916 692 2924
rect 748 2836 756 2844
rect 476 2756 484 2764
rect 476 2716 484 2724
rect 604 2716 612 2724
rect 652 2716 660 2724
rect 700 2716 708 2724
rect 412 2616 420 2624
rect 924 3056 932 3064
rect 908 2956 916 2964
rect 828 2916 836 2924
rect 524 2696 532 2704
rect 556 2696 564 2704
rect 636 2696 644 2704
rect 732 2696 740 2704
rect 492 2676 500 2684
rect 540 2676 548 2684
rect 604 2676 612 2684
rect 684 2676 692 2684
rect 748 2676 756 2684
rect 444 2656 452 2664
rect 556 2656 564 2664
rect 524 2636 532 2644
rect 428 2576 436 2584
rect 412 2556 420 2564
rect 444 2556 452 2564
rect 460 2556 468 2564
rect 428 2536 436 2544
rect 540 2536 548 2544
rect 396 2456 404 2464
rect 412 2456 420 2464
rect 396 2376 404 2384
rect 380 2356 388 2364
rect 380 2336 388 2344
rect 364 2296 372 2304
rect 492 2516 500 2524
rect 460 2476 468 2484
rect 476 2456 484 2464
rect 508 2496 516 2504
rect 572 2636 580 2644
rect 588 2496 596 2504
rect 572 2456 580 2464
rect 588 2456 596 2464
rect 460 2416 468 2424
rect 492 2416 500 2424
rect 444 2316 452 2324
rect 396 2276 404 2284
rect 380 2156 388 2164
rect 428 2216 436 2224
rect 364 2136 372 2144
rect 396 2136 404 2144
rect 492 2396 500 2404
rect 476 2296 484 2304
rect 508 2356 516 2364
rect 524 2356 532 2364
rect 508 2276 516 2284
rect 348 2116 356 2124
rect 396 2116 404 2124
rect 444 2116 452 2124
rect 476 2116 484 2124
rect 380 2096 388 2104
rect 380 2036 388 2044
rect 332 1996 340 2004
rect 316 1956 324 1964
rect 316 1936 324 1944
rect 220 1896 228 1904
rect 172 1880 180 1884
rect 172 1876 180 1880
rect 156 1696 164 1704
rect 140 1516 148 1524
rect 220 1856 228 1864
rect 204 1796 212 1804
rect 268 1876 276 1884
rect 284 1816 292 1824
rect 284 1796 292 1804
rect 236 1776 244 1784
rect 220 1756 228 1764
rect 204 1736 212 1744
rect 300 1736 308 1744
rect 188 1516 196 1524
rect 172 1496 180 1504
rect 348 1916 356 1924
rect 348 1876 356 1884
rect 332 1716 340 1724
rect 284 1636 292 1644
rect 252 1536 260 1544
rect 284 1496 292 1504
rect 204 1456 212 1464
rect 124 1416 132 1424
rect 204 1396 212 1404
rect 156 1356 164 1364
rect 188 1336 196 1344
rect 172 1316 180 1324
rect 284 1416 292 1424
rect 268 1316 276 1324
rect 284 1316 292 1324
rect 44 1216 52 1224
rect 220 1276 228 1284
rect 252 1276 260 1284
rect 220 1256 228 1264
rect 380 1756 388 1764
rect 364 1736 372 1744
rect 460 2096 468 2104
rect 428 2056 436 2064
rect 444 2056 452 2064
rect 428 2016 436 2024
rect 348 1636 356 1644
rect 364 1536 372 1544
rect 364 1516 372 1524
rect 316 1456 324 1464
rect 332 1376 340 1384
rect 364 1356 372 1364
rect 332 1336 340 1344
rect 540 2256 548 2264
rect 556 2196 564 2204
rect 684 2656 692 2664
rect 748 2656 756 2664
rect 620 2616 628 2624
rect 636 2556 644 2564
rect 732 2576 740 2584
rect 764 2556 772 2564
rect 812 2556 820 2564
rect 860 2676 868 2684
rect 876 2656 884 2664
rect 700 2536 708 2544
rect 748 2536 756 2544
rect 636 2516 644 2524
rect 668 2516 676 2524
rect 700 2516 708 2524
rect 652 2476 660 2484
rect 620 2456 628 2464
rect 604 2336 612 2344
rect 700 2376 708 2384
rect 684 2336 692 2344
rect 732 2396 740 2404
rect 764 2456 772 2464
rect 748 2376 756 2384
rect 732 2336 740 2344
rect 716 2316 724 2324
rect 604 2296 612 2304
rect 652 2296 660 2304
rect 620 2256 628 2264
rect 652 2176 660 2184
rect 636 2136 644 2144
rect 524 2096 532 2104
rect 508 2016 516 2024
rect 620 2076 628 2084
rect 636 2056 644 2064
rect 604 2016 612 2024
rect 636 2016 644 2024
rect 572 1976 580 1984
rect 540 1956 548 1964
rect 524 1936 532 1944
rect 492 1896 500 1904
rect 444 1856 452 1864
rect 476 1856 484 1864
rect 492 1856 500 1864
rect 428 1756 436 1764
rect 428 1736 436 1744
rect 428 1676 436 1684
rect 412 1656 420 1664
rect 460 1716 468 1724
rect 444 1616 452 1624
rect 428 1556 436 1564
rect 412 1476 420 1484
rect 396 1456 404 1464
rect 412 1336 420 1344
rect 348 1316 356 1324
rect 316 1276 324 1284
rect 332 1276 340 1284
rect 156 1156 164 1164
rect 204 1156 212 1164
rect 140 1136 148 1144
rect 188 1136 196 1144
rect 44 1116 52 1124
rect 60 1116 68 1124
rect 108 1116 116 1124
rect 172 1116 180 1124
rect 12 896 20 904
rect 44 1076 52 1084
rect 44 876 52 884
rect 28 656 36 664
rect 140 1096 148 1104
rect 76 1076 84 1084
rect 140 956 148 964
rect 156 936 164 944
rect 124 876 132 884
rect 76 736 84 744
rect 92 696 100 704
rect 60 676 68 684
rect 124 696 132 704
rect 156 896 164 904
rect 172 896 180 904
rect 300 1216 308 1224
rect 284 1136 292 1144
rect 252 1116 260 1124
rect 268 1116 276 1124
rect 316 1116 324 1124
rect 220 1096 228 1104
rect 380 1296 388 1304
rect 236 956 244 964
rect 204 916 212 924
rect 236 916 244 924
rect 220 896 228 904
rect 236 896 244 904
rect 188 876 196 884
rect 204 876 212 884
rect 156 816 164 824
rect 188 656 196 664
rect 108 576 116 584
rect 332 1056 340 1064
rect 316 1016 324 1024
rect 284 976 292 984
rect 268 916 276 924
rect 252 876 260 884
rect 300 936 308 944
rect 300 876 308 884
rect 332 976 340 984
rect 412 1276 420 1284
rect 412 1076 420 1084
rect 396 956 404 964
rect 444 1536 452 1544
rect 524 1836 532 1844
rect 588 1916 596 1924
rect 620 1996 628 2004
rect 636 1996 644 2004
rect 572 1856 580 1864
rect 524 1816 532 1824
rect 556 1816 564 1824
rect 540 1796 548 1804
rect 572 1776 580 1784
rect 492 1696 500 1704
rect 588 1636 596 1644
rect 572 1616 580 1624
rect 492 1596 500 1604
rect 508 1536 516 1544
rect 524 1516 532 1524
rect 508 1456 516 1464
rect 444 1296 452 1304
rect 476 1296 484 1304
rect 444 1016 452 1024
rect 604 1536 612 1544
rect 684 2176 692 2184
rect 780 2336 788 2344
rect 844 2336 852 2344
rect 876 2336 884 2344
rect 828 2316 836 2324
rect 796 2296 804 2304
rect 860 2296 868 2304
rect 796 2236 804 2244
rect 860 2236 868 2244
rect 780 2176 788 2184
rect 764 2116 772 2124
rect 716 2096 724 2104
rect 812 2096 820 2104
rect 748 2036 756 2044
rect 700 1996 708 2004
rect 732 1996 740 2004
rect 988 3096 996 3104
rect 1116 3276 1124 3284
rect 1068 3216 1076 3224
rect 1052 3136 1060 3144
rect 1084 3116 1092 3124
rect 1100 3116 1108 3124
rect 1219 3206 1227 3214
rect 1229 3206 1237 3214
rect 1239 3206 1247 3214
rect 1249 3206 1257 3214
rect 1259 3206 1267 3214
rect 1269 3206 1277 3214
rect 1292 3116 1300 3124
rect 1148 3096 1156 3104
rect 1212 3096 1220 3104
rect 1116 3056 1124 3064
rect 1084 2976 1092 2984
rect 1228 3056 1236 3064
rect 1196 2996 1204 3004
rect 1196 2976 1204 2984
rect 1516 3416 1524 3424
rect 2492 3756 2500 3764
rect 2732 3756 2740 3764
rect 3020 3756 3028 3764
rect 3148 3756 3156 3764
rect 1756 3716 1764 3724
rect 1724 3696 1732 3704
rect 1708 3476 1716 3484
rect 1564 3416 1572 3424
rect 1644 3416 1652 3424
rect 1532 3396 1540 3404
rect 1404 3296 1412 3304
rect 1596 3336 1604 3344
rect 1692 3336 1700 3344
rect 1516 3216 1524 3224
rect 1564 3216 1572 3224
rect 1596 3196 1604 3204
rect 1676 3196 1684 3204
rect 1484 3176 1492 3184
rect 1404 3136 1412 3144
rect 1308 3036 1316 3044
rect 1372 3116 1380 3124
rect 1356 3096 1364 3104
rect 1356 3056 1364 3064
rect 1340 2996 1348 3004
rect 1676 3176 1684 3184
rect 1644 3096 1652 3104
rect 1452 3076 1460 3084
rect 1564 3036 1572 3044
rect 1612 3056 1620 3064
rect 1532 2936 1540 2944
rect 1580 2936 1588 2944
rect 1596 2936 1604 2944
rect 1164 2916 1172 2924
rect 1260 2916 1268 2924
rect 1372 2916 1380 2924
rect 1420 2916 1428 2924
rect 1500 2916 1508 2924
rect 1548 2916 1556 2924
rect 1868 3696 1876 3704
rect 1772 3396 1780 3404
rect 2364 3736 2372 3744
rect 2428 3736 2436 3744
rect 2476 3736 2484 3744
rect 2284 3716 2292 3724
rect 2348 3716 2356 3724
rect 2156 3696 2164 3704
rect 2220 3696 2228 3704
rect 2268 3696 2276 3704
rect 2332 3696 2340 3704
rect 2460 3716 2468 3724
rect 1932 3616 1940 3624
rect 1996 3616 2004 3624
rect 2300 3676 2308 3684
rect 2332 3676 2340 3684
rect 2364 3676 2372 3684
rect 2444 3696 2452 3704
rect 2508 3676 2516 3684
rect 2396 3656 2404 3664
rect 2412 3656 2420 3664
rect 2524 3656 2532 3664
rect 2556 3656 2564 3664
rect 2188 3636 2196 3644
rect 2460 3636 2468 3644
rect 2540 3636 2548 3644
rect 2540 3576 2548 3584
rect 2156 3516 2164 3524
rect 2492 3556 2500 3564
rect 2540 3556 2548 3564
rect 2060 3496 2068 3504
rect 2092 3496 2100 3504
rect 2204 3496 2212 3504
rect 2428 3496 2436 3504
rect 1932 3456 1940 3464
rect 1932 3416 1940 3424
rect 1964 3416 1972 3424
rect 1996 3416 2004 3424
rect 1916 3396 1924 3404
rect 1948 3376 1956 3384
rect 1740 3316 1748 3324
rect 1756 3296 1764 3304
rect 1724 3176 1732 3184
rect 1756 3136 1764 3144
rect 1724 3116 1732 3124
rect 1772 3116 1780 3124
rect 1692 3096 1700 3104
rect 1692 3016 1700 3024
rect 1628 2976 1636 2984
rect 1644 2936 1652 2944
rect 1020 2836 1028 2844
rect 1084 2836 1092 2844
rect 1228 2896 1236 2904
rect 1324 2896 1332 2904
rect 1292 2876 1300 2884
rect 1219 2806 1227 2814
rect 1229 2806 1237 2814
rect 1239 2806 1247 2814
rect 1249 2806 1257 2814
rect 1259 2806 1267 2814
rect 1269 2806 1277 2814
rect 1148 2716 1156 2724
rect 1340 2836 1348 2844
rect 1356 2836 1364 2844
rect 1484 2876 1492 2884
rect 1452 2756 1460 2764
rect 1500 2736 1508 2744
rect 1452 2716 1460 2724
rect 1388 2696 1396 2704
rect 1036 2636 1044 2644
rect 908 2596 916 2604
rect 972 2596 980 2604
rect 1068 2596 1076 2604
rect 1004 2516 1012 2524
rect 1228 2676 1236 2684
rect 1196 2596 1204 2604
rect 1100 2476 1108 2484
rect 1148 2476 1156 2484
rect 1036 2396 1044 2404
rect 1020 2376 1028 2384
rect 1004 2356 1012 2364
rect 924 2296 932 2304
rect 1020 2276 1028 2284
rect 972 2236 980 2244
rect 956 2176 964 2184
rect 892 2136 900 2144
rect 924 2136 932 2144
rect 876 2116 884 2124
rect 924 2116 932 2124
rect 828 1976 836 1984
rect 972 2136 980 2144
rect 1340 2656 1348 2664
rect 1324 2556 1332 2564
rect 1212 2516 1220 2524
rect 1372 2616 1380 2624
rect 1420 2696 1428 2704
rect 1420 2636 1428 2644
rect 1404 2616 1412 2624
rect 1436 2556 1444 2564
rect 1228 2496 1236 2504
rect 1340 2476 1348 2484
rect 1219 2406 1227 2414
rect 1229 2406 1237 2414
rect 1239 2406 1247 2414
rect 1249 2406 1257 2414
rect 1259 2406 1267 2414
rect 1269 2406 1277 2414
rect 1052 2296 1058 2304
rect 1058 2296 1060 2304
rect 1356 2456 1364 2464
rect 1404 2476 1412 2484
rect 1388 2276 1396 2284
rect 1132 2236 1140 2244
rect 1244 2236 1252 2244
rect 1292 2136 1300 2144
rect 1004 2096 1012 2104
rect 988 1996 996 2004
rect 988 1976 996 1984
rect 668 1916 676 1924
rect 956 1956 964 1964
rect 988 1956 996 1964
rect 908 1916 916 1924
rect 652 1876 660 1884
rect 796 1876 804 1884
rect 732 1776 740 1784
rect 828 1776 836 1784
rect 924 1856 932 1864
rect 764 1756 772 1764
rect 860 1756 868 1764
rect 908 1756 916 1764
rect 636 1556 644 1564
rect 652 1516 660 1524
rect 588 1476 596 1484
rect 620 1476 628 1484
rect 652 1476 660 1484
rect 972 1716 980 1724
rect 956 1676 964 1684
rect 908 1616 916 1624
rect 668 1456 676 1464
rect 732 1456 740 1464
rect 716 1416 724 1424
rect 780 1356 788 1364
rect 588 1296 596 1304
rect 700 1336 708 1344
rect 572 1196 580 1204
rect 604 1196 612 1204
rect 668 1196 676 1204
rect 524 1076 532 1084
rect 700 1096 708 1104
rect 908 1476 916 1484
rect 876 1456 884 1464
rect 972 1436 980 1444
rect 892 1416 900 1424
rect 1004 1736 1012 1744
rect 1084 2096 1092 2104
rect 1052 2076 1060 2084
rect 1219 2006 1227 2014
rect 1229 2006 1237 2014
rect 1239 2006 1247 2014
rect 1249 2006 1257 2014
rect 1259 2006 1267 2014
rect 1269 2006 1277 2014
rect 1292 1920 1300 1924
rect 1292 1916 1300 1920
rect 1228 1876 1236 1884
rect 1628 2836 1636 2844
rect 1612 2736 1620 2744
rect 1564 2696 1572 2704
rect 1692 2876 1700 2884
rect 1676 2816 1684 2824
rect 1676 2736 1684 2744
rect 1660 2696 1668 2704
rect 1484 2676 1492 2684
rect 1516 2676 1524 2684
rect 1548 2676 1556 2684
rect 1628 2676 1636 2684
rect 1516 2636 1524 2644
rect 1676 2616 1684 2624
rect 1660 2596 1668 2604
rect 1580 2556 1588 2564
rect 1580 2536 1588 2544
rect 1612 2536 1620 2544
rect 1756 3056 1764 3064
rect 1868 3336 1876 3344
rect 1884 3296 1892 3304
rect 1820 3216 1828 3224
rect 1820 3176 1828 3184
rect 1820 3116 1828 3124
rect 1804 3096 1812 3104
rect 1932 3336 1940 3344
rect 2012 3336 2020 3344
rect 2060 3316 2068 3324
rect 1916 3176 1924 3184
rect 1804 3056 1812 3064
rect 1788 3016 1796 3024
rect 1740 2896 1748 2904
rect 1724 2836 1732 2844
rect 1708 2796 1716 2804
rect 1740 2776 1748 2784
rect 1788 2816 1796 2824
rect 1724 2736 1732 2744
rect 1756 2736 1764 2744
rect 1852 3016 1860 3024
rect 1868 2936 1876 2944
rect 1948 3096 1956 3104
rect 2044 3296 2052 3304
rect 2124 3296 2132 3304
rect 1996 3156 2004 3164
rect 2012 3116 2020 3124
rect 1916 3056 1924 3064
rect 2060 3216 2068 3224
rect 2124 3216 2132 3224
rect 2108 3176 2116 3184
rect 2092 3136 2100 3144
rect 2028 3096 2036 3104
rect 2284 3456 2292 3464
rect 2316 3436 2324 3444
rect 2956 3736 2964 3744
rect 3004 3736 3012 3744
rect 3196 3736 3204 3744
rect 2988 3716 2996 3724
rect 2972 3696 2980 3704
rect 2924 3636 2932 3644
rect 2988 3616 2996 3624
rect 3020 3596 3028 3604
rect 3052 3656 3060 3664
rect 3036 3556 3044 3564
rect 2812 3536 2820 3544
rect 3308 3756 3316 3764
rect 3356 3756 3364 3764
rect 3420 3756 3428 3764
rect 3100 3716 3108 3724
rect 3148 3716 3156 3724
rect 3180 3716 3188 3724
rect 3228 3716 3236 3724
rect 3132 3676 3140 3684
rect 3084 3656 3092 3664
rect 3068 3616 3076 3624
rect 3116 3656 3124 3664
rect 3100 3556 3108 3564
rect 3116 3536 3124 3544
rect 2508 3516 2516 3524
rect 2556 3516 2564 3524
rect 2668 3516 2676 3524
rect 2700 3516 2708 3524
rect 3036 3516 3044 3524
rect 2572 3476 2580 3484
rect 2652 3436 2660 3444
rect 2284 3356 2292 3364
rect 2364 3356 2372 3364
rect 2476 3356 2484 3364
rect 2204 3316 2212 3324
rect 2284 3316 2292 3324
rect 2140 3176 2148 3184
rect 2188 3136 2196 3144
rect 2156 3116 2164 3124
rect 2172 3116 2180 3124
rect 2332 3196 2340 3204
rect 2268 3176 2276 3184
rect 2140 3096 2148 3104
rect 1996 3016 2004 3024
rect 2028 3016 2036 3024
rect 1916 2936 1924 2944
rect 1916 2916 1924 2924
rect 1820 2876 1828 2884
rect 1932 2836 1940 2844
rect 1852 2796 1860 2804
rect 1804 2716 1812 2724
rect 1692 2516 1700 2524
rect 1500 2496 1508 2504
rect 1468 2456 1476 2464
rect 1580 2476 1588 2484
rect 1516 2416 1524 2424
rect 1500 2336 1508 2344
rect 1452 2316 1460 2324
rect 1612 2336 1620 2344
rect 1532 2316 1540 2324
rect 1580 2316 1588 2324
rect 1452 2256 1460 2264
rect 1468 2196 1476 2204
rect 1628 2316 1636 2324
rect 1660 2316 1668 2324
rect 1596 2296 1604 2304
rect 1580 2276 1588 2284
rect 1596 2216 1604 2224
rect 1628 2216 1636 2224
rect 1580 2136 1588 2144
rect 1596 2136 1604 2144
rect 1548 2116 1556 2124
rect 1772 2696 1780 2704
rect 1756 2676 1764 2684
rect 1740 2636 1748 2644
rect 1788 2656 1796 2664
rect 1820 2696 1828 2704
rect 1788 2636 1796 2644
rect 1772 2576 1780 2584
rect 1820 2476 1828 2484
rect 1772 2336 1780 2344
rect 1804 2336 1812 2344
rect 1708 2316 1716 2324
rect 1788 2316 1796 2324
rect 1692 2296 1700 2304
rect 1660 2276 1668 2284
rect 1740 2276 1748 2284
rect 1692 2236 1700 2244
rect 1724 2236 1732 2244
rect 1676 2196 1684 2204
rect 1756 2236 1764 2244
rect 1788 2256 1796 2264
rect 1788 2216 1796 2224
rect 1692 2136 1700 2144
rect 1612 2116 1620 2124
rect 1516 2096 1524 2104
rect 1660 2096 1668 2104
rect 1500 1996 1508 2004
rect 1420 1956 1428 1964
rect 1484 1916 1492 1924
rect 1196 1776 1204 1784
rect 1340 1776 1348 1784
rect 1052 1736 1060 1744
rect 1068 1716 1076 1724
rect 1219 1606 1227 1614
rect 1229 1606 1237 1614
rect 1239 1606 1247 1614
rect 1249 1606 1257 1614
rect 1259 1606 1267 1614
rect 1269 1606 1277 1614
rect 1196 1576 1204 1584
rect 1036 1556 1044 1564
rect 1084 1556 1092 1564
rect 1100 1556 1108 1564
rect 1020 1516 1028 1524
rect 1068 1516 1076 1524
rect 988 1416 996 1424
rect 844 1356 852 1364
rect 924 1356 932 1364
rect 860 1296 868 1304
rect 860 1216 868 1224
rect 828 1116 836 1124
rect 796 1076 804 1084
rect 844 1076 852 1084
rect 636 1056 644 1064
rect 812 1036 820 1044
rect 444 976 452 984
rect 460 976 468 984
rect 492 976 500 984
rect 396 916 404 924
rect 460 956 468 964
rect 412 896 420 904
rect 380 876 388 884
rect 364 716 372 724
rect 396 716 404 724
rect 220 696 228 704
rect 268 696 276 704
rect 284 696 292 704
rect 460 696 468 704
rect 252 636 260 644
rect 220 576 228 584
rect 44 556 52 564
rect 92 556 100 564
rect 124 556 132 564
rect 204 556 212 564
rect 12 536 20 544
rect 28 536 36 544
rect 44 536 52 544
rect 44 496 52 504
rect 108 536 116 544
rect 172 536 180 544
rect 236 536 244 544
rect 188 516 196 524
rect 268 516 276 524
rect 300 676 308 684
rect 316 676 324 684
rect 428 676 436 684
rect 796 956 804 964
rect 508 936 516 944
rect 588 936 596 944
rect 492 696 500 704
rect 828 916 836 924
rect 620 816 628 824
rect 652 816 660 824
rect 524 736 532 744
rect 588 716 596 724
rect 1148 1536 1156 1544
rect 1212 1556 1220 1564
rect 1196 1496 1204 1504
rect 1372 1736 1380 1744
rect 1468 1696 1476 1704
rect 1452 1556 1460 1564
rect 1356 1496 1364 1504
rect 1180 1456 1188 1464
rect 1164 1436 1172 1444
rect 1052 1416 1060 1424
rect 1020 1396 1028 1404
rect 972 1316 980 1324
rect 940 1216 948 1224
rect 1436 1436 1444 1444
rect 1116 1356 1124 1364
rect 1148 1356 1156 1364
rect 1340 1356 1348 1364
rect 1420 1356 1428 1364
rect 1116 1316 1124 1324
rect 1020 1176 1028 1184
rect 908 1116 916 1124
rect 876 1096 884 1104
rect 1004 1056 1012 1064
rect 972 1036 980 1044
rect 1228 1336 1236 1344
rect 1468 1436 1476 1444
rect 1164 1236 1172 1244
rect 1196 1216 1204 1224
rect 1219 1206 1227 1214
rect 1229 1206 1237 1214
rect 1239 1206 1247 1214
rect 1249 1206 1257 1214
rect 1259 1206 1267 1214
rect 1269 1206 1277 1214
rect 1164 1096 1172 1104
rect 1276 1096 1284 1104
rect 1308 1116 1316 1124
rect 1340 1116 1348 1124
rect 1532 1696 1540 1704
rect 1596 1856 1604 1864
rect 1676 1856 1684 1864
rect 1756 1996 1764 2004
rect 1884 2776 1892 2784
rect 1868 2736 1876 2744
rect 1900 2736 1908 2744
rect 1932 2736 1940 2744
rect 1980 2956 1988 2964
rect 1980 2936 1988 2944
rect 2012 2996 2020 3004
rect 2124 2956 2132 2964
rect 2044 2936 2052 2944
rect 1964 2916 1972 2924
rect 2028 2916 2036 2924
rect 2012 2896 2020 2904
rect 1996 2736 2004 2744
rect 1884 2696 1892 2704
rect 1932 2696 1940 2704
rect 1948 2696 1956 2704
rect 1980 2696 1988 2704
rect 1884 2636 1892 2644
rect 1852 2556 1860 2564
rect 1852 2396 1860 2404
rect 1884 2336 1892 2344
rect 1932 2656 1940 2664
rect 2076 2896 2084 2904
rect 2076 2776 2084 2784
rect 2060 2756 2068 2764
rect 2108 2736 2116 2744
rect 2028 2716 2036 2724
rect 2092 2716 2100 2724
rect 2028 2696 2036 2704
rect 2220 3096 2228 3104
rect 2300 3156 2308 3164
rect 2284 3116 2292 3124
rect 2204 3056 2212 3064
rect 2188 2956 2196 2964
rect 2396 3336 2404 3344
rect 2556 3336 2564 3344
rect 2444 3216 2452 3224
rect 2380 3176 2388 3184
rect 2364 3156 2372 3164
rect 2364 3096 2372 3104
rect 2380 3056 2388 3064
rect 2428 2976 2436 2984
rect 2140 2896 2148 2904
rect 2060 2656 2068 2664
rect 1932 2576 1940 2584
rect 2012 2576 2020 2584
rect 1948 2556 1956 2564
rect 2076 2576 2084 2584
rect 2236 2936 2244 2944
rect 2348 2956 2356 2964
rect 2316 2936 2324 2944
rect 2396 2936 2404 2944
rect 2204 2916 2212 2924
rect 2284 2916 2292 2924
rect 2364 2916 2372 2924
rect 2332 2896 2340 2904
rect 2316 2876 2324 2884
rect 2252 2796 2260 2804
rect 2252 2716 2260 2724
rect 2348 2736 2356 2744
rect 2492 3096 2500 3104
rect 2540 3096 2548 3104
rect 2476 3056 2484 3064
rect 2460 2976 2468 2984
rect 2412 2916 2420 2924
rect 2380 2736 2388 2744
rect 2268 2696 2276 2704
rect 2364 2696 2372 2704
rect 2444 2876 2452 2884
rect 2428 2736 2436 2744
rect 2316 2676 2324 2684
rect 2444 2676 2452 2684
rect 2108 2656 2116 2664
rect 2140 2656 2148 2664
rect 2204 2656 2212 2664
rect 2268 2656 2276 2664
rect 2140 2576 2148 2584
rect 2060 2556 2068 2564
rect 2092 2556 2100 2564
rect 2236 2556 2244 2564
rect 2236 2536 2244 2544
rect 2268 2536 2276 2544
rect 2348 2536 2356 2544
rect 2124 2416 2132 2424
rect 1948 2336 1956 2344
rect 1916 2316 1924 2324
rect 2028 2316 2036 2324
rect 2092 2316 2100 2324
rect 1916 2296 1924 2304
rect 1996 2296 2004 2304
rect 1980 2276 1988 2284
rect 1868 2236 1876 2244
rect 2044 2256 2052 2264
rect 1852 2216 1860 2224
rect 1964 2216 1972 2224
rect 1836 2156 1844 2164
rect 1996 2196 2004 2204
rect 1948 2156 1956 2164
rect 1884 2136 1892 2144
rect 1804 2116 1812 2124
rect 1836 2116 1844 2124
rect 1916 2116 1924 2124
rect 2012 2156 2020 2164
rect 1964 2136 1972 2144
rect 1996 2136 2004 2144
rect 1980 2116 1988 2124
rect 1916 2076 1924 2084
rect 2044 2116 2052 2124
rect 2124 2276 2132 2284
rect 2428 2656 2436 2664
rect 2412 2416 2420 2424
rect 2348 2296 2356 2304
rect 2508 3036 2516 3044
rect 2684 3496 2692 3504
rect 2972 3496 2974 3504
rect 2974 3496 2980 3504
rect 3068 3496 3076 3504
rect 3100 3496 3108 3504
rect 2668 3156 2676 3164
rect 2780 3456 2788 3464
rect 2812 3436 2820 3444
rect 2908 3436 2916 3444
rect 3068 3436 3076 3444
rect 2723 3406 2731 3414
rect 2733 3406 2741 3414
rect 2743 3406 2751 3414
rect 2753 3406 2761 3414
rect 2763 3406 2771 3414
rect 2773 3406 2781 3414
rect 2908 3376 2916 3384
rect 3084 3376 3092 3384
rect 3068 3256 3076 3264
rect 3068 3196 3076 3204
rect 2876 3176 2884 3184
rect 2588 3036 2596 3044
rect 2723 3006 2731 3014
rect 2733 3006 2741 3014
rect 2743 3006 2751 3014
rect 2753 3006 2761 3014
rect 2763 3006 2771 3014
rect 2773 3006 2781 3014
rect 2668 2956 2676 2964
rect 2492 2916 2500 2924
rect 2476 2896 2484 2904
rect 2540 2816 2548 2824
rect 2636 2916 2644 2924
rect 2668 2896 2676 2904
rect 2764 2836 2772 2844
rect 3276 3696 3284 3704
rect 3292 3696 3300 3704
rect 3212 3656 3220 3664
rect 3244 3576 3252 3584
rect 3212 3536 3220 3544
rect 3228 3536 3236 3544
rect 3148 3516 3156 3524
rect 3212 3516 3220 3524
rect 3148 3496 3156 3504
rect 3212 3496 3220 3504
rect 3228 3476 3236 3484
rect 3180 3456 3188 3464
rect 3260 3436 3268 3444
rect 3372 3736 3380 3744
rect 3404 3736 3412 3744
rect 3468 3736 3476 3744
rect 3372 3716 3380 3724
rect 3452 3716 3460 3724
rect 3340 3696 3348 3704
rect 3324 3676 3332 3684
rect 3468 3576 3476 3584
rect 3388 3536 3396 3544
rect 3372 3516 3380 3524
rect 3372 3496 3380 3504
rect 3292 3436 3300 3444
rect 3388 3476 3396 3484
rect 3420 3496 3428 3504
rect 3468 3496 3476 3504
rect 3340 3456 3348 3464
rect 3404 3456 3412 3464
rect 3276 3396 3284 3404
rect 3260 3376 3268 3384
rect 3100 3316 3108 3324
rect 3148 3216 3156 3224
rect 3180 3216 3188 3224
rect 3324 3196 3332 3204
rect 3308 3176 3316 3184
rect 3260 3136 3268 3144
rect 3228 3116 3236 3124
rect 3052 3016 3060 3024
rect 2924 2976 2932 2984
rect 2924 2956 2932 2964
rect 2956 2956 2964 2964
rect 2812 2796 2820 2804
rect 2956 2796 2964 2804
rect 2524 2716 2532 2724
rect 2556 2716 2564 2724
rect 2508 2696 2516 2704
rect 2540 2696 2548 2704
rect 2476 2656 2484 2664
rect 2492 2656 2500 2664
rect 2460 2616 2468 2624
rect 2252 2256 2260 2264
rect 2204 2216 2212 2224
rect 2444 2256 2452 2264
rect 2268 2196 2276 2204
rect 2380 2196 2388 2204
rect 2220 2156 2228 2164
rect 2236 2156 2244 2164
rect 2092 2136 2100 2144
rect 2204 2136 2212 2144
rect 2060 2096 2068 2104
rect 2028 2076 2036 2084
rect 1804 1976 1812 1984
rect 1836 1976 1844 1984
rect 1756 1896 1764 1904
rect 1916 1896 1924 1904
rect 1740 1816 1748 1824
rect 1644 1756 1652 1764
rect 1788 1736 1796 1744
rect 1644 1716 1652 1724
rect 1676 1716 1684 1724
rect 1612 1476 1620 1484
rect 1724 1456 1732 1464
rect 1612 1436 1620 1444
rect 1516 1336 1524 1344
rect 1612 1336 1620 1344
rect 1596 1316 1604 1324
rect 1628 1316 1636 1324
rect 1564 1296 1572 1304
rect 1596 1276 1604 1284
rect 1660 1336 1668 1344
rect 1676 1336 1684 1344
rect 1724 1336 1732 1344
rect 1692 1296 1700 1304
rect 1644 1216 1652 1224
rect 1596 1156 1604 1164
rect 1484 1096 1492 1104
rect 1148 1056 1156 1064
rect 1036 996 1044 1004
rect 1084 996 1092 1004
rect 876 956 884 964
rect 908 936 916 944
rect 1116 936 1124 944
rect 908 916 916 924
rect 956 916 964 924
rect 972 916 980 924
rect 1219 806 1227 814
rect 1229 806 1237 814
rect 1239 806 1247 814
rect 1249 806 1257 814
rect 1259 806 1267 814
rect 1269 806 1277 814
rect 844 736 852 744
rect 540 696 548 704
rect 780 696 788 704
rect 300 616 308 624
rect 300 556 308 564
rect 348 656 356 664
rect 396 656 404 664
rect 364 636 372 644
rect 380 636 388 644
rect 348 616 356 624
rect 444 636 452 644
rect 316 536 324 544
rect 156 496 164 504
rect 252 496 260 504
rect 220 396 228 404
rect 268 396 276 404
rect 204 376 212 384
rect 620 676 628 684
rect 748 676 756 684
rect 764 676 772 684
rect 492 596 500 604
rect 540 436 548 444
rect 572 436 580 444
rect 316 296 324 304
rect 460 296 468 304
rect 28 196 36 204
rect 92 196 100 204
rect 188 156 196 164
rect 220 136 228 144
rect 748 296 756 304
rect 572 276 580 284
rect 604 216 612 224
rect 668 216 676 224
rect 524 156 532 164
rect 492 136 500 144
rect 700 136 708 144
rect 684 116 686 124
rect 686 116 692 124
rect 876 696 884 704
rect 1308 696 1316 704
rect 1116 676 1124 684
rect 876 656 884 664
rect 1084 656 1092 664
rect 812 576 820 584
rect 796 296 804 304
rect 1036 556 1044 564
rect 924 236 932 244
rect 908 216 916 224
rect 940 216 948 224
rect 1004 216 1012 224
rect 876 156 884 164
rect 828 136 836 144
rect 1452 1076 1460 1084
rect 1484 1076 1492 1084
rect 1404 1056 1412 1064
rect 1404 1036 1412 1044
rect 1388 996 1396 1004
rect 1436 1016 1444 1024
rect 1372 956 1380 964
rect 1420 956 1428 964
rect 1468 1056 1476 1064
rect 1500 1016 1508 1024
rect 1356 936 1364 944
rect 1500 916 1508 924
rect 1548 1096 1556 1104
rect 1548 1076 1556 1084
rect 1644 1136 1652 1144
rect 1724 1296 1732 1304
rect 1676 1116 1684 1124
rect 1676 1096 1684 1104
rect 1708 1096 1716 1104
rect 1756 1496 1764 1504
rect 1804 1436 1812 1444
rect 2172 2096 2180 2104
rect 2140 2036 2148 2044
rect 2220 2116 2228 2124
rect 2332 2156 2340 2164
rect 2252 2096 2260 2104
rect 2188 1936 2196 1944
rect 2188 1896 2196 1904
rect 1932 1756 1940 1764
rect 1996 1756 2004 1764
rect 1868 1736 1876 1744
rect 2188 1876 2196 1884
rect 2236 1896 2244 1904
rect 2220 1856 2228 1864
rect 2236 1836 2244 1844
rect 2284 2076 2292 2084
rect 2284 2056 2292 2064
rect 2284 1936 2292 1944
rect 2332 2076 2340 2084
rect 2284 1916 2292 1924
rect 2316 1916 2324 1924
rect 2300 1876 2308 1884
rect 2348 1896 2356 1904
rect 2460 2116 2468 2124
rect 2396 2096 2404 2104
rect 2412 2096 2420 2104
rect 2396 2076 2404 2084
rect 2428 2076 2436 2084
rect 2300 1856 2308 1864
rect 2268 1816 2276 1824
rect 2220 1736 2228 1744
rect 2188 1716 2196 1724
rect 1964 1696 1972 1704
rect 1996 1696 2004 1704
rect 1836 1516 1844 1524
rect 1884 1516 1892 1524
rect 1788 1296 1796 1304
rect 2188 1636 2196 1644
rect 2012 1516 2020 1524
rect 1932 1496 1940 1504
rect 1836 1316 1842 1324
rect 1842 1316 1844 1324
rect 1932 1476 1940 1484
rect 2204 1616 2212 1624
rect 2044 1496 2052 1504
rect 2076 1496 2084 1504
rect 2060 1476 2068 1484
rect 2156 1476 2164 1484
rect 1948 1456 1956 1464
rect 2028 1456 2036 1464
rect 2076 1456 2084 1464
rect 2108 1456 2116 1464
rect 1852 1276 1860 1284
rect 1804 1156 1812 1164
rect 1788 1136 1796 1144
rect 1740 1076 1748 1084
rect 1836 1076 1844 1084
rect 1740 1056 1748 1064
rect 1772 1056 1780 1064
rect 1612 1036 1620 1044
rect 1756 1036 1764 1044
rect 1532 976 1540 984
rect 1740 976 1748 984
rect 2028 1336 2036 1344
rect 2188 1336 2196 1344
rect 2172 1316 2180 1324
rect 1964 1216 1972 1224
rect 1996 1216 2004 1224
rect 1932 1076 1940 1084
rect 2076 1056 2084 1064
rect 1884 996 1892 1004
rect 1532 916 1540 924
rect 1532 896 1540 904
rect 1612 896 1620 904
rect 1548 876 1556 884
rect 1340 796 1348 804
rect 1452 796 1460 804
rect 1628 716 1636 724
rect 1340 676 1348 684
rect 1532 676 1540 684
rect 1596 676 1604 684
rect 1324 596 1332 604
rect 1500 656 1508 664
rect 1484 616 1492 624
rect 1388 576 1396 584
rect 1356 556 1364 564
rect 1372 556 1380 564
rect 1436 556 1444 564
rect 1308 536 1316 544
rect 1228 516 1230 524
rect 1230 516 1236 524
rect 1219 406 1227 414
rect 1229 406 1237 414
rect 1239 406 1247 414
rect 1249 406 1257 414
rect 1259 406 1267 414
rect 1269 406 1277 414
rect 1148 296 1156 304
rect 1196 296 1204 304
rect 1196 236 1204 244
rect 1228 236 1236 244
rect 1068 216 1076 224
rect 1036 196 1044 204
rect 1212 196 1220 204
rect 1004 156 1012 164
rect 972 136 980 144
rect 796 116 804 124
rect 1164 116 1166 124
rect 1166 116 1172 124
rect 1452 516 1460 524
rect 1708 916 1716 924
rect 1756 916 1764 924
rect 1804 916 1812 924
rect 1676 716 1684 724
rect 1932 936 1940 944
rect 1852 856 1860 864
rect 1772 716 1780 724
rect 1644 656 1652 664
rect 1692 576 1700 584
rect 1708 576 1716 584
rect 1596 556 1604 564
rect 1548 516 1556 524
rect 1580 516 1588 524
rect 1628 536 1636 544
rect 1740 536 1748 544
rect 1628 516 1636 524
rect 1340 496 1348 504
rect 1356 336 1364 344
rect 1356 236 1364 244
rect 1772 496 1780 504
rect 1660 416 1668 424
rect 1692 416 1700 424
rect 1628 396 1636 404
rect 1660 396 1668 404
rect 1628 296 1636 304
rect 1532 236 1540 244
rect 1500 216 1508 224
rect 1548 216 1556 224
rect 1420 136 1428 144
rect 1580 136 1588 144
rect 1852 796 1860 804
rect 1932 796 1940 804
rect 1964 696 1972 704
rect 2092 976 2100 984
rect 2076 956 2084 964
rect 2044 936 2052 944
rect 1996 896 2004 904
rect 2044 876 2052 884
rect 2332 1796 2340 1804
rect 2300 1676 2308 1684
rect 2380 1876 2388 1884
rect 2348 1656 2356 1664
rect 2380 1736 2388 1744
rect 2380 1716 2388 1724
rect 2364 1636 2372 1644
rect 2380 1636 2388 1644
rect 2220 1496 2228 1504
rect 2252 1496 2260 1504
rect 2348 1476 2356 1484
rect 2412 1716 2420 1724
rect 2700 2676 2706 2684
rect 2706 2676 2708 2684
rect 2892 2676 2900 2684
rect 2588 2656 2596 2664
rect 2604 2656 2612 2664
rect 2892 2656 2900 2664
rect 2556 2636 2564 2644
rect 2723 2606 2731 2614
rect 2733 2606 2741 2614
rect 2743 2606 2751 2614
rect 2753 2606 2761 2614
rect 2763 2606 2771 2614
rect 2773 2606 2781 2614
rect 2524 2596 2532 2604
rect 2860 2596 2868 2604
rect 3068 2796 3076 2804
rect 3228 3096 3236 3104
rect 3308 3076 3316 3084
rect 3180 3016 3188 3024
rect 3228 3016 3236 3024
rect 3308 2976 3316 2984
rect 3116 2936 3124 2944
rect 3228 2916 3236 2924
rect 3276 2916 3284 2924
rect 3084 2656 3092 2664
rect 3052 2616 3060 2624
rect 3292 2876 3300 2884
rect 3196 2656 3204 2664
rect 3180 2616 3188 2624
rect 3276 2616 3284 2624
rect 3052 2596 3060 2604
rect 3100 2596 3108 2604
rect 3164 2596 3172 2604
rect 2636 2556 2644 2564
rect 2860 2556 2868 2564
rect 2764 2496 2772 2504
rect 2572 2416 2580 2424
rect 2636 2416 2644 2424
rect 2668 2416 2676 2424
rect 2492 2336 2500 2344
rect 2492 2296 2500 2304
rect 3228 2596 3236 2604
rect 3212 2556 3220 2564
rect 3180 2496 3188 2504
rect 3084 2396 3092 2404
rect 3020 2376 3028 2384
rect 3052 2376 3060 2384
rect 2764 2316 2772 2324
rect 2700 2296 2708 2304
rect 2764 2296 2772 2304
rect 2604 2276 2612 2284
rect 2828 2276 2836 2284
rect 3116 2320 3124 2324
rect 3116 2316 3124 2320
rect 2764 2256 2772 2264
rect 3052 2256 3060 2264
rect 2844 2216 2852 2224
rect 2723 2206 2731 2214
rect 2733 2206 2741 2214
rect 2743 2206 2751 2214
rect 2753 2206 2761 2214
rect 2763 2206 2771 2214
rect 2773 2206 2781 2214
rect 2572 2196 2580 2204
rect 2636 2196 2644 2204
rect 2508 2176 2516 2184
rect 2556 2176 2564 2184
rect 2476 2056 2484 2064
rect 2476 1916 2484 1924
rect 2444 1776 2452 1784
rect 2444 1756 2452 1764
rect 2460 1736 2468 1744
rect 2492 1856 2500 1864
rect 2764 2116 2772 2124
rect 2668 2096 2676 2104
rect 2556 2056 2564 2064
rect 2524 1896 2532 1904
rect 2588 2016 2596 2024
rect 2684 1896 2690 1904
rect 2690 1896 2692 1904
rect 2668 1876 2676 1884
rect 3020 2216 3028 2224
rect 3084 2216 3092 2224
rect 2892 2196 2900 2204
rect 2924 2156 2932 2164
rect 2860 2136 2868 2144
rect 3116 2136 3124 2144
rect 3228 2536 3236 2544
rect 3292 2536 3300 2544
rect 3292 2516 3300 2524
rect 3212 2296 3220 2304
rect 3276 2296 3284 2304
rect 3452 3476 3460 3484
rect 3452 3416 3460 3424
rect 3372 3396 3380 3404
rect 3420 3396 3428 3404
rect 3500 3796 3508 3804
rect 3420 3376 3428 3384
rect 3484 3376 3492 3384
rect 3436 3316 3444 3324
rect 3356 3136 3364 3144
rect 3372 3136 3380 3144
rect 3356 3096 3364 3104
rect 3404 3076 3412 3084
rect 3404 3056 3412 3064
rect 3468 3176 3476 3184
rect 3484 3136 3492 3144
rect 3484 3116 3492 3124
rect 3468 3096 3476 3104
rect 3484 3096 3492 3104
rect 3436 2996 3444 3004
rect 3468 3076 3476 3084
rect 3468 3036 3476 3044
rect 3452 2976 3460 2984
rect 3372 2936 3380 2944
rect 3468 2936 3476 2944
rect 3356 2896 3364 2904
rect 3404 2896 3412 2904
rect 3452 2896 3460 2904
rect 3436 2856 3444 2864
rect 3356 2736 3364 2744
rect 3388 2716 3396 2724
rect 3324 2696 3332 2704
rect 3372 2596 3380 2604
rect 3436 2696 3444 2704
rect 3404 2616 3412 2624
rect 3420 2596 3428 2604
rect 3404 2576 3412 2584
rect 3340 2536 3348 2544
rect 3388 2536 3396 2544
rect 3308 2356 3316 2364
rect 3308 2316 3316 2324
rect 3196 2276 3204 2284
rect 3228 2276 3236 2284
rect 3244 2276 3252 2284
rect 3196 2216 3204 2224
rect 3228 2216 3236 2224
rect 3180 2116 3188 2124
rect 2924 2036 2932 2044
rect 2956 1956 2964 1964
rect 2876 1876 2884 1884
rect 2620 1856 2628 1864
rect 2604 1796 2612 1804
rect 2572 1736 2580 1744
rect 2428 1616 2436 1624
rect 2460 1616 2468 1624
rect 2396 1576 2404 1584
rect 2524 1716 2532 1724
rect 2620 1716 2628 1724
rect 2508 1696 2516 1704
rect 2572 1696 2580 1704
rect 2332 1416 2340 1424
rect 2492 1416 2500 1424
rect 2284 1396 2292 1404
rect 2268 1336 2276 1344
rect 2556 1536 2564 1544
rect 2428 1356 2436 1364
rect 2460 1356 2468 1364
rect 2524 1356 2532 1364
rect 2380 1336 2388 1344
rect 2492 1336 2500 1344
rect 2524 1336 2532 1344
rect 2300 1316 2308 1324
rect 2332 1316 2340 1324
rect 2540 1316 2548 1324
rect 2204 1296 2212 1304
rect 2220 1296 2228 1304
rect 2140 1196 2148 1204
rect 2220 1176 2228 1184
rect 2140 1156 2148 1164
rect 2124 1116 2132 1124
rect 2204 1096 2212 1104
rect 2156 1076 2164 1084
rect 2252 1096 2260 1104
rect 2252 1056 2260 1064
rect 2220 996 2228 1004
rect 2188 976 2196 984
rect 2252 976 2260 984
rect 2332 1296 2340 1304
rect 2492 1296 2500 1304
rect 2460 1136 2468 1144
rect 2396 1116 2404 1124
rect 2476 1116 2484 1124
rect 2364 1096 2372 1104
rect 2332 1056 2340 1064
rect 2508 1176 2516 1184
rect 2524 1136 2532 1144
rect 2588 1656 2596 1664
rect 2604 1496 2612 1504
rect 2620 1476 2628 1484
rect 2572 1356 2580 1364
rect 2684 1836 2692 1844
rect 2668 1756 2676 1764
rect 2652 1736 2660 1744
rect 2700 1816 2708 1824
rect 2723 1806 2731 1814
rect 2733 1806 2741 1814
rect 2743 1806 2751 1814
rect 2753 1806 2761 1814
rect 2763 1806 2771 1814
rect 2773 1806 2781 1814
rect 2716 1776 2724 1784
rect 2732 1736 2740 1744
rect 2908 1756 2916 1764
rect 2828 1736 2836 1744
rect 2892 1736 2900 1744
rect 2700 1716 2708 1724
rect 2844 1716 2852 1724
rect 2652 1676 2660 1684
rect 2876 1696 2884 1704
rect 2924 1696 2932 1704
rect 2860 1676 2868 1684
rect 2908 1576 2916 1584
rect 2716 1536 2724 1544
rect 2796 1536 2804 1544
rect 2700 1496 2708 1504
rect 3292 2256 3300 2264
rect 3260 2196 3268 2204
rect 3260 2156 3268 2164
rect 3324 2296 3332 2304
rect 3884 3776 3892 3784
rect 4108 3756 4116 3764
rect 4540 3756 4548 3764
rect 4876 3756 4884 3764
rect 5292 3756 5300 3764
rect 3612 3736 3620 3744
rect 3516 3656 3524 3664
rect 3868 3736 3876 3744
rect 3932 3736 3940 3744
rect 3820 3716 3828 3724
rect 3916 3716 3924 3724
rect 3644 3636 3652 3644
rect 3612 3616 3620 3624
rect 3692 3616 3700 3624
rect 3724 3576 3732 3584
rect 3788 3556 3796 3564
rect 3756 3536 3764 3544
rect 3788 3536 3796 3544
rect 3532 3496 3540 3504
rect 3516 3476 3524 3484
rect 3516 3436 3524 3444
rect 3724 3496 3732 3504
rect 3740 3496 3748 3504
rect 3548 3396 3556 3404
rect 3564 3396 3572 3404
rect 3564 3356 3572 3364
rect 3532 3336 3540 3344
rect 3548 3316 3556 3324
rect 3516 3296 3524 3304
rect 3580 3296 3588 3304
rect 3596 3296 3604 3304
rect 3564 3256 3572 3264
rect 3532 3216 3540 3224
rect 3644 3456 3652 3464
rect 3660 3436 3668 3444
rect 3676 3436 3684 3444
rect 3644 3416 3652 3424
rect 3708 3436 3716 3444
rect 3628 3376 3636 3384
rect 3644 3356 3652 3364
rect 3740 3356 3748 3364
rect 3756 3356 3764 3364
rect 3628 3316 3636 3324
rect 3756 3316 3764 3324
rect 3596 3276 3604 3284
rect 3612 3276 3620 3284
rect 3756 3276 3764 3284
rect 3692 3236 3700 3244
rect 3708 3236 3716 3244
rect 3644 3216 3652 3224
rect 3660 3216 3668 3224
rect 3692 3216 3700 3224
rect 3612 3116 3620 3124
rect 3596 3096 3604 3104
rect 3532 3076 3540 3084
rect 3516 3056 3524 3064
rect 3756 3196 3764 3204
rect 3708 3136 3716 3144
rect 3756 3136 3764 3144
rect 3692 3076 3700 3084
rect 3644 3056 3652 3064
rect 3612 3036 3620 3044
rect 3628 3036 3636 3044
rect 3596 2976 3604 2984
rect 3756 3096 3764 3104
rect 3820 3576 3828 3584
rect 3884 3676 3892 3684
rect 3900 3676 3908 3684
rect 4076 3676 4084 3684
rect 3996 3656 4004 3664
rect 4268 3736 4270 3744
rect 4270 3736 4276 3744
rect 4460 3736 4468 3744
rect 4380 3716 4386 3724
rect 4386 3716 4388 3724
rect 4108 3636 4116 3644
rect 3900 3616 3908 3624
rect 3916 3616 3924 3624
rect 3948 3616 3956 3624
rect 4124 3616 4132 3624
rect 3884 3596 3892 3604
rect 3868 3556 3876 3564
rect 3836 3536 3844 3544
rect 3932 3596 3940 3604
rect 3980 3596 3988 3604
rect 4060 3596 4068 3604
rect 3964 3576 3972 3584
rect 3964 3516 3972 3524
rect 3852 3456 3860 3464
rect 4092 3556 4100 3564
rect 3996 3536 4004 3544
rect 4012 3536 4020 3544
rect 4060 3536 4068 3544
rect 4076 3536 4084 3544
rect 4028 3516 4036 3524
rect 3948 3436 3956 3444
rect 3964 3436 3972 3444
rect 4076 3516 4084 3524
rect 4044 3496 4052 3504
rect 4060 3496 4068 3504
rect 4012 3436 4020 3444
rect 3820 3376 3828 3384
rect 3996 3376 4004 3384
rect 3916 3356 3924 3364
rect 3980 3356 3988 3364
rect 3820 3316 3828 3324
rect 3788 3256 3796 3264
rect 3788 3096 3796 3104
rect 3836 3296 3844 3304
rect 3884 3296 3892 3304
rect 3948 3296 3956 3304
rect 3932 3236 3940 3244
rect 3996 3276 4004 3284
rect 4012 3256 4020 3264
rect 4227 3606 4235 3614
rect 4237 3606 4245 3614
rect 4247 3606 4255 3614
rect 4257 3606 4265 3614
rect 4267 3606 4275 3614
rect 4277 3606 4285 3614
rect 4412 3576 4420 3584
rect 4124 3536 4132 3544
rect 4844 3736 4852 3744
rect 5020 3736 5028 3744
rect 5068 3736 5076 3744
rect 5084 3736 5092 3744
rect 4636 3716 4644 3724
rect 4748 3716 4756 3724
rect 4956 3716 4964 3724
rect 4444 3536 4452 3544
rect 4492 3536 4500 3544
rect 4540 3536 4548 3544
rect 4204 3516 4212 3524
rect 4348 3516 4356 3524
rect 4396 3516 4404 3524
rect 4508 3516 4516 3524
rect 4620 3516 4628 3524
rect 4124 3496 4132 3504
rect 4220 3496 4228 3504
rect 4108 3476 4116 3484
rect 4204 3456 4212 3464
rect 4092 3436 4100 3444
rect 4108 3436 4116 3444
rect 4124 3376 4132 3384
rect 4172 3356 4180 3364
rect 4220 3356 4228 3364
rect 4092 3296 4100 3304
rect 4076 3276 4084 3284
rect 4044 3256 4052 3264
rect 4124 3236 4132 3244
rect 4076 3216 4084 3224
rect 4028 3196 4036 3204
rect 4092 3196 4100 3204
rect 3868 3136 3876 3144
rect 3980 3136 3988 3144
rect 4012 3136 4020 3144
rect 4060 3136 4068 3144
rect 3836 3116 3844 3124
rect 4076 3116 4084 3124
rect 3948 3096 3956 3104
rect 3996 3096 4004 3104
rect 3820 3076 3828 3084
rect 3852 3076 3860 3084
rect 3900 3076 3908 3084
rect 3756 3056 3764 3064
rect 3772 3056 3780 3064
rect 3724 3036 3732 3044
rect 3900 2996 3908 3004
rect 4060 3076 4068 3084
rect 4076 3076 4084 3084
rect 3996 3056 4004 3064
rect 4092 2996 4100 3004
rect 3740 2976 3748 2984
rect 3788 2976 3796 2984
rect 3836 2976 3844 2984
rect 3964 2976 3972 2984
rect 3980 2976 3988 2984
rect 3660 2956 3668 2964
rect 3692 2956 3700 2964
rect 3532 2936 3540 2944
rect 3500 2856 3508 2864
rect 3468 2716 3476 2724
rect 3484 2616 3492 2624
rect 3468 2556 3476 2564
rect 3452 2516 3460 2524
rect 3452 2476 3460 2484
rect 3356 2336 3364 2344
rect 3372 2316 3380 2324
rect 3388 2296 3396 2304
rect 3324 2276 3332 2284
rect 3340 2276 3348 2284
rect 3372 2276 3380 2284
rect 3388 2196 3396 2204
rect 3340 2156 3348 2164
rect 3324 2136 3332 2144
rect 3308 2116 3316 2124
rect 3356 2116 3364 2124
rect 3340 1956 3348 1964
rect 2972 1816 2980 1824
rect 3372 1936 3380 1944
rect 3372 1896 3380 1904
rect 3356 1856 3364 1864
rect 3388 1856 3396 1864
rect 3244 1816 3252 1824
rect 3324 1816 3332 1824
rect 3148 1776 3156 1784
rect 3228 1776 3236 1784
rect 3036 1756 3044 1764
rect 3324 1796 3332 1804
rect 3340 1756 3348 1764
rect 3116 1636 3124 1644
rect 3036 1516 3044 1524
rect 3292 1696 3300 1704
rect 3292 1516 3300 1524
rect 2812 1496 2820 1504
rect 2956 1496 2962 1504
rect 2962 1496 2964 1504
rect 2668 1476 2676 1484
rect 2876 1476 2884 1484
rect 3148 1476 3156 1484
rect 2620 1456 2628 1464
rect 2636 1456 2644 1464
rect 2668 1456 2676 1464
rect 2604 1336 2612 1344
rect 2636 1316 2644 1324
rect 2556 1096 2564 1104
rect 2460 1076 2468 1084
rect 2492 1076 2500 1084
rect 2508 1076 2516 1084
rect 2364 1056 2372 1064
rect 2396 1056 2404 1064
rect 2348 1016 2356 1024
rect 2220 956 2228 964
rect 2268 956 2276 964
rect 2348 956 2356 964
rect 2124 936 2132 944
rect 2188 936 2196 944
rect 2236 936 2244 944
rect 2252 936 2260 944
rect 2284 936 2292 944
rect 2316 936 2324 944
rect 2364 936 2372 944
rect 2124 896 2132 904
rect 2220 896 2228 904
rect 2268 896 2276 904
rect 2444 1056 2452 1064
rect 2428 956 2436 964
rect 2412 916 2420 924
rect 2604 1296 2612 1304
rect 3100 1416 3108 1424
rect 2723 1406 2731 1414
rect 2733 1406 2741 1414
rect 2743 1406 2751 1414
rect 2753 1406 2761 1414
rect 2763 1406 2771 1414
rect 2773 1406 2781 1414
rect 2732 1356 2740 1364
rect 2748 1276 2756 1284
rect 2668 1196 2676 1204
rect 2588 1096 2596 1104
rect 2572 1056 2580 1064
rect 2540 1036 2548 1044
rect 2460 996 2468 1004
rect 2508 1016 2516 1024
rect 2924 1336 2932 1344
rect 3068 1336 3076 1344
rect 3100 1316 3108 1324
rect 3068 1296 3076 1304
rect 2748 1096 2754 1104
rect 2754 1096 2756 1104
rect 2940 1076 2948 1084
rect 2908 1056 2916 1064
rect 2620 996 2628 1004
rect 2620 976 2628 984
rect 2492 956 2500 964
rect 2604 956 2612 964
rect 2476 916 2484 924
rect 2380 876 2388 884
rect 2284 796 2292 804
rect 2316 796 2324 804
rect 2108 696 2116 704
rect 2172 696 2180 704
rect 2476 736 2484 744
rect 1884 656 1892 664
rect 1980 656 1988 664
rect 2252 656 2260 664
rect 2140 596 2148 604
rect 2188 596 2196 604
rect 2300 596 2308 604
rect 1900 516 1908 524
rect 1804 496 1812 504
rect 2028 536 2036 544
rect 1852 416 1860 424
rect 1932 416 1940 424
rect 1788 396 1796 404
rect 1804 396 1812 404
rect 1948 396 1956 404
rect 2156 516 2164 524
rect 2220 516 2228 524
rect 2076 316 2084 324
rect 2188 316 2196 324
rect 2220 316 2228 324
rect 2124 296 2132 304
rect 2220 296 2228 304
rect 1884 276 1892 284
rect 2044 276 2052 284
rect 2348 556 2356 564
rect 2268 516 2276 524
rect 2364 516 2370 524
rect 2370 516 2372 524
rect 2252 496 2260 504
rect 2460 676 2468 684
rect 2428 656 2436 664
rect 2572 916 2580 924
rect 2604 816 2612 824
rect 2524 716 2532 724
rect 2572 716 2580 724
rect 2723 1006 2731 1014
rect 2733 1006 2741 1014
rect 2743 1006 2751 1014
rect 2753 1006 2761 1014
rect 2763 1006 2771 1014
rect 2773 1006 2781 1014
rect 2860 996 2868 1004
rect 2908 996 2916 1004
rect 2636 936 2644 944
rect 2636 856 2644 864
rect 2732 696 2740 704
rect 2892 936 2900 944
rect 3036 1036 3044 1044
rect 3084 976 3092 984
rect 3036 956 3044 964
rect 3068 956 3076 964
rect 2860 796 2868 804
rect 2908 796 2916 804
rect 2700 676 2708 684
rect 2620 656 2628 664
rect 2636 656 2644 664
rect 2668 656 2676 664
rect 2556 636 2564 644
rect 2492 596 2500 604
rect 2428 576 2436 584
rect 2556 556 2564 564
rect 2332 496 2340 504
rect 2396 496 2404 504
rect 2723 606 2731 614
rect 2733 606 2741 614
rect 2743 606 2751 614
rect 2753 606 2761 614
rect 2763 606 2771 614
rect 2773 606 2781 614
rect 2828 676 2836 684
rect 2620 500 2628 504
rect 2620 496 2628 500
rect 2796 496 2804 504
rect 2476 416 2484 424
rect 2524 416 2532 424
rect 2268 316 2276 324
rect 1852 216 1860 224
rect 1980 216 1988 224
rect 2028 216 2036 224
rect 2236 256 2244 264
rect 2268 256 2276 264
rect 1948 136 1956 144
rect 2236 136 2244 144
rect 2268 136 2276 144
rect 2252 116 2260 124
rect 1660 96 1668 104
rect 1852 96 1860 104
rect 2700 296 2708 304
rect 2812 296 2820 304
rect 2700 276 2708 284
rect 2796 276 2804 284
rect 2476 256 2484 264
rect 2348 236 2356 244
rect 2508 236 2516 244
rect 2332 216 2340 224
rect 2316 176 2324 184
rect 2444 216 2452 224
rect 2380 176 2388 184
rect 2396 156 2404 164
rect 2620 196 2628 204
rect 2460 176 2468 184
rect 2444 136 2452 144
rect 2716 236 2724 244
rect 2700 216 2708 224
rect 2668 196 2676 204
rect 2652 176 2660 184
rect 2668 176 2676 184
rect 2668 156 2676 164
rect 2556 136 2564 144
rect 2572 136 2580 144
rect 2636 136 2644 144
rect 2428 116 2436 124
rect 2556 116 2564 124
rect 2723 206 2731 214
rect 2733 206 2741 214
rect 2743 206 2751 214
rect 2753 206 2761 214
rect 2763 206 2771 214
rect 2773 206 2781 214
rect 2684 136 2692 144
rect 2796 136 2804 144
rect 2220 96 2228 104
rect 2300 96 2308 104
rect 2492 96 2500 104
rect 2540 96 2548 104
rect 2652 116 2660 124
rect 2716 116 2724 124
rect 2748 96 2756 104
rect 2780 96 2788 104
rect 2252 76 2260 84
rect 2284 76 2292 84
rect 2364 76 2372 84
rect 2396 76 2404 84
rect 2540 76 2548 84
rect 1219 6 1227 14
rect 1229 6 1237 14
rect 1239 6 1247 14
rect 1249 6 1257 14
rect 1259 6 1267 14
rect 1269 6 1277 14
rect 3212 1436 3220 1444
rect 3180 1396 3188 1404
rect 3148 1356 3156 1364
rect 3148 1316 3156 1324
rect 3164 1296 3172 1304
rect 3132 1116 3140 1124
rect 3116 1056 3124 1064
rect 3132 1036 3140 1044
rect 3100 816 3108 824
rect 3084 796 3092 804
rect 3052 756 3060 764
rect 2940 656 2948 664
rect 3196 1356 3204 1364
rect 3292 1476 3300 1484
rect 3436 2276 3444 2284
rect 3420 2256 3428 2264
rect 3420 2176 3428 2184
rect 3436 2176 3444 2184
rect 3468 2096 3476 2104
rect 3676 2936 3684 2944
rect 3772 2936 3780 2944
rect 3756 2916 3764 2924
rect 3772 2896 3780 2904
rect 3564 2876 3572 2884
rect 3724 2876 3732 2884
rect 3548 2756 3556 2764
rect 3548 2696 3556 2704
rect 3644 2656 3652 2664
rect 3612 2616 3620 2624
rect 3756 2596 3764 2604
rect 3628 2556 3636 2564
rect 3660 2556 3668 2564
rect 3548 2496 3556 2504
rect 3564 2416 3572 2424
rect 3644 2376 3652 2384
rect 3516 2356 3524 2364
rect 3612 2356 3620 2364
rect 3500 2256 3508 2264
rect 3420 1996 3428 2004
rect 3484 1996 3492 2004
rect 3452 1876 3460 1884
rect 3420 1856 3428 1864
rect 3436 1856 3444 1864
rect 3420 1776 3428 1784
rect 3372 1556 3380 1564
rect 3340 1536 3348 1544
rect 3420 1696 3428 1704
rect 3404 1516 3412 1524
rect 3372 1496 3380 1504
rect 3308 1456 3316 1464
rect 3452 1516 3460 1524
rect 3436 1496 3444 1504
rect 3436 1436 3444 1444
rect 3324 1416 3332 1424
rect 3388 1416 3396 1424
rect 3484 1756 3492 1764
rect 3484 1696 3492 1704
rect 3500 1676 3508 1684
rect 3596 2316 3604 2324
rect 3564 2296 3572 2304
rect 3532 2276 3540 2284
rect 3548 2176 3556 2184
rect 3660 2356 3668 2364
rect 3948 2936 3956 2944
rect 3836 2916 3844 2924
rect 3884 2896 3892 2904
rect 3820 2876 3828 2884
rect 3916 2876 3924 2884
rect 3964 2916 3972 2924
rect 4124 3076 4132 3084
rect 4364 3496 4372 3504
rect 4428 3496 4436 3504
rect 4492 3496 4500 3504
rect 4428 3456 4436 3464
rect 4364 3376 4372 3384
rect 4284 3256 4292 3264
rect 4227 3206 4235 3214
rect 4237 3206 4245 3214
rect 4247 3206 4255 3214
rect 4257 3206 4265 3214
rect 4267 3206 4275 3214
rect 4277 3206 4285 3214
rect 4300 3116 4308 3124
rect 4300 3056 4308 3064
rect 3996 2936 4004 2944
rect 3996 2896 4004 2904
rect 4076 2896 4084 2904
rect 4028 2876 4036 2884
rect 3804 2856 3812 2864
rect 3884 2856 3892 2864
rect 3932 2856 3940 2864
rect 3868 2696 3876 2704
rect 3804 2576 3812 2584
rect 3676 2316 3684 2324
rect 3708 2316 3716 2324
rect 3660 2296 3668 2304
rect 3708 2276 3716 2284
rect 3724 2256 3732 2264
rect 3740 2236 3748 2244
rect 3692 2196 3700 2204
rect 3708 2176 3716 2184
rect 3580 2096 3588 2104
rect 3676 2116 3684 2124
rect 3644 2076 3652 2084
rect 3724 2116 3732 2124
rect 3772 2296 3780 2304
rect 3788 2256 3796 2264
rect 3788 2236 3796 2244
rect 3804 2136 3812 2144
rect 3708 2076 3716 2084
rect 3756 2076 3764 2084
rect 3692 2036 3700 2044
rect 3596 1876 3604 1884
rect 3596 1856 3604 1864
rect 3532 1816 3540 1824
rect 3548 1776 3556 1784
rect 3532 1756 3540 1764
rect 3516 1576 3524 1584
rect 3516 1516 3524 1524
rect 3564 1736 3572 1744
rect 3628 1836 3636 1844
rect 4156 2956 4164 2964
rect 4140 2916 4148 2924
rect 4188 2916 4196 2924
rect 4220 2916 4228 2924
rect 4348 3316 4356 3324
rect 4412 3296 4420 3304
rect 4380 3236 4388 3244
rect 4348 3156 4356 3164
rect 4332 3096 4340 3104
rect 4316 3036 4324 3044
rect 4364 3116 4372 3124
rect 4412 3216 4420 3224
rect 4396 3076 4404 3084
rect 4396 3036 4404 3044
rect 4380 2976 4388 2984
rect 4364 2936 4372 2944
rect 4476 3396 4484 3404
rect 4444 3356 4452 3364
rect 4588 3496 4596 3504
rect 4620 3496 4628 3504
rect 4524 3476 4532 3484
rect 4540 3456 4548 3464
rect 4604 3436 4612 3444
rect 4556 3416 4564 3424
rect 4572 3416 4580 3424
rect 4876 3596 4884 3604
rect 4796 3576 4804 3584
rect 4732 3556 4740 3564
rect 4764 3556 4772 3564
rect 4748 3536 4756 3544
rect 4652 3516 4660 3524
rect 4652 3496 4660 3504
rect 4668 3476 4676 3484
rect 4716 3476 4724 3484
rect 4684 3456 4692 3464
rect 4732 3456 4740 3464
rect 4732 3416 4740 3424
rect 4700 3396 4708 3404
rect 4828 3536 4836 3544
rect 4780 3496 4788 3504
rect 4796 3496 4804 3504
rect 4844 3496 4852 3504
rect 4988 3556 4996 3564
rect 4924 3536 4932 3544
rect 4940 3536 4948 3544
rect 5004 3536 5012 3544
rect 4924 3496 4932 3504
rect 4972 3496 4980 3504
rect 4988 3496 4996 3504
rect 4876 3476 4884 3484
rect 4796 3456 4804 3464
rect 4652 3356 4660 3364
rect 4716 3336 4724 3344
rect 4476 3316 4484 3324
rect 4556 3316 4564 3324
rect 4460 3296 4468 3304
rect 4524 3276 4532 3284
rect 4428 3176 4436 3184
rect 4316 2916 4324 2924
rect 4332 2916 4340 2924
rect 4284 2856 4292 2864
rect 4227 2806 4235 2814
rect 4237 2806 4245 2814
rect 4247 2806 4255 2814
rect 4257 2806 4265 2814
rect 4267 2806 4275 2814
rect 4277 2806 4285 2814
rect 4220 2756 4228 2764
rect 4092 2696 4100 2704
rect 3964 2676 3972 2684
rect 4188 2696 4196 2704
rect 3996 2656 4004 2664
rect 4172 2656 4180 2664
rect 4300 2656 4308 2664
rect 3948 2556 3956 2564
rect 4060 2556 4068 2564
rect 3980 2276 3988 2284
rect 3852 2236 3860 2244
rect 3900 2216 3908 2224
rect 4028 2216 4036 2224
rect 3884 2176 3892 2184
rect 3996 2176 4004 2184
rect 3964 2156 3972 2164
rect 3852 2136 3860 2144
rect 3948 2136 3956 2144
rect 3916 2116 3924 2124
rect 3980 2116 3988 2124
rect 3820 2096 3828 2104
rect 3804 2076 3812 2084
rect 3804 2056 3812 2064
rect 3788 1976 3796 1984
rect 3884 2016 3892 2024
rect 4012 2136 4020 2144
rect 4188 2516 4196 2524
rect 4188 2436 4196 2444
rect 4732 3176 4740 3184
rect 4540 3076 4548 3084
rect 4444 3056 4452 3064
rect 4572 3056 4580 3064
rect 4780 3216 4788 3224
rect 4860 3436 4868 3444
rect 4876 3436 4884 3444
rect 4860 3296 4868 3304
rect 4844 3196 4852 3204
rect 4684 3056 4692 3064
rect 4748 3056 4756 3064
rect 4604 2996 4612 3004
rect 4652 2996 4660 3004
rect 4492 2936 4500 2944
rect 4716 2916 4724 2924
rect 4540 2856 4548 2864
rect 4460 2836 4468 2844
rect 4524 2836 4532 2844
rect 4348 2696 4356 2704
rect 4364 2676 4372 2684
rect 4332 2576 4340 2584
rect 4300 2536 4308 2544
rect 4316 2536 4324 2544
rect 4348 2536 4354 2544
rect 4354 2536 4356 2544
rect 4220 2496 4228 2504
rect 4316 2456 4324 2464
rect 4332 2416 4340 2424
rect 4227 2406 4235 2414
rect 4237 2406 4245 2414
rect 4247 2406 4255 2414
rect 4257 2406 4265 2414
rect 4267 2406 4275 2414
rect 4277 2406 4285 2414
rect 4204 2376 4212 2384
rect 4156 2316 4164 2324
rect 4188 2316 4196 2324
rect 4124 2256 4132 2264
rect 4108 2236 4116 2244
rect 4124 2236 4132 2244
rect 4140 2216 4148 2224
rect 4124 2176 4132 2184
rect 4108 2156 4116 2164
rect 4188 2276 4196 2284
rect 4172 2256 4180 2264
rect 4316 2336 4324 2344
rect 4284 2316 4292 2324
rect 4300 2296 4308 2304
rect 4316 2276 4324 2284
rect 4236 2236 4244 2244
rect 4028 2076 4036 2084
rect 3996 2036 4004 2044
rect 3900 1936 3908 1944
rect 3916 1936 3924 1944
rect 3948 1936 3956 1944
rect 3772 1916 3780 1924
rect 3788 1896 3790 1904
rect 3790 1896 3796 1904
rect 3884 1896 3892 1904
rect 3868 1876 3876 1884
rect 3804 1856 3812 1864
rect 3852 1856 3860 1864
rect 3804 1836 3812 1844
rect 3628 1776 3636 1784
rect 3676 1776 3684 1784
rect 3708 1776 3716 1784
rect 3564 1596 3572 1604
rect 3884 1816 3892 1824
rect 3756 1556 3764 1564
rect 3692 1536 3700 1544
rect 3628 1516 3636 1524
rect 3708 1516 3716 1524
rect 3500 1496 3508 1504
rect 3532 1496 3540 1504
rect 3564 1496 3572 1504
rect 3676 1496 3684 1504
rect 3484 1476 3492 1484
rect 3452 1396 3460 1404
rect 3484 1356 3492 1364
rect 3564 1356 3572 1364
rect 3356 1316 3364 1324
rect 3180 1116 3188 1124
rect 3164 1076 3172 1084
rect 3356 1296 3364 1304
rect 3212 1096 3220 1104
rect 3244 1056 3252 1064
rect 3196 996 3204 1004
rect 3276 936 3284 944
rect 3148 916 3156 924
rect 3132 736 3140 744
rect 3084 696 3092 704
rect 3100 696 3108 704
rect 3116 656 3124 664
rect 2940 636 2948 644
rect 3036 636 3044 644
rect 2908 596 2916 604
rect 2972 596 2980 604
rect 3260 836 3268 844
rect 3164 816 3172 824
rect 3148 696 3156 704
rect 3212 776 3220 784
rect 3260 756 3268 764
rect 3340 756 3348 764
rect 3180 696 3188 704
rect 3228 696 3236 704
rect 3212 676 3220 684
rect 3196 656 3204 664
rect 3212 636 3220 644
rect 2844 496 2852 504
rect 3148 496 3156 504
rect 2876 296 2884 304
rect 2860 276 2868 284
rect 2876 276 2884 284
rect 3084 276 3092 284
rect 3052 256 3060 264
rect 3068 196 3076 204
rect 2892 176 2900 184
rect 2908 116 2914 124
rect 2914 116 2916 124
rect 2876 96 2884 104
rect 3100 76 3108 84
rect 3180 536 3188 544
rect 3308 716 3316 724
rect 3372 1236 3380 1244
rect 3980 1896 3988 1904
rect 4012 1936 4020 1944
rect 4012 1916 4020 1924
rect 3996 1876 4004 1884
rect 4012 1876 4020 1884
rect 3948 1856 3956 1864
rect 3916 1776 3924 1784
rect 4012 1776 4020 1784
rect 4044 2056 4052 2064
rect 4092 2116 4100 2124
rect 4156 2116 4164 2124
rect 4124 2096 4132 2104
rect 4076 2076 4084 2084
rect 4108 2076 4116 2084
rect 4108 1996 4116 2004
rect 4172 2056 4180 2064
rect 4076 1936 4084 1944
rect 4124 1936 4132 1944
rect 4044 1896 4052 1904
rect 4060 1856 4068 1864
rect 4284 2096 4292 2104
rect 4227 2006 4235 2014
rect 4237 2006 4245 2014
rect 4247 2006 4255 2014
rect 4257 2006 4265 2014
rect 4267 2006 4275 2014
rect 4277 2006 4285 2014
rect 4188 1976 4196 1984
rect 4156 1936 4164 1944
rect 4188 1936 4196 1944
rect 4108 1916 4116 1924
rect 4140 1916 4148 1924
rect 4108 1876 4116 1884
rect 4124 1856 4132 1864
rect 4108 1796 4116 1804
rect 4044 1736 4052 1744
rect 4060 1716 4068 1724
rect 4108 1716 4116 1724
rect 3980 1676 3988 1684
rect 4028 1676 4036 1684
rect 3996 1636 4004 1644
rect 3900 1616 3908 1624
rect 3964 1616 3972 1624
rect 3804 1576 3812 1584
rect 3788 1556 3796 1564
rect 3788 1496 3796 1504
rect 3644 1476 3652 1484
rect 3708 1416 3716 1424
rect 3740 1396 3748 1404
rect 3612 1356 3620 1364
rect 3628 1356 3636 1364
rect 3708 1356 3716 1364
rect 3724 1356 3732 1364
rect 3612 1336 3620 1344
rect 3644 1336 3652 1344
rect 3660 1336 3668 1344
rect 3756 1336 3764 1344
rect 3596 1296 3604 1304
rect 3580 1196 3588 1204
rect 3676 1316 3684 1324
rect 3644 1156 3652 1164
rect 3692 1096 3700 1104
rect 3388 1056 3396 1064
rect 3372 996 3380 1004
rect 3356 696 3364 704
rect 3276 676 3284 684
rect 3244 656 3252 664
rect 3356 636 3364 644
rect 3276 596 3284 604
rect 3324 576 3332 584
rect 3244 556 3252 564
rect 3516 1076 3524 1084
rect 3548 1056 3556 1064
rect 3420 996 3428 1004
rect 3788 1216 3796 1224
rect 3772 1176 3780 1184
rect 3788 1096 3796 1104
rect 3772 1076 3780 1084
rect 3724 1036 3732 1044
rect 3740 1016 3748 1024
rect 3708 996 3716 1004
rect 3676 976 3684 984
rect 3548 956 3556 964
rect 3452 936 3460 944
rect 3532 936 3540 944
rect 3436 916 3444 924
rect 3484 916 3492 924
rect 3516 916 3524 924
rect 3420 836 3428 844
rect 3532 816 3540 824
rect 3708 956 3716 964
rect 3580 736 3588 744
rect 3788 836 3796 844
rect 3788 796 3796 804
rect 3724 756 3732 764
rect 3692 696 3700 704
rect 3388 656 3396 664
rect 3548 636 3556 644
rect 3372 616 3380 624
rect 3436 616 3444 624
rect 3676 616 3684 624
rect 3676 576 3684 584
rect 3548 556 3556 564
rect 3580 556 3588 564
rect 3580 536 3588 544
rect 3756 736 3764 744
rect 3772 736 3780 744
rect 3740 696 3748 704
rect 3820 1516 3828 1524
rect 3884 1516 3892 1524
rect 3836 1496 3844 1504
rect 3868 1496 3876 1504
rect 3868 1476 3876 1484
rect 3836 1456 3844 1464
rect 3820 1316 3828 1324
rect 3820 1216 3828 1224
rect 3852 1116 3860 1124
rect 3852 1036 3860 1044
rect 3836 996 3844 1004
rect 3948 1536 3956 1544
rect 3980 1536 3988 1544
rect 3932 1496 3940 1504
rect 3964 1516 3972 1524
rect 4012 1496 4020 1504
rect 3932 1456 3940 1464
rect 3964 1436 3972 1444
rect 4012 1436 4020 1444
rect 3884 1276 3892 1284
rect 3900 1196 3908 1204
rect 3932 1156 3940 1164
rect 3916 1056 3924 1064
rect 3980 1296 3988 1304
rect 3996 1076 4004 1084
rect 3964 1056 3972 1064
rect 3948 1036 3956 1044
rect 3948 1016 3956 1024
rect 3932 996 3940 1004
rect 3900 956 3908 964
rect 3900 916 3908 924
rect 3868 896 3876 904
rect 3900 896 3908 904
rect 3932 896 3940 904
rect 3852 716 3860 724
rect 3916 736 3924 744
rect 3964 936 3972 944
rect 3980 936 3988 944
rect 4076 1636 4084 1644
rect 4060 1596 4068 1604
rect 4044 1536 4052 1544
rect 4076 1536 4084 1544
rect 4092 1516 4100 1524
rect 4172 1556 4180 1564
rect 4140 1516 4148 1524
rect 4236 1916 4244 1924
rect 4412 2696 4420 2704
rect 4428 2696 4436 2704
rect 4396 2676 4404 2684
rect 4732 2696 4740 2704
rect 4492 2676 4500 2684
rect 4508 2656 4516 2664
rect 4444 2616 4452 2624
rect 4476 2596 4484 2604
rect 4508 2556 4516 2564
rect 4428 2516 4436 2524
rect 4508 2456 4516 2464
rect 4412 2416 4420 2424
rect 4380 2396 4388 2404
rect 4412 2396 4420 2404
rect 4444 2376 4452 2384
rect 4396 2336 4404 2344
rect 4412 2316 4420 2324
rect 4364 2296 4372 2304
rect 4348 2276 4356 2284
rect 4332 2256 4340 2264
rect 4380 2236 4388 2244
rect 4332 2216 4340 2224
rect 4348 2176 4356 2184
rect 4460 2316 4468 2324
rect 4796 2676 4804 2684
rect 4700 2656 4708 2664
rect 4652 2616 4660 2624
rect 4668 2616 4676 2624
rect 4732 2576 4740 2584
rect 4764 2536 4772 2544
rect 4716 2516 4724 2524
rect 4684 2496 4692 2504
rect 4700 2496 4708 2504
rect 4748 2496 4756 2504
rect 4556 2376 4564 2384
rect 4588 2376 4596 2384
rect 4604 2336 4612 2344
rect 4668 2336 4676 2344
rect 4572 2316 4580 2324
rect 4636 2316 4644 2324
rect 4652 2316 4660 2324
rect 4556 2296 4564 2304
rect 4508 2276 4516 2284
rect 4508 2256 4516 2264
rect 4492 2176 4500 2184
rect 4364 2156 4372 2164
rect 4444 2156 4452 2164
rect 4476 2156 4484 2164
rect 4348 2116 4356 2124
rect 4332 1916 4340 1924
rect 4412 2036 4420 2044
rect 4364 1936 4372 1944
rect 4364 1916 4372 1924
rect 4476 2096 4484 2104
rect 4492 2096 4500 2104
rect 4444 2076 4452 2084
rect 4460 2076 4468 2084
rect 4428 1996 4436 2004
rect 4492 2076 4500 2084
rect 4460 1936 4468 1944
rect 4348 1896 4356 1904
rect 4332 1876 4340 1884
rect 4316 1856 4324 1864
rect 4348 1836 4356 1844
rect 4316 1796 4324 1804
rect 4227 1606 4235 1614
rect 4237 1606 4245 1614
rect 4247 1606 4255 1614
rect 4257 1606 4265 1614
rect 4267 1606 4275 1614
rect 4277 1606 4285 1614
rect 4332 1556 4340 1564
rect 4076 1496 4084 1504
rect 4124 1456 4132 1464
rect 4028 1236 4036 1244
rect 4188 1476 4196 1484
rect 4156 1436 4164 1444
rect 4172 1436 4180 1444
rect 4204 1436 4212 1444
rect 4124 1356 4132 1364
rect 4236 1516 4244 1524
rect 4252 1496 4260 1504
rect 4268 1356 4276 1364
rect 4124 1336 4132 1344
rect 4220 1336 4228 1344
rect 4076 1216 4084 1224
rect 4044 1116 4052 1124
rect 4252 1256 4260 1264
rect 4227 1206 4235 1214
rect 4237 1206 4245 1214
rect 4247 1206 4255 1214
rect 4257 1206 4265 1214
rect 4267 1206 4275 1214
rect 4277 1206 4285 1214
rect 4204 1196 4212 1204
rect 4316 1196 4324 1204
rect 4156 1156 4164 1164
rect 4140 1116 4148 1124
rect 4124 1096 4132 1104
rect 4204 1116 4212 1124
rect 4476 1876 4484 1884
rect 4476 1816 4484 1824
rect 4460 1776 4468 1784
rect 4524 2216 4532 2224
rect 4588 2276 4596 2284
rect 4604 2276 4612 2284
rect 4572 2256 4580 2264
rect 4524 2136 4532 2144
rect 4540 2136 4548 2144
rect 4492 1796 4500 1804
rect 4460 1516 4468 1524
rect 4428 1396 4436 1404
rect 4412 1376 4420 1384
rect 4060 1076 4068 1084
rect 4044 1056 4052 1064
rect 4092 976 4100 984
rect 4108 956 4116 964
rect 4028 936 4036 944
rect 4044 936 4052 944
rect 4076 936 4084 944
rect 3964 896 3972 904
rect 4044 896 4052 904
rect 4076 896 4084 904
rect 4028 856 4036 864
rect 3916 716 3924 724
rect 3964 716 3972 724
rect 3884 696 3892 704
rect 3804 676 3812 684
rect 3868 676 3876 684
rect 3932 676 3940 684
rect 3996 676 4004 684
rect 4124 896 4132 904
rect 3708 656 3716 664
rect 3548 516 3556 524
rect 3596 516 3604 524
rect 3644 516 3652 524
rect 3692 516 3700 524
rect 3692 496 3700 504
rect 3244 296 3250 304
rect 3250 296 3252 304
rect 3948 636 3956 644
rect 3772 616 3780 624
rect 3804 616 3812 624
rect 3724 556 3732 564
rect 3916 596 3924 604
rect 3868 536 3876 544
rect 3356 216 3364 224
rect 3436 216 3444 224
rect 3676 216 3684 224
rect 3404 196 3412 204
rect 3548 196 3556 204
rect 3596 196 3604 204
rect 3244 136 3252 144
rect 3308 136 3316 144
rect 3292 116 3300 124
rect 3580 116 3588 124
rect 3324 96 3332 104
rect 3388 96 3396 104
rect 3852 276 3860 284
rect 3772 216 3780 224
rect 3868 196 3876 204
rect 3900 216 3908 224
rect 3868 156 3876 164
rect 4044 636 4052 644
rect 4108 536 4116 544
rect 4076 336 4084 344
rect 4028 276 4036 284
rect 3980 216 3988 224
rect 4124 516 4132 524
rect 4172 1096 4180 1104
rect 4316 1096 4324 1104
rect 4236 1076 4244 1084
rect 4332 1076 4340 1084
rect 4316 1036 4324 1044
rect 4220 1016 4228 1024
rect 4156 976 4164 984
rect 4428 1336 4436 1344
rect 4364 1296 4372 1304
rect 4396 1316 4404 1324
rect 4540 1816 4548 1824
rect 4780 2436 4788 2444
rect 4764 2316 4772 2324
rect 4780 2316 4788 2324
rect 4940 3296 4948 3304
rect 4972 3316 4980 3324
rect 4956 3096 4964 3104
rect 4908 3036 4916 3044
rect 5052 3696 5060 3704
rect 5036 3596 5044 3604
rect 5068 3676 5076 3684
rect 5324 3736 5332 3744
rect 5212 3716 5220 3724
rect 5292 3716 5300 3724
rect 5324 3716 5332 3724
rect 5100 3696 5108 3704
rect 5084 3516 5092 3524
rect 5020 3436 5028 3444
rect 5132 3496 5140 3504
rect 5068 3436 5076 3444
rect 5036 3376 5044 3384
rect 5068 3376 5076 3384
rect 5036 3356 5044 3364
rect 5084 3336 5092 3344
rect 5020 3296 5028 3304
rect 5100 3316 5108 3324
rect 5036 3276 5044 3284
rect 5068 3276 5076 3284
rect 4988 3216 4996 3224
rect 4988 3196 4996 3204
rect 4940 3056 4948 3064
rect 4972 3056 4980 3064
rect 5036 3056 5044 3064
rect 4924 3016 4932 3024
rect 4940 2976 4948 2984
rect 4924 2956 4932 2964
rect 4892 2936 4900 2944
rect 4956 2916 4964 2924
rect 4892 2776 4900 2784
rect 4860 2716 4868 2724
rect 4828 2696 4836 2704
rect 4812 2656 4820 2664
rect 4812 2636 4820 2644
rect 4796 2296 4804 2304
rect 4700 2276 4708 2284
rect 4732 2276 4740 2284
rect 4700 2236 4708 2244
rect 4732 2236 4740 2244
rect 4748 2236 4756 2244
rect 4620 2136 4628 2144
rect 4636 2116 4644 2124
rect 4652 2116 4660 2124
rect 4604 2016 4612 2024
rect 4652 1996 4660 2004
rect 4796 2256 4804 2264
rect 5228 3536 5236 3544
rect 5164 3416 5172 3424
rect 5148 3376 5156 3384
rect 5244 3416 5252 3424
rect 5228 3376 5236 3384
rect 5164 3356 5172 3364
rect 5212 3356 5220 3364
rect 5164 3336 5172 3344
rect 5244 3316 5252 3324
rect 5308 3316 5316 3324
rect 5132 3276 5140 3284
rect 5116 3196 5124 3204
rect 5100 3096 5108 3104
rect 5116 3096 5124 3104
rect 5084 3076 5092 3084
rect 5068 3036 5076 3044
rect 5052 3016 5060 3024
rect 5004 2996 5012 3004
rect 5020 2976 5028 2984
rect 4988 2956 4996 2964
rect 5036 2936 5044 2944
rect 5132 3076 5140 3084
rect 5116 3016 5124 3024
rect 5100 2976 5108 2984
rect 4988 2916 4996 2924
rect 4972 2776 4980 2784
rect 4972 2696 4980 2704
rect 5212 3296 5220 3304
rect 5308 3096 5316 3104
rect 5212 3076 5220 3084
rect 5260 3076 5268 3084
rect 5292 3076 5300 3084
rect 5372 3376 5380 3384
rect 5356 3336 5364 3344
rect 5340 3296 5348 3304
rect 5340 3116 5348 3124
rect 5436 3356 5444 3364
rect 5372 3296 5380 3304
rect 5452 3296 5460 3304
rect 5404 3276 5412 3284
rect 5372 3116 5380 3124
rect 5420 3116 5428 3124
rect 5244 2996 5252 3004
rect 5356 3076 5364 3084
rect 5372 3036 5380 3044
rect 5180 2956 5188 2964
rect 5164 2936 5172 2944
rect 5084 2676 5092 2684
rect 5148 2676 5156 2684
rect 4908 2656 4916 2664
rect 4908 2636 4916 2644
rect 4956 2636 4964 2644
rect 5052 2636 5060 2644
rect 5148 2556 5156 2564
rect 4924 2536 4932 2544
rect 4828 2436 4836 2444
rect 4860 2356 4868 2364
rect 4844 2296 4852 2304
rect 4940 2336 4948 2344
rect 4876 2316 4884 2324
rect 4716 2116 4724 2124
rect 4780 2116 4788 2124
rect 4748 2096 4756 2104
rect 4684 1976 4692 1984
rect 4588 1956 4596 1964
rect 4604 1936 4612 1944
rect 4636 1936 4644 1944
rect 4588 1876 4596 1884
rect 4572 1796 4580 1804
rect 4620 1876 4628 1884
rect 4652 1896 4660 1904
rect 4668 1896 4676 1904
rect 4748 1876 4756 1884
rect 4908 2216 4916 2224
rect 5116 2516 5118 2524
rect 5118 2516 5124 2524
rect 5196 2916 5204 2924
rect 5228 2916 5236 2924
rect 5276 2816 5284 2824
rect 5308 2816 5316 2824
rect 5308 2796 5316 2804
rect 5244 2656 5252 2664
rect 5276 2636 5284 2644
rect 5164 2436 5172 2444
rect 5164 2296 5172 2304
rect 4972 2276 4978 2284
rect 4978 2276 4980 2284
rect 4956 2256 4964 2264
rect 4940 2196 4948 2204
rect 5308 2436 5316 2444
rect 5356 2316 5364 2324
rect 5404 2316 5412 2324
rect 5436 2436 5444 2444
rect 5132 2256 5140 2264
rect 5228 2256 5236 2264
rect 5372 2256 5380 2264
rect 5420 2256 5428 2264
rect 4972 2116 4980 2124
rect 4780 2056 4788 2064
rect 4892 2056 4900 2064
rect 4812 1996 4820 2004
rect 4892 1976 4900 1984
rect 5084 2216 5092 2224
rect 5068 2116 5076 2124
rect 5372 2236 5380 2244
rect 5324 2196 5332 2204
rect 5148 2176 5156 2184
rect 5132 2156 5140 2164
rect 5308 2156 5316 2164
rect 5276 2136 5284 2144
rect 5180 2116 5188 2124
rect 5180 2016 5188 2024
rect 5228 2016 5236 2024
rect 5004 1916 5012 1924
rect 5164 1916 5172 1924
rect 5196 1916 5204 1924
rect 5116 1896 5124 1904
rect 5132 1896 5140 1904
rect 4988 1876 4996 1884
rect 5052 1876 5060 1884
rect 4860 1836 4868 1844
rect 4780 1816 4788 1824
rect 4876 1816 4884 1824
rect 4764 1796 4772 1804
rect 4908 1796 4916 1804
rect 4604 1756 4612 1764
rect 4684 1756 4692 1764
rect 4700 1756 4708 1764
rect 4860 1756 4868 1764
rect 4636 1736 4644 1744
rect 4524 1596 4532 1604
rect 4572 1696 4580 1704
rect 4588 1556 4596 1564
rect 4556 1536 4564 1544
rect 4540 1516 4548 1524
rect 4508 1496 4516 1504
rect 4524 1496 4532 1504
rect 4556 1496 4564 1504
rect 4524 1476 4532 1484
rect 4540 1456 4548 1464
rect 4508 1436 4516 1444
rect 4540 1416 4548 1424
rect 4620 1636 4628 1644
rect 4620 1596 4628 1604
rect 4652 1716 4660 1724
rect 4716 1716 4724 1724
rect 4780 1716 4788 1724
rect 4812 1716 4820 1724
rect 4700 1696 4708 1704
rect 4668 1656 4676 1664
rect 4684 1656 4692 1664
rect 4684 1636 4692 1644
rect 4636 1576 4644 1584
rect 4636 1536 4644 1544
rect 4620 1516 4628 1524
rect 4828 1696 4836 1704
rect 4796 1676 4804 1684
rect 4844 1676 4852 1684
rect 4860 1676 4868 1684
rect 4892 1676 4900 1684
rect 4748 1656 4756 1664
rect 4764 1656 4772 1664
rect 5004 1856 5012 1864
rect 4972 1716 4980 1724
rect 4956 1696 4964 1704
rect 4940 1676 4948 1684
rect 4972 1676 4980 1684
rect 4908 1656 4916 1664
rect 4972 1656 4980 1664
rect 4812 1576 4820 1584
rect 4700 1516 4708 1524
rect 4716 1516 4724 1524
rect 4796 1516 4804 1524
rect 4956 1596 4964 1604
rect 4876 1556 4884 1564
rect 4876 1536 4884 1544
rect 4940 1536 4948 1544
rect 4876 1496 4884 1504
rect 4988 1536 4996 1544
rect 4860 1456 4868 1464
rect 4892 1456 4900 1464
rect 4908 1456 4916 1464
rect 4636 1416 4644 1424
rect 4780 1416 4788 1424
rect 4828 1416 4836 1424
rect 4892 1396 4900 1404
rect 4812 1356 4820 1364
rect 4700 1336 4708 1344
rect 4556 1316 4564 1324
rect 4492 1296 4500 1304
rect 4476 1276 4484 1284
rect 4540 1276 4548 1284
rect 4540 1256 4548 1264
rect 4428 1176 4436 1184
rect 4396 1116 4404 1124
rect 4476 1096 4484 1104
rect 4492 1076 4500 1084
rect 4460 1036 4468 1044
rect 4412 1016 4420 1024
rect 4460 996 4468 1004
rect 4380 956 4388 964
rect 4156 916 4164 924
rect 4220 916 4228 924
rect 4812 1296 4820 1304
rect 4700 1276 4708 1284
rect 4620 1236 4628 1244
rect 4556 1196 4564 1204
rect 4604 1136 4612 1144
rect 4572 1096 4580 1104
rect 4556 1076 4564 1084
rect 4588 1076 4596 1084
rect 4556 976 4564 984
rect 4524 956 4532 964
rect 4380 936 4388 944
rect 4412 936 4420 944
rect 4492 916 4500 924
rect 4492 896 4500 904
rect 4556 896 4564 904
rect 4396 876 4404 884
rect 4172 856 4180 864
rect 4300 856 4308 864
rect 4364 856 4372 864
rect 4428 856 4436 864
rect 4188 836 4196 844
rect 4332 836 4340 844
rect 4412 836 4420 844
rect 4364 816 4372 824
rect 4227 806 4235 814
rect 4237 806 4245 814
rect 4247 806 4255 814
rect 4257 806 4265 814
rect 4267 806 4275 814
rect 4277 806 4285 814
rect 4252 716 4260 724
rect 4188 556 4196 564
rect 4204 556 4212 564
rect 4252 536 4260 544
rect 4300 536 4308 544
rect 4172 516 4180 524
rect 4188 516 4196 524
rect 4156 476 4164 484
rect 4188 476 4196 484
rect 4300 476 4308 484
rect 4227 406 4235 414
rect 4237 406 4245 414
rect 4247 406 4255 414
rect 4257 406 4265 414
rect 4267 406 4275 414
rect 4277 406 4285 414
rect 4124 156 4132 164
rect 4444 836 4452 844
rect 4476 736 4484 744
rect 4508 736 4516 744
rect 4588 976 4596 984
rect 4588 936 4596 944
rect 4844 1136 4852 1144
rect 4876 1136 4884 1144
rect 4716 1116 4724 1124
rect 4732 1116 4740 1124
rect 4620 1096 4628 1104
rect 4636 1096 4644 1104
rect 4668 1096 4676 1104
rect 4764 1096 4772 1104
rect 4796 1096 4804 1104
rect 4828 1096 4836 1104
rect 4732 1076 4740 1084
rect 4716 1056 4724 1064
rect 4684 1016 4692 1024
rect 4668 996 4676 1004
rect 4652 956 4660 964
rect 4684 956 4692 964
rect 4652 936 4660 944
rect 4636 916 4644 924
rect 4460 696 4468 704
rect 4540 696 4548 704
rect 4604 696 4612 704
rect 4492 656 4500 664
rect 4476 636 4484 644
rect 4428 516 4436 524
rect 4364 496 4372 504
rect 4284 216 4292 224
rect 4332 156 4340 164
rect 4508 636 4516 644
rect 4668 776 4676 784
rect 4748 976 4756 984
rect 4780 976 4788 984
rect 4828 1076 4836 1084
rect 4860 1076 4868 1084
rect 4812 1056 4820 1064
rect 4796 936 4804 944
rect 4924 1156 4932 1164
rect 5020 1756 5028 1764
rect 5020 1736 5028 1744
rect 5084 1816 5092 1824
rect 5052 1736 5060 1744
rect 5068 1736 5076 1744
rect 5052 1716 5060 1724
rect 5036 1656 5044 1664
rect 5020 1636 5028 1644
rect 5004 1496 5012 1504
rect 4972 1456 4980 1464
rect 5036 1416 5044 1424
rect 4972 1296 4980 1304
rect 5004 1136 5012 1144
rect 4956 1116 4964 1124
rect 4972 1116 4980 1124
rect 4908 1096 4916 1104
rect 4924 1076 4932 1084
rect 4988 1076 4996 1084
rect 4892 1056 4900 1064
rect 4908 1056 4916 1064
rect 5004 1056 5012 1064
rect 4972 996 4980 1004
rect 5116 1816 5124 1824
rect 5148 1876 5156 1884
rect 5132 1736 5140 1744
rect 5100 1716 5108 1724
rect 5100 1656 5108 1664
rect 5084 1636 5092 1644
rect 5116 1616 5124 1624
rect 5180 1876 5188 1884
rect 5068 1536 5076 1544
rect 5116 1536 5124 1544
rect 5164 1536 5172 1544
rect 5084 1516 5092 1524
rect 5100 1516 5108 1524
rect 5164 1496 5172 1504
rect 5100 1476 5108 1484
rect 5116 1476 5124 1484
rect 5180 1476 5188 1484
rect 5148 1456 5156 1464
rect 5068 1316 5076 1324
rect 5132 1296 5140 1304
rect 5052 1256 5060 1264
rect 5052 1136 5060 1144
rect 5148 1196 5156 1204
rect 5132 1136 5140 1144
rect 5052 1116 5060 1124
rect 5212 1836 5220 1844
rect 5420 2136 5428 2144
rect 5404 2116 5412 2124
rect 5276 1816 5284 1824
rect 5388 1796 5396 1804
rect 5420 1836 5428 1844
rect 5228 1716 5236 1724
rect 5196 1296 5204 1304
rect 5148 1076 5156 1084
rect 5036 996 5044 1004
rect 5116 1056 5124 1064
rect 5020 976 5028 984
rect 5084 976 5092 984
rect 4988 956 4996 964
rect 4876 916 4884 924
rect 4732 896 4740 904
rect 4780 896 4788 904
rect 4716 736 4724 744
rect 4700 716 4708 724
rect 4844 776 4852 784
rect 4844 736 4852 744
rect 5116 916 5124 924
rect 5180 976 5188 984
rect 4988 756 4996 764
rect 5036 756 5044 764
rect 5068 756 5076 764
rect 5148 756 5156 764
rect 4908 716 4916 724
rect 4588 676 4596 684
rect 4652 676 4660 684
rect 4588 656 4596 664
rect 4556 636 4564 644
rect 4508 616 4516 624
rect 4540 616 4548 624
rect 4748 676 4756 684
rect 4684 616 4692 624
rect 4604 596 4612 604
rect 4668 596 4676 604
rect 4716 576 4724 584
rect 4620 556 4628 564
rect 4764 556 4772 564
rect 4492 516 4500 524
rect 4476 476 4484 484
rect 4764 536 4772 544
rect 4652 416 4660 424
rect 4492 256 4500 264
rect 4684 256 4692 264
rect 3964 116 3972 124
rect 3996 116 4004 124
rect 4716 236 4724 244
rect 4828 676 4836 684
rect 4796 636 4804 644
rect 4876 596 4884 604
rect 4908 696 4916 704
rect 4924 696 4932 704
rect 4972 696 4980 704
rect 5052 716 5060 724
rect 5020 676 5028 684
rect 5036 656 5044 664
rect 4940 576 4948 584
rect 4924 556 4932 564
rect 5004 576 5012 584
rect 4972 536 4980 544
rect 5020 536 5028 544
rect 4828 516 4836 524
rect 4844 516 4852 524
rect 4780 456 4788 464
rect 4764 336 4772 344
rect 4972 436 4980 444
rect 4828 376 4836 384
rect 4876 376 4884 384
rect 4796 336 4804 344
rect 4764 296 4772 304
rect 4828 256 4836 264
rect 5100 736 5108 744
rect 5084 716 5092 724
rect 5100 676 5108 684
rect 5164 676 5170 684
rect 5170 676 5172 684
rect 5068 576 5076 584
rect 5116 536 5124 544
rect 5084 516 5092 524
rect 5100 516 5108 524
rect 5148 556 5156 564
rect 5212 496 5220 504
rect 5196 376 5204 384
rect 5180 316 5188 324
rect 4988 256 4996 264
rect 4988 236 4996 244
rect 5020 236 5028 244
rect 5036 216 5044 224
rect 5180 276 5188 284
rect 5244 1456 5252 1464
rect 5308 1436 5316 1444
rect 5356 1416 5364 1424
rect 5340 1396 5348 1404
rect 5484 3436 5492 3444
rect 5468 2576 5476 2584
rect 5516 3076 5524 3084
rect 5516 2696 5524 2704
rect 5484 2436 5492 2444
rect 5516 2396 5524 2404
rect 5468 2256 5476 2264
rect 5468 1916 5476 1924
rect 5500 1896 5508 1904
rect 5452 1516 5460 1524
rect 5516 1496 5524 1504
rect 5420 1196 5428 1204
rect 5372 1056 5380 1064
rect 5372 996 5380 1004
rect 5340 956 5348 964
rect 5260 916 5268 924
rect 5420 816 5428 824
rect 5452 816 5460 824
rect 5356 656 5364 664
rect 5340 536 5348 544
rect 5340 516 5348 524
rect 5308 496 5316 504
rect 5468 496 5476 504
rect 5308 376 5316 384
rect 5276 336 5284 344
rect 5324 316 5332 324
rect 5244 296 5252 304
rect 5212 256 5220 264
rect 4588 116 4596 124
rect 4620 116 4628 124
rect 5452 116 5460 124
rect 5516 96 5524 104
rect 3260 36 3268 44
rect 3292 36 3300 44
rect 3708 36 3716 44
rect 5164 36 5172 44
rect 5356 36 5364 44
rect 3260 16 3268 24
rect 3516 16 3524 24
rect 4227 6 4235 14
rect 4237 6 4245 14
rect 4247 6 4255 14
rect 4257 6 4265 14
rect 4267 6 4275 14
rect 4277 6 4285 14
rect 4700 16 4708 24
<< metal3 >>
rect 2068 3817 2092 3823
rect 3412 3817 3484 3823
rect 2722 3814 2782 3816
rect 2722 3806 2723 3814
rect 2732 3806 2733 3814
rect 2771 3806 2772 3814
rect 2781 3806 2782 3814
rect 2722 3804 2782 3806
rect 3444 3797 3500 3803
rect 1972 3777 2188 3783
rect 3284 3777 3884 3783
rect 196 3757 524 3763
rect 532 3757 892 3763
rect 1348 3757 2492 3763
rect 2740 3757 3020 3763
rect 3156 3757 3308 3763
rect 3364 3757 3420 3763
rect 4116 3757 4540 3763
rect 4884 3757 5292 3763
rect 228 3737 268 3743
rect 932 3737 2364 3743
rect 2436 3737 2476 3743
rect 2964 3737 3004 3743
rect 3204 3737 3372 3743
rect 3412 3737 3468 3743
rect 3604 3737 3612 3743
rect 3876 3737 3932 3743
rect 3940 3737 4268 3743
rect 4468 3737 4844 3743
rect 5028 3737 5068 3743
rect 5092 3737 5324 3743
rect 324 3717 380 3723
rect 1620 3717 1756 3723
rect 2292 3717 2348 3723
rect 2356 3717 2460 3723
rect 2468 3717 2988 3723
rect 3108 3717 3148 3723
rect 3188 3717 3228 3723
rect 3380 3717 3452 3723
rect 3460 3717 3820 3723
rect 3924 3717 4380 3723
rect 4644 3717 4748 3723
rect 4964 3717 5212 3723
rect 5300 3717 5324 3723
rect 1732 3697 1868 3703
rect 2164 3697 2220 3703
rect 2276 3697 2332 3703
rect 2340 3697 2444 3703
rect 2452 3697 2972 3703
rect 2980 3697 3276 3703
rect 3300 3697 3340 3703
rect 5060 3697 5100 3703
rect 740 3677 2300 3683
rect 2340 3677 2364 3683
rect 2516 3677 3132 3683
rect 3197 3677 3324 3683
rect 932 3657 1148 3663
rect 1156 3657 2396 3663
rect 2420 3657 2524 3663
rect 2564 3657 3052 3663
rect 3060 3657 3084 3663
rect 3197 3663 3203 3677
rect 3668 3677 3884 3683
rect 3908 3677 4076 3683
rect 5076 3677 5260 3683
rect 3124 3657 3203 3663
rect 3220 3657 3516 3663
rect 3524 3657 3996 3663
rect 692 3637 716 3643
rect 2196 3637 2460 3643
rect 2548 3637 2924 3643
rect 3252 3637 3644 3643
rect 3652 3637 4108 3643
rect 1940 3617 1996 3623
rect 2996 3617 3068 3623
rect 3076 3617 3612 3623
rect 3700 3617 3900 3623
rect 3924 3617 3948 3623
rect 3965 3617 4124 3623
rect 1218 3614 1278 3616
rect 1218 3606 1219 3614
rect 1228 3606 1229 3614
rect 1267 3606 1268 3614
rect 1277 3606 1278 3614
rect 1218 3604 1278 3606
rect 3028 3597 3884 3603
rect 3965 3603 3971 3617
rect 4226 3614 4286 3616
rect 4226 3606 4227 3614
rect 4236 3606 4237 3614
rect 4275 3606 4276 3614
rect 4285 3606 4286 3614
rect 4226 3604 4286 3606
rect 3940 3597 3971 3603
rect 3988 3597 4060 3603
rect 4884 3597 5036 3603
rect 388 3577 444 3583
rect 452 3577 492 3583
rect 500 3577 732 3583
rect 980 3577 2540 3583
rect 3252 3577 3468 3583
rect 3476 3577 3724 3583
rect 3828 3577 3964 3583
rect 3988 3577 4412 3583
rect 4436 3577 4796 3583
rect 2500 3557 2540 3563
rect 2548 3557 3036 3563
rect 3108 3557 3788 3563
rect 3876 3557 4092 3563
rect 4109 3557 4732 3563
rect 2820 3537 3116 3543
rect 3124 3537 3212 3543
rect 3236 3537 3388 3543
rect 3764 3537 3788 3543
rect 3844 3537 3996 3543
rect 4020 3537 4060 3543
rect 4109 3543 4115 3557
rect 4772 3557 4988 3563
rect 4084 3537 4115 3543
rect 4132 3537 4428 3543
rect 4452 3537 4492 3543
rect 4548 3537 4748 3543
rect 4836 3537 4924 3543
rect 4948 3537 5004 3543
rect 5012 3537 5228 3543
rect 436 3517 476 3523
rect 484 3517 540 3523
rect 548 3517 2156 3523
rect 2516 3517 2556 3523
rect 2676 3517 2700 3523
rect 3044 3517 3148 3523
rect 3220 3517 3372 3523
rect 3380 3517 3964 3523
rect 3972 3517 4028 3523
rect 4084 3517 4204 3523
rect 4356 3517 4396 3523
rect 4404 3517 4508 3523
rect 4516 3517 4620 3523
rect 4660 3517 5084 3523
rect 836 3497 1004 3503
rect 1236 3497 1404 3503
rect 1412 3497 1436 3503
rect 2068 3497 2092 3503
rect 2100 3497 2204 3503
rect 2436 3497 2684 3503
rect 2980 3497 3068 3503
rect 3108 3497 3148 3503
rect 3156 3497 3212 3503
rect 3380 3497 3420 3503
rect 3476 3497 3532 3503
rect 3748 3497 4044 3503
rect 4068 3497 4108 3503
rect 4132 3497 4220 3503
rect 4372 3497 4428 3503
rect 4596 3497 4620 3503
rect 4660 3497 4780 3503
rect 4804 3497 4844 3503
rect 4932 3497 4972 3503
rect 4996 3497 5132 3503
rect 228 3477 444 3483
rect 1124 3477 1708 3483
rect 2580 3477 3228 3483
rect 3245 3477 3388 3483
rect 1940 3457 2284 3463
rect 2788 3457 2860 3463
rect 3245 3463 3251 3477
rect 3396 3477 3452 3483
rect 3524 3477 4108 3483
rect 4116 3477 4524 3483
rect 4532 3477 4668 3483
rect 4676 3477 4716 3483
rect 4724 3477 4876 3483
rect 3188 3457 3251 3463
rect 3348 3457 3404 3463
rect 3412 3457 3644 3463
rect 3652 3457 3852 3463
rect 3860 3457 4204 3463
rect 4093 3444 4099 3457
rect 4436 3457 4540 3463
rect 4660 3457 4684 3463
rect 4740 3457 4796 3463
rect 36 3437 396 3443
rect 756 3437 892 3443
rect 2324 3437 2380 3443
rect 2660 3437 2812 3443
rect 2820 3437 2908 3443
rect 3076 3437 3260 3443
rect 3300 3437 3516 3443
rect 3524 3437 3660 3443
rect 3684 3437 3708 3443
rect 3716 3437 3948 3443
rect 3972 3437 4012 3443
rect 4612 3437 4860 3443
rect 4884 3437 5020 3443
rect 5076 3437 5228 3443
rect 5396 3437 5484 3443
rect 516 3417 684 3423
rect 1124 3417 1148 3423
rect 1156 3417 1292 3423
rect 1300 3417 1516 3423
rect 1524 3417 1564 3423
rect 1572 3417 1644 3423
rect 1652 3417 1932 3423
rect 1972 3417 1996 3423
rect 3460 3417 3644 3423
rect 3661 3423 3667 3436
rect 3661 3417 4556 3423
rect 4580 3417 4732 3423
rect 5172 3417 5244 3423
rect 2722 3414 2782 3416
rect 2722 3406 2723 3414
rect 2732 3406 2733 3414
rect 2771 3406 2772 3414
rect 2781 3406 2782 3414
rect 2722 3404 2782 3406
rect 196 3397 220 3403
rect 532 3397 812 3403
rect 1780 3397 1916 3403
rect 3284 3397 3372 3403
rect 3428 3397 3548 3403
rect 3572 3397 3660 3403
rect 3668 3397 4476 3403
rect 4692 3397 4700 3403
rect 580 3377 732 3383
rect 740 3377 956 3383
rect 1533 3383 1539 3396
rect 1533 3377 1948 3383
rect 2916 3377 3084 3383
rect 3092 3377 3244 3383
rect 3252 3377 3260 3383
rect 3428 3377 3484 3383
rect 3636 3377 3820 3383
rect 4004 3377 4124 3383
rect 4132 3377 4364 3383
rect 4596 3377 5036 3383
rect 5076 3377 5148 3383
rect 5236 3377 5372 3383
rect 500 3357 748 3363
rect 2292 3357 2364 3363
rect 2484 3357 3564 3363
rect 3652 3357 3740 3363
rect 3764 3357 3916 3363
rect 3988 3357 4172 3363
rect 4228 3357 4444 3363
rect 4452 3357 4652 3363
rect 4660 3357 4748 3363
rect 5044 3357 5164 3363
rect 5220 3357 5436 3363
rect 468 3337 524 3343
rect 804 3337 892 3343
rect 900 3337 972 3343
rect 1604 3337 1692 3343
rect 1876 3337 1932 3343
rect 1940 3337 2012 3343
rect 2404 3337 2556 3343
rect 3540 3337 4012 3343
rect 4221 3343 4227 3356
rect 4020 3337 4227 3343
rect 4372 3337 4716 3343
rect 5092 3337 5164 3343
rect 5172 3337 5356 3343
rect 420 3317 572 3323
rect 644 3317 668 3323
rect 836 3317 876 3323
rect 884 3317 908 3323
rect 1748 3317 2060 3323
rect 2068 3317 2092 3323
rect 2212 3317 2284 3323
rect 3108 3317 3372 3323
rect 3380 3317 3436 3323
rect 3556 3317 3628 3323
rect 3636 3317 3756 3323
rect 3828 3317 4348 3323
rect 4484 3317 4492 3323
rect 4500 3317 4556 3323
rect 4980 3317 5100 3323
rect 5252 3317 5308 3323
rect 260 3297 444 3303
rect 516 3297 588 3303
rect 708 3297 748 3303
rect 756 3297 860 3303
rect 868 3297 1036 3303
rect 1156 3297 1404 3303
rect 1764 3297 1804 3303
rect 1892 3297 2044 3303
rect 2052 3297 2124 3303
rect 3524 3297 3580 3303
rect 3588 3297 3596 3303
rect 3604 3297 3724 3303
rect 3732 3297 3836 3303
rect 3844 3297 3884 3303
rect 3892 3297 3948 3303
rect 3956 3297 4076 3303
rect 4100 3297 4364 3303
rect 4420 3297 4460 3303
rect 4868 3297 4940 3303
rect 5028 3297 5212 3303
rect 5348 3297 5372 3303
rect 5460 3297 5555 3303
rect 436 3277 652 3283
rect 948 3277 1116 3283
rect 3620 3277 3756 3283
rect 3988 3277 3996 3283
rect 4052 3277 4076 3283
rect 4084 3277 4524 3283
rect 5044 3277 5068 3283
rect 5140 3277 5404 3283
rect 484 3257 524 3263
rect 532 3257 924 3263
rect 3076 3257 3564 3263
rect 3572 3257 3788 3263
rect 3805 3257 4012 3263
rect 2868 3237 3692 3243
rect 3805 3243 3811 3257
rect 4052 3257 4284 3263
rect 3716 3237 3811 3243
rect 3940 3237 4124 3243
rect 4205 3237 4380 3243
rect 276 3217 300 3223
rect 724 3217 1068 3223
rect 1524 3217 1564 3223
rect 1828 3217 2060 3223
rect 2068 3217 2124 3223
rect 2388 3217 2444 3223
rect 3156 3217 3180 3223
rect 3540 3217 3644 3223
rect 3668 3217 3692 3223
rect 3764 3217 3916 3223
rect 4205 3223 4211 3237
rect 4084 3217 4211 3223
rect 4420 3217 4780 3223
rect 4788 3217 4988 3223
rect 1218 3214 1278 3216
rect 1218 3206 1219 3214
rect 1228 3206 1229 3214
rect 1267 3206 1268 3214
rect 1277 3206 1278 3214
rect 1218 3204 1278 3206
rect 4226 3214 4286 3216
rect 4226 3206 4227 3214
rect 4236 3206 4237 3214
rect 4275 3206 4276 3214
rect 4285 3206 4286 3214
rect 4226 3204 4286 3206
rect 1604 3197 1676 3203
rect 2109 3197 2332 3203
rect 2109 3184 2115 3197
rect 3076 3197 3324 3203
rect 3764 3197 4028 3203
rect 4036 3197 4092 3203
rect 4852 3197 4988 3203
rect 4996 3197 5116 3203
rect 36 3177 172 3183
rect 180 3177 252 3183
rect 260 3177 316 3183
rect 1492 3177 1676 3183
rect 1732 3177 1820 3183
rect 1924 3177 2108 3183
rect 2148 3177 2268 3183
rect 2276 3177 2380 3183
rect 2884 3177 3308 3183
rect 3476 3177 4428 3183
rect 4740 3177 4748 3183
rect 484 3157 524 3163
rect 548 3157 556 3163
rect 564 3157 604 3163
rect 2004 3157 2300 3163
rect 2372 3157 2668 3163
rect 3709 3157 4348 3163
rect 3709 3144 3715 3157
rect 100 3137 124 3143
rect 244 3137 380 3143
rect 420 3137 572 3143
rect 740 3137 1052 3143
rect 1412 3137 1756 3143
rect 2100 3137 2188 3143
rect 3268 3137 3356 3143
rect 3380 3137 3484 3143
rect 3492 3137 3708 3143
rect 3876 3137 3980 3143
rect 3988 3137 4012 3143
rect 4020 3137 4060 3143
rect 20 3117 60 3123
rect 125 3123 131 3136
rect 125 3117 428 3123
rect 452 3117 668 3123
rect 964 3117 1084 3123
rect 1108 3117 1292 3123
rect 1300 3117 1372 3123
rect 1732 3117 1772 3123
rect 1828 3117 2012 3123
rect 2020 3117 2156 3123
rect 2164 3117 2172 3123
rect 2205 3117 2284 3123
rect 84 3097 188 3103
rect 196 3097 236 3103
rect 244 3097 556 3103
rect 596 3097 620 3103
rect 660 3097 988 3103
rect 1156 3097 1212 3103
rect 1220 3097 1356 3103
rect 1652 3097 1692 3103
rect 1812 3097 1948 3103
rect 2036 3097 2140 3103
rect 2205 3103 2211 3117
rect 3236 3117 3484 3123
rect 3620 3117 3836 3123
rect 3949 3117 4076 3123
rect 3949 3104 3955 3117
rect 4308 3117 4364 3123
rect 5348 3117 5372 3123
rect 5428 3117 5555 3123
rect 2148 3097 2211 3103
rect 2228 3097 2364 3103
rect 2372 3097 2492 3103
rect 2548 3097 3228 3103
rect 3364 3097 3468 3103
rect 3492 3097 3596 3103
rect 3764 3097 3788 3103
rect 4004 3097 4332 3103
rect 4964 3097 5100 3103
rect 5124 3097 5308 3103
rect 308 3077 444 3083
rect 500 3077 732 3083
rect 788 3077 1452 3083
rect 2541 3083 2547 3096
rect 1460 3077 2547 3083
rect 3316 3077 3404 3083
rect 3412 3077 3468 3083
rect 3540 3077 3692 3083
rect 3700 3077 3820 3083
rect 3860 3077 3900 3083
rect 4052 3077 4060 3083
rect 4084 3077 4124 3083
rect 4404 3077 4540 3083
rect 5092 3077 5132 3083
rect 5140 3077 5212 3083
rect 5220 3077 5260 3083
rect 5300 3077 5356 3083
rect 5524 3077 5555 3083
rect 52 3057 140 3063
rect 148 3057 220 3063
rect 340 3057 348 3063
rect 356 3057 508 3063
rect 676 3057 764 3063
rect 772 3057 796 3063
rect 884 3057 924 3063
rect 1124 3057 1228 3063
rect 1364 3057 1612 3063
rect 1764 3057 1772 3063
rect 1780 3057 1804 3063
rect 1924 3057 2204 3063
rect 2388 3057 2476 3063
rect 3412 3057 3516 3063
rect 3652 3057 3756 3063
rect 3780 3057 3996 3063
rect 4308 3057 4444 3063
rect 4580 3057 4684 3063
rect 4692 3057 4748 3063
rect 4948 3057 4972 3063
rect 4980 3057 5036 3063
rect 116 3037 332 3043
rect 468 3037 540 3043
rect 660 3037 684 3043
rect 724 3037 748 3043
rect 1316 3037 1427 3043
rect 404 3017 620 3023
rect 676 3017 716 3023
rect 1421 3023 1427 3037
rect 1572 3037 2508 3043
rect 2516 3037 2588 3043
rect 3476 3037 3612 3043
rect 3636 3037 3660 3043
rect 3668 3037 3724 3043
rect 4324 3037 4396 3043
rect 4916 3037 5036 3043
rect 5044 3037 5068 3043
rect 5076 3037 5372 3043
rect 1421 3017 1692 3023
rect 1700 3017 1788 3023
rect 1796 3017 1852 3023
rect 2004 3017 2028 3023
rect 3060 3017 3180 3023
rect 3236 3017 4924 3023
rect 4932 3017 4940 3023
rect 5060 3017 5116 3023
rect 2722 3014 2782 3016
rect 2722 3006 2723 3014
rect 2732 3006 2733 3014
rect 2771 3006 2772 3014
rect 2781 3006 2782 3014
rect 2722 3004 2782 3006
rect 436 2997 492 3003
rect 532 2997 572 3003
rect 1204 2997 1324 3003
rect 1332 2997 1340 3003
rect 1812 2997 2012 3003
rect 3444 2997 3900 3003
rect 3908 2997 4092 3003
rect 4612 2997 4652 3003
rect 5012 2997 5244 3003
rect 5252 2997 5324 3003
rect 196 2977 332 2983
rect 1092 2977 1196 2983
rect 1636 2977 2428 2983
rect 2468 2977 2924 2983
rect 2932 2977 3308 2983
rect 3316 2977 3340 2983
rect 3460 2977 3468 2983
rect 3604 2977 3740 2983
rect 3796 2977 3836 2983
rect 3844 2977 3964 2983
rect 3988 2977 4380 2983
rect 4948 2977 5020 2983
rect 5028 2977 5100 2983
rect 132 2957 140 2963
rect 148 2957 188 2963
rect 212 2957 364 2963
rect 372 2957 412 2963
rect 564 2957 748 2963
rect 756 2957 908 2963
rect 1988 2957 2124 2963
rect 2196 2957 2348 2963
rect 2676 2957 2924 2963
rect 2964 2957 3660 2963
rect 3700 2957 3852 2963
rect 3965 2963 3971 2976
rect 3965 2957 4156 2963
rect 4493 2957 4924 2963
rect 4493 2944 4499 2957
rect 4996 2957 5180 2963
rect 5188 2957 5356 2963
rect 340 2937 700 2943
rect 1540 2937 1580 2943
rect 1588 2937 1596 2943
rect 1604 2937 1644 2943
rect 1876 2937 1916 2943
rect 1924 2937 1980 2943
rect 2052 2937 2236 2943
rect 2244 2937 2316 2943
rect 2324 2937 2396 2943
rect 3124 2937 3372 2943
rect 3476 2937 3532 2943
rect 3684 2937 3772 2943
rect 3956 2937 3996 2943
rect 4372 2937 4492 2943
rect 4788 2937 4892 2943
rect 5044 2937 5164 2943
rect 116 2917 220 2923
rect 228 2917 380 2923
rect 692 2917 828 2923
rect 1172 2917 1260 2923
rect 1380 2917 1420 2923
rect 1508 2917 1548 2923
rect 1924 2917 1964 2923
rect 2036 2917 2204 2923
rect 2212 2917 2284 2923
rect 2292 2917 2364 2923
rect 2500 2917 2636 2923
rect 3220 2917 3228 2923
rect 3284 2917 3372 2923
rect 3380 2917 3747 2923
rect 36 2897 60 2903
rect 68 2897 140 2903
rect 1236 2897 1324 2903
rect 1748 2897 1900 2903
rect 2020 2897 2076 2903
rect 2084 2897 2140 2903
rect 2340 2897 2348 2903
rect 2484 2897 2668 2903
rect 3364 2897 3404 2903
rect 3412 2897 3452 2903
rect 3741 2903 3747 2917
rect 3764 2917 3836 2923
rect 3860 2917 3964 2923
rect 4148 2917 4188 2923
rect 4228 2917 4316 2923
rect 4340 2917 4428 2923
rect 4724 2917 4956 2923
rect 4996 2917 5004 2923
rect 5204 2917 5228 2923
rect 3741 2897 3756 2903
rect 3764 2897 3772 2903
rect 3780 2897 3884 2903
rect 4004 2897 4012 2903
rect 196 2877 252 2883
rect 260 2877 348 2883
rect 1300 2877 1484 2883
rect 1700 2877 1820 2883
rect 2324 2877 2444 2883
rect 3300 2877 3564 2883
rect 3572 2877 3724 2883
rect 3732 2877 3820 2883
rect 3828 2877 3916 2883
rect 3924 2877 4028 2883
rect 404 2857 444 2863
rect 3293 2863 3299 2876
rect 1108 2857 3299 2863
rect 3444 2857 3500 2863
rect 3812 2857 3884 2863
rect 3892 2857 3932 2863
rect 4292 2857 4540 2863
rect 756 2837 1020 2843
rect 1092 2837 1340 2843
rect 1364 2837 1628 2843
rect 1732 2837 1932 2843
rect 2068 2837 2764 2843
rect 4468 2837 4524 2843
rect 196 2817 556 2823
rect 1684 2817 1788 2823
rect 1796 2817 2540 2823
rect 5284 2817 5308 2823
rect 1218 2814 1278 2816
rect 1218 2806 1219 2814
rect 1228 2806 1229 2814
rect 1267 2806 1268 2814
rect 1277 2806 1278 2814
rect 1218 2804 1278 2806
rect 4226 2814 4286 2816
rect 4226 2806 4227 2814
rect 4236 2806 4237 2814
rect 4275 2806 4276 2814
rect 4285 2806 4286 2814
rect 4226 2804 4286 2806
rect 1716 2797 1852 2803
rect 2820 2797 2828 2803
rect 2836 2797 2956 2803
rect 2964 2797 3068 2803
rect 5268 2797 5308 2803
rect 1588 2777 1740 2783
rect 1892 2777 2076 2783
rect 4900 2777 4972 2783
rect 308 2757 476 2763
rect 1460 2757 1740 2763
rect 2068 2757 2156 2763
rect 2964 2757 3548 2763
rect 3556 2757 4220 2763
rect 228 2737 380 2743
rect 1508 2737 1612 2743
rect 1684 2737 1724 2743
rect 1764 2737 1868 2743
rect 1908 2737 1932 2743
rect 2004 2737 2108 2743
rect 2356 2737 2380 2743
rect 2436 2737 2476 2743
rect 2484 2737 3356 2743
rect 3364 2737 3532 2743
rect 292 2717 300 2723
rect 372 2717 476 2723
rect 612 2717 652 2723
rect 660 2717 700 2723
rect 1156 2717 1452 2723
rect 1460 2717 1804 2723
rect 1812 2717 2028 2723
rect 2100 2717 2252 2723
rect 2532 2717 2556 2723
rect 3396 2717 3468 2723
rect 4084 2717 4860 2723
rect 388 2697 396 2703
rect 532 2697 556 2703
rect 644 2697 732 2703
rect 1364 2697 1388 2703
rect 1572 2697 1660 2703
rect 1780 2697 1820 2703
rect 1892 2697 1932 2703
rect 1956 2697 1980 2703
rect 1988 2697 2028 2703
rect 2276 2697 2364 2703
rect 2516 2697 2540 2703
rect 3332 2697 3436 2703
rect 3556 2697 3868 2703
rect 4100 2697 4188 2703
rect 4356 2697 4412 2703
rect 4436 2697 4732 2703
rect 4836 2697 4972 2703
rect 5524 2697 5555 2703
rect 388 2677 492 2683
rect 548 2677 604 2683
rect 692 2677 748 2683
rect 756 2677 860 2683
rect 1236 2677 1324 2683
rect 1332 2677 1484 2683
rect 1524 2677 1548 2683
rect 1636 2677 1756 2683
rect 1780 2677 2316 2683
rect 2452 2677 2700 2683
rect 3972 2677 4364 2683
rect 4404 2677 4492 2683
rect 4500 2677 4796 2683
rect 5092 2677 5148 2683
rect 372 2657 444 2663
rect 452 2657 460 2663
rect 692 2657 716 2663
rect 756 2657 876 2663
rect 1348 2657 1788 2663
rect 1940 2657 2060 2663
rect 2068 2657 2108 2663
rect 2148 2657 2204 2663
rect 2212 2657 2268 2663
rect 2436 2657 2476 2663
rect 2500 2657 2588 2663
rect 2612 2657 2892 2663
rect 2900 2657 3020 2663
rect 3092 2657 3196 2663
rect 3204 2657 3644 2663
rect 3652 2657 3996 2663
rect 4180 2657 4300 2663
rect 4516 2657 4700 2663
rect 4708 2657 4812 2663
rect 4916 2657 5244 2663
rect 532 2637 572 2643
rect 1044 2637 1404 2643
rect 1428 2637 1516 2643
rect 1748 2637 1788 2643
rect 1892 2637 2556 2643
rect 4820 2637 4908 2643
rect 4964 2637 5052 2643
rect 5060 2637 5276 2643
rect 420 2617 620 2623
rect 1380 2617 1404 2623
rect 1460 2617 1676 2623
rect 1684 2617 2460 2623
rect 3060 2617 3180 2623
rect 3284 2617 3404 2623
rect 3492 2617 3612 2623
rect 4452 2617 4652 2623
rect 4676 2617 4684 2623
rect 2722 2614 2782 2616
rect 2722 2606 2723 2614
rect 2732 2606 2733 2614
rect 2771 2606 2772 2614
rect 2781 2606 2782 2614
rect 2722 2604 2782 2606
rect 916 2597 972 2603
rect 980 2597 1068 2603
rect 1076 2597 1196 2603
rect 1668 2597 1676 2603
rect 1748 2597 2524 2603
rect 2868 2597 3052 2603
rect 3060 2597 3100 2603
rect 3172 2597 3228 2603
rect 3380 2597 3420 2603
rect 3428 2597 3756 2603
rect 4468 2597 4476 2603
rect 436 2577 732 2583
rect 1780 2577 1932 2583
rect 2020 2577 2076 2583
rect 2084 2577 2140 2583
rect 2420 2577 3404 2583
rect 3412 2577 3804 2583
rect 3812 2577 3820 2583
rect 4340 2577 4556 2583
rect 4564 2577 4732 2583
rect 4820 2577 5420 2583
rect 5428 2577 5468 2583
rect 20 2557 92 2563
rect 100 2557 140 2563
rect 324 2557 332 2563
rect 420 2557 444 2563
rect 644 2557 764 2563
rect 772 2557 812 2563
rect 1332 2557 1436 2563
rect 1444 2557 1580 2563
rect 1860 2557 1948 2563
rect 2068 2557 2092 2563
rect 2244 2557 2636 2563
rect 2644 2557 2860 2563
rect 2900 2557 3212 2563
rect 3476 2557 3628 2563
rect 3668 2557 3948 2563
rect 3956 2557 4060 2563
rect 4068 2557 4508 2563
rect 4948 2557 5148 2563
rect 77 2537 204 2543
rect 77 2524 83 2537
rect 260 2537 364 2543
rect 436 2537 540 2543
rect 708 2537 748 2543
rect 1620 2537 2236 2543
rect 2276 2537 2348 2543
rect 3236 2537 3292 2543
rect 3348 2537 3388 2543
rect 4308 2537 4316 2543
rect 4324 2537 4348 2543
rect 4772 2537 4924 2543
rect 52 2517 76 2523
rect 132 2517 140 2523
rect 148 2517 156 2523
rect 244 2517 268 2523
rect 276 2517 316 2523
rect 356 2517 492 2523
rect 644 2517 668 2523
rect 708 2517 1004 2523
rect 1220 2517 1692 2523
rect 3300 2517 3452 2523
rect 4196 2517 4428 2523
rect 4724 2517 5100 2523
rect 5108 2517 5116 2523
rect 516 2497 524 2503
rect 596 2497 620 2503
rect 628 2497 684 2503
rect 1236 2497 1500 2503
rect 2772 2497 2828 2503
rect 3188 2497 3548 2503
rect 4228 2497 4684 2503
rect 4708 2497 4748 2503
rect 116 2477 380 2483
rect 468 2477 652 2483
rect 1108 2477 1148 2483
rect 1156 2477 1340 2483
rect 1348 2477 1404 2483
rect 1412 2477 1580 2483
rect 1588 2477 1820 2483
rect 3460 2477 3468 2483
rect 3668 2477 4428 2483
rect 196 2457 204 2463
rect 308 2457 396 2463
rect 420 2457 476 2463
rect 580 2457 588 2463
rect 596 2457 620 2463
rect 628 2457 764 2463
rect 1364 2457 1468 2463
rect 3188 2457 3212 2463
rect 4324 2457 4508 2463
rect 4196 2437 4780 2443
rect 4788 2437 4828 2443
rect 4836 2437 5164 2443
rect 5172 2437 5308 2443
rect 5444 2437 5484 2443
rect 468 2417 492 2423
rect 1524 2417 1548 2423
rect 2132 2417 2412 2423
rect 2580 2417 2636 2423
rect 2676 2417 3564 2423
rect 4340 2417 4412 2423
rect 1218 2414 1278 2416
rect 1218 2406 1219 2414
rect 1228 2406 1229 2414
rect 1267 2406 1268 2414
rect 1277 2406 1278 2414
rect 1218 2404 1278 2406
rect 4226 2414 4286 2416
rect 4226 2406 4227 2414
rect 4236 2406 4237 2414
rect 4275 2406 4276 2414
rect 4285 2406 4286 2414
rect 4226 2404 4286 2406
rect 500 2397 732 2403
rect 740 2397 1036 2403
rect 1716 2397 1852 2403
rect 1860 2397 2092 2403
rect 2100 2397 3075 2403
rect 404 2377 700 2383
rect 708 2377 748 2383
rect 1028 2377 2060 2383
rect 3028 2377 3052 2383
rect 3069 2383 3075 2397
rect 3092 2397 3596 2403
rect 4388 2397 4412 2403
rect 5524 2397 5555 2403
rect 3069 2377 3644 2383
rect 3652 2377 3660 2383
rect 4212 2377 4444 2383
rect 4564 2377 4588 2383
rect 388 2357 508 2363
rect 532 2357 1004 2363
rect 1844 2357 3308 2363
rect 3316 2357 3516 2363
rect 3620 2357 3660 2363
rect 4301 2357 4860 2363
rect 388 2337 604 2343
rect 612 2337 684 2343
rect 692 2337 732 2343
rect 788 2337 844 2343
rect 852 2337 876 2343
rect 1508 2337 1612 2343
rect 1780 2337 1804 2343
rect 1812 2337 1884 2343
rect 1892 2337 1948 2343
rect 1956 2337 2492 2343
rect 4301 2343 4307 2357
rect 4868 2357 5516 2363
rect 3364 2337 4307 2343
rect 4324 2337 4396 2343
rect 4404 2337 4604 2343
rect 4612 2337 4668 2343
rect 5549 2343 5555 2363
rect 4948 2337 5555 2343
rect 228 2317 444 2323
rect 724 2317 828 2323
rect 1460 2317 1532 2323
rect 1588 2317 1628 2323
rect 1668 2317 1676 2323
rect 1684 2317 1708 2323
rect 1780 2317 1788 2323
rect 1796 2317 1916 2323
rect 2036 2317 2092 2323
rect 2772 2317 3116 2323
rect 3316 2317 3372 2323
rect 3604 2317 3676 2323
rect 3716 2317 4156 2323
rect 4164 2317 4188 2323
rect 4292 2317 4412 2323
rect 4420 2317 4460 2323
rect 4468 2317 4572 2323
rect 4580 2317 4636 2323
rect 4660 2317 4764 2323
rect 4788 2317 4876 2323
rect 5364 2317 5404 2323
rect 5412 2317 5555 2323
rect 52 2297 364 2303
rect 468 2297 476 2303
rect 612 2297 652 2303
rect 804 2297 860 2303
rect 868 2297 924 2303
rect 932 2297 1052 2303
rect 1604 2297 1692 2303
rect 1924 2297 1996 2303
rect 2356 2297 2492 2303
rect 2708 2297 2764 2303
rect 3220 2297 3276 2303
rect 3284 2297 3324 2303
rect 3332 2297 3388 2303
rect 3396 2297 3564 2303
rect 3572 2297 3660 2303
rect 3780 2297 4291 2303
rect 196 2277 227 2283
rect 221 2264 227 2277
rect 404 2277 508 2283
rect 628 2277 1020 2283
rect 1332 2277 1388 2283
rect 1396 2277 1580 2283
rect 1588 2277 1660 2283
rect 1668 2277 1740 2283
rect 1748 2277 1980 2283
rect 1988 2277 2124 2283
rect 2836 2277 3196 2283
rect 3204 2277 3228 2283
rect 3252 2277 3324 2283
rect 3348 2277 3372 2283
rect 3380 2277 3436 2283
rect 3540 2277 3708 2283
rect 3988 2277 4188 2283
rect 4285 2283 4291 2297
rect 4308 2297 4364 2303
rect 4564 2297 4796 2303
rect 4852 2297 5164 2303
rect 4285 2277 4316 2283
rect 4324 2277 4348 2283
rect 4516 2277 4579 2283
rect 196 2257 204 2263
rect 397 2263 403 2276
rect 4573 2264 4579 2277
rect 4612 2277 4700 2283
rect 4724 2277 4732 2283
rect 4756 2277 4972 2283
rect 5524 2277 5555 2283
rect 340 2257 403 2263
rect 548 2257 620 2263
rect 1460 2257 1788 2263
rect 2052 2257 2252 2263
rect 2452 2257 2764 2263
rect 3060 2257 3292 2263
rect 3428 2257 3500 2263
rect 3508 2257 3724 2263
rect 3796 2257 4124 2263
rect 4180 2257 4332 2263
rect 4436 2257 4508 2263
rect 4580 2257 4796 2263
rect 4964 2257 5132 2263
rect 5236 2257 5260 2263
rect 5380 2257 5420 2263
rect 5428 2257 5468 2263
rect 308 2237 796 2243
rect 868 2237 972 2243
rect 1140 2237 1244 2243
rect 1652 2237 1692 2243
rect 1700 2237 1724 2243
rect 1764 2237 1868 2243
rect 3748 2237 3788 2243
rect 3860 2237 4108 2243
rect 4132 2237 4236 2243
rect 4244 2237 4380 2243
rect 4388 2237 4700 2243
rect 4708 2237 4732 2243
rect 4740 2237 4748 2243
rect 4756 2237 5372 2243
rect 68 2217 428 2223
rect 1604 2217 1628 2223
rect 1636 2217 1788 2223
rect 1796 2217 1852 2223
rect 1972 2217 2204 2223
rect 2852 2217 3020 2223
rect 3028 2217 3084 2223
rect 3092 2217 3196 2223
rect 3236 2217 3900 2223
rect 4036 2217 4140 2223
rect 4340 2217 4524 2223
rect 4596 2217 4908 2223
rect 5092 2217 5228 2223
rect 2722 2214 2782 2216
rect 2722 2206 2723 2214
rect 2732 2206 2733 2214
rect 2771 2206 2772 2214
rect 2781 2206 2782 2214
rect 2722 2204 2782 2206
rect 228 2197 284 2203
rect 292 2197 316 2203
rect 324 2197 556 2203
rect 1476 2197 1676 2203
rect 1684 2197 1996 2203
rect 2276 2197 2380 2203
rect 2580 2197 2636 2203
rect 2900 2197 3260 2203
rect 3268 2197 3372 2203
rect 3396 2197 3692 2203
rect 3700 2197 4940 2203
rect 4957 2197 5324 2203
rect 164 2177 652 2183
rect 660 2177 684 2183
rect 788 2177 956 2183
rect 1364 2177 2508 2183
rect 2564 2177 3420 2183
rect 3444 2177 3548 2183
rect 3556 2177 3708 2183
rect 3764 2177 3884 2183
rect 4004 2177 4124 2183
rect 4356 2177 4492 2183
rect 4957 2183 4963 2197
rect 4500 2177 4963 2183
rect 5012 2177 5148 2183
rect 84 2157 172 2163
rect 180 2157 268 2163
rect 308 2157 380 2163
rect 1844 2157 1948 2163
rect 2020 2157 2220 2163
rect 2244 2157 2332 2163
rect 2932 2157 3260 2163
rect 3268 2157 3340 2163
rect 3380 2157 3964 2163
rect 3997 2157 4076 2163
rect 100 2137 156 2143
rect 164 2137 188 2143
rect 372 2137 396 2143
rect 644 2137 892 2143
rect 932 2137 972 2143
rect 1300 2137 1580 2143
rect 1604 2137 1692 2143
rect 1805 2137 1884 2143
rect 1805 2124 1811 2137
rect 1892 2137 1964 2143
rect 2004 2137 2092 2143
rect 2212 2137 2860 2143
rect 3124 2137 3324 2143
rect 3812 2137 3852 2143
rect 3997 2143 4003 2157
rect 4372 2157 4444 2163
rect 4468 2157 4476 2163
rect 5140 2157 5308 2163
rect 3956 2137 4003 2143
rect 4020 2137 4524 2143
rect 4548 2137 4556 2143
rect 4628 2137 4659 2143
rect 4653 2124 4659 2137
rect 5284 2137 5420 2143
rect 180 2117 348 2123
rect 404 2117 444 2123
rect 484 2117 764 2123
rect 884 2117 924 2123
rect 1556 2117 1612 2123
rect 1620 2117 1804 2123
rect 1844 2117 1916 2123
rect 1988 2117 2044 2123
rect 2228 2117 2460 2123
rect 2772 2117 3180 2123
rect 3316 2117 3356 2123
rect 3684 2117 3724 2123
rect 3732 2117 3916 2123
rect 3924 2117 3980 2123
rect 4100 2117 4156 2123
rect 4356 2117 4636 2123
rect 4724 2117 4780 2123
rect 4788 2117 4876 2123
rect 4980 2117 5068 2123
rect 5076 2117 5180 2123
rect 5364 2117 5404 2123
rect 276 2097 380 2103
rect 468 2097 524 2103
rect 724 2097 812 2103
rect 1012 2097 1084 2103
rect 1524 2097 1660 2103
rect 2068 2097 2172 2103
rect 2260 2097 2396 2103
rect 2420 2097 2668 2103
rect 3476 2097 3500 2103
rect 3588 2097 3756 2103
rect 3828 2097 4124 2103
rect 4292 2097 4476 2103
rect 4500 2097 4748 2103
rect 132 2077 252 2083
rect 436 2077 620 2083
rect 692 2077 1052 2083
rect 1924 2077 2028 2083
rect 2292 2077 2332 2083
rect 2404 2077 2428 2083
rect 3652 2077 3708 2083
rect 3716 2077 3756 2083
rect 3764 2077 3804 2083
rect 3828 2077 4028 2083
rect 4084 2077 4108 2083
rect 4148 2077 4444 2083
rect 4468 2077 4492 2083
rect 244 2057 428 2063
rect 452 2057 636 2063
rect 2260 2057 2284 2063
rect 2324 2057 2348 2063
rect 2484 2057 2556 2063
rect 3812 2057 4044 2063
rect 4052 2057 4172 2063
rect 4180 2057 4556 2063
rect 4564 2057 4780 2063
rect 4788 2057 4892 2063
rect 388 2037 748 2043
rect 2148 2037 2508 2043
rect 2516 2037 2924 2043
rect 3700 2037 3996 2043
rect 4420 2037 4588 2043
rect 4596 2037 5228 2043
rect 436 2017 508 2023
rect 612 2017 636 2023
rect 2596 2017 2604 2023
rect 3892 2017 4140 2023
rect 4612 2017 4620 2023
rect 5188 2017 5228 2023
rect 1218 2014 1278 2016
rect 1218 2006 1219 2014
rect 1228 2006 1229 2014
rect 1267 2006 1268 2014
rect 1277 2006 1278 2014
rect 1218 2004 1278 2006
rect 4226 2014 4286 2016
rect 4226 2006 4227 2014
rect 4236 2006 4237 2014
rect 4275 2006 4276 2014
rect 4285 2006 4286 2014
rect 4226 2004 4286 2006
rect 340 1997 620 2003
rect 644 1997 700 2003
rect 740 1997 940 2003
rect 996 1997 1004 2003
rect 1508 1997 1756 2003
rect 3428 1997 3484 2003
rect 3956 1997 4108 2003
rect 4436 1997 4652 2003
rect 4820 1997 5004 2003
rect 500 1977 572 1983
rect 580 1977 828 1983
rect 996 1977 1100 1983
rect 1812 1977 1836 1983
rect 3796 1977 4188 1983
rect 4692 1977 4892 1983
rect 324 1957 540 1963
rect 964 1957 988 1963
rect 1428 1957 2956 1963
rect 3348 1957 4588 1963
rect 324 1937 332 1943
rect 468 1937 524 1943
rect 2196 1937 2252 1943
rect 2292 1937 3372 1943
rect 3540 1937 3900 1943
rect 3924 1937 3948 1943
rect 4020 1937 4076 1943
rect 4132 1937 4156 1943
rect 4196 1937 4339 1943
rect 4333 1924 4339 1937
rect 4468 1937 4604 1943
rect 4612 1937 4636 1943
rect 68 1917 108 1923
rect 356 1917 588 1923
rect 596 1917 668 1923
rect 916 1917 1292 1923
rect 1300 1917 1484 1923
rect 2292 1917 2316 1923
rect 2324 1917 2476 1923
rect 2484 1917 2828 1923
rect 3780 1917 4012 1923
rect 4116 1917 4140 1923
rect 4148 1917 4236 1923
rect 4340 1917 4364 1923
rect 5012 1917 5164 1923
rect 5204 1917 5324 1923
rect 5332 1917 5468 1923
rect 52 1897 60 1903
rect 68 1897 220 1903
rect 500 1897 812 1903
rect 1764 1897 1916 1903
rect 2196 1897 2236 1903
rect 2356 1897 2524 1903
rect 2532 1897 2684 1903
rect 3380 1897 3756 1903
rect 3764 1897 3788 1903
rect 3892 1897 3980 1903
rect 4052 1897 4348 1903
rect 4676 1897 4812 1903
rect 5044 1897 5116 1903
rect 5140 1897 5500 1903
rect 20 1877 172 1883
rect 276 1877 348 1883
rect 660 1877 796 1883
rect 1236 1877 1324 1883
rect 2196 1877 2300 1883
rect 2308 1877 2380 1883
rect 2676 1877 2876 1883
rect 3460 1877 3596 1883
rect 3876 1877 3996 1883
rect 4020 1877 4099 1883
rect 100 1857 140 1863
rect 148 1857 220 1863
rect 228 1857 300 1863
rect 452 1857 476 1863
rect 500 1857 572 1863
rect 580 1857 924 1863
rect 1604 1857 1676 1863
rect 2228 1857 2300 1863
rect 2500 1857 2620 1863
rect 3364 1857 3388 1863
rect 3396 1857 3420 1863
rect 3428 1857 3436 1863
rect 3444 1857 3596 1863
rect 3604 1857 3804 1863
rect 3860 1857 3948 1863
rect 4068 1857 4076 1863
rect 4093 1863 4099 1877
rect 4116 1877 4332 1883
rect 4340 1877 4476 1883
rect 4596 1877 4620 1883
rect 4756 1877 4988 1883
rect 4996 1877 5052 1883
rect 5156 1877 5180 1883
rect 5188 1877 5388 1883
rect 4093 1857 4124 1863
rect 4324 1857 5004 1863
rect 2244 1837 2684 1843
rect 3636 1837 3804 1843
rect 3812 1837 4348 1843
rect 4356 1837 4860 1843
rect 5220 1837 5420 1843
rect 276 1817 284 1823
rect 532 1817 556 1823
rect 1748 1817 2124 1823
rect 2276 1817 2700 1823
rect 2980 1817 3244 1823
rect 3252 1817 3324 1823
rect 3332 1817 3532 1823
rect 3540 1817 3884 1823
rect 3892 1817 4476 1823
rect 4484 1817 4540 1823
rect 4548 1817 4780 1823
rect 4884 1817 5084 1823
rect 5124 1817 5276 1823
rect 2722 1814 2782 1816
rect 2722 1806 2723 1814
rect 2732 1806 2733 1814
rect 2771 1806 2772 1814
rect 2781 1806 2782 1814
rect 2722 1804 2782 1806
rect 212 1797 284 1803
rect 292 1797 540 1803
rect 2340 1797 2604 1803
rect 3332 1797 4108 1803
rect 4180 1797 4316 1803
rect 4500 1797 4572 1803
rect 4692 1797 4764 1803
rect 4788 1797 4812 1803
rect 4916 1797 5379 1803
rect 244 1777 572 1783
rect 740 1777 828 1783
rect 836 1777 1196 1783
rect 1204 1777 1340 1783
rect 2452 1777 2675 1783
rect 2669 1764 2675 1777
rect 2724 1777 3148 1783
rect 3236 1777 3420 1783
rect 3508 1777 3548 1783
rect 3604 1777 3628 1783
rect 3684 1777 3708 1783
rect 3924 1777 4012 1783
rect 4020 1777 4460 1783
rect 5373 1783 5379 1797
rect 5396 1797 5452 1803
rect 5549 1783 5555 1803
rect 5373 1777 5555 1783
rect 52 1757 92 1763
rect 116 1757 220 1763
rect 228 1757 380 1763
rect 436 1757 764 1763
rect 868 1757 908 1763
rect 1652 1757 1932 1763
rect 2004 1757 2284 1763
rect 2452 1757 2476 1763
rect 2676 1757 2908 1763
rect 3044 1757 3340 1763
rect 3492 1757 3532 1763
rect 4612 1757 4684 1763
rect 4708 1757 4860 1763
rect 4980 1757 5020 1763
rect 5332 1757 5555 1763
rect 212 1737 300 1743
rect 372 1737 428 1743
rect 948 1737 1004 1743
rect 1060 1737 1372 1743
rect 1796 1737 1868 1743
rect 2228 1737 2380 1743
rect 2468 1737 2572 1743
rect 2660 1737 2732 1743
rect 2836 1737 2892 1743
rect 3028 1737 3564 1743
rect 4020 1737 4044 1743
rect 4644 1737 4716 1743
rect 4788 1737 5020 1743
rect 5028 1737 5052 1743
rect 5076 1737 5132 1743
rect 100 1717 332 1723
rect 340 1717 460 1723
rect 980 1717 1068 1723
rect 1652 1717 1676 1723
rect 1684 1717 2188 1723
rect 2196 1717 2380 1723
rect 2420 1717 2524 1723
rect 2628 1717 2700 1723
rect 2708 1717 2844 1723
rect 4068 1717 4108 1723
rect 4660 1717 4716 1723
rect 4724 1717 4780 1723
rect 4788 1717 4812 1723
rect 4820 1717 4972 1723
rect 5060 1717 5100 1723
rect 5236 1717 5260 1723
rect 164 1697 492 1703
rect 1476 1697 1532 1703
rect 1972 1697 1996 1703
rect 2413 1703 2419 1716
rect 2004 1697 2419 1703
rect 2516 1697 2572 1703
rect 2884 1697 2924 1703
rect 3092 1697 3292 1703
rect 3428 1697 3484 1703
rect 3492 1697 4076 1703
rect 4580 1697 4700 1703
rect 4708 1697 4828 1703
rect 4836 1697 4956 1703
rect 4964 1697 5324 1703
rect 5373 1697 5555 1703
rect 884 1677 956 1683
rect 2308 1677 2652 1683
rect 2660 1677 2860 1683
rect 3284 1677 3500 1683
rect 3988 1677 4028 1683
rect 4804 1677 4844 1683
rect 4868 1677 4892 1683
rect 4900 1677 4940 1683
rect 5373 1683 5379 1697
rect 4980 1677 5379 1683
rect 308 1657 412 1663
rect 2356 1657 2588 1663
rect 3348 1657 3971 1663
rect 292 1637 348 1643
rect 356 1637 588 1643
rect 2196 1637 2364 1643
rect 2388 1637 3116 1643
rect 3965 1643 3971 1657
rect 3988 1657 4668 1663
rect 4692 1657 4748 1663
rect 4772 1657 4908 1663
rect 5044 1657 5100 1663
rect 3965 1637 3996 1643
rect 4084 1637 4595 1643
rect 452 1617 572 1623
rect 580 1617 908 1623
rect 2212 1617 2428 1623
rect 2436 1617 2460 1623
rect 3908 1617 3964 1623
rect 4589 1623 4595 1637
rect 4628 1637 4684 1643
rect 4765 1643 4771 1656
rect 4692 1637 4771 1643
rect 5028 1637 5084 1643
rect 4589 1617 5116 1623
rect 1218 1614 1278 1616
rect 1218 1606 1219 1614
rect 1228 1606 1229 1614
rect 1267 1606 1268 1614
rect 1277 1606 1278 1614
rect 1218 1604 1278 1606
rect 4226 1614 4286 1616
rect 4226 1606 4227 1614
rect 4236 1606 4237 1614
rect 4275 1606 4276 1614
rect 4285 1606 4286 1614
rect 4226 1604 4286 1606
rect 3572 1597 4060 1603
rect 4532 1597 4620 1603
rect 4660 1597 4956 1603
rect 52 1577 1196 1583
rect 2404 1577 2412 1583
rect 2420 1577 2908 1583
rect 3524 1577 3724 1583
rect 3812 1577 3980 1583
rect 4157 1577 4636 1583
rect 436 1557 636 1563
rect 1044 1557 1084 1563
rect 1108 1557 1212 1563
rect 1220 1557 1452 1563
rect 3380 1557 3756 1563
rect 4157 1563 4163 1577
rect 4644 1577 4812 1583
rect 3796 1557 4163 1563
rect 4180 1557 4332 1563
rect 4340 1557 4588 1563
rect 4596 1557 4876 1563
rect 84 1537 252 1543
rect 372 1537 428 1543
rect 436 1537 444 1543
rect 516 1537 604 1543
rect 820 1537 1148 1543
rect 2564 1537 2716 1543
rect 2724 1537 2796 1543
rect 3348 1537 3692 1543
rect 3956 1537 3980 1543
rect 3988 1537 4044 1543
rect 4084 1537 4556 1543
rect 4644 1537 4723 1543
rect 4717 1524 4723 1537
rect 4884 1537 4940 1543
rect 4996 1537 5068 1543
rect 5076 1537 5116 1543
rect 5172 1537 5196 1543
rect 36 1517 44 1523
rect 52 1517 60 1523
rect 148 1517 188 1523
rect 196 1517 364 1523
rect 532 1517 652 1523
rect 660 1517 1020 1523
rect 1028 1517 1068 1523
rect 1844 1517 1884 1523
rect 2020 1517 2156 1523
rect 2164 1517 3036 1523
rect 3300 1517 3404 1523
rect 3460 1517 3516 1523
rect 3524 1517 3628 1523
rect 3716 1517 3820 1523
rect 3828 1517 3884 1523
rect 3972 1517 4092 1523
rect 4148 1517 4236 1523
rect 4468 1517 4540 1523
rect 4628 1517 4700 1523
rect 4724 1517 4796 1523
rect 4877 1517 5084 1523
rect 4877 1504 4883 1517
rect 5108 1517 5452 1523
rect -35 1497 12 1503
rect 84 1497 172 1503
rect 180 1497 284 1503
rect 1204 1497 1356 1503
rect 1764 1497 1932 1503
rect 1940 1497 2044 1503
rect 2052 1497 2076 1503
rect 2228 1497 2252 1503
rect 2612 1497 2700 1503
rect 2708 1497 2812 1503
rect 2964 1497 3372 1503
rect 3444 1497 3500 1503
rect 3508 1497 3532 1503
rect 3540 1497 3564 1503
rect 3684 1497 3788 1503
rect 3844 1497 3868 1503
rect 3940 1497 4012 1503
rect 4020 1497 4076 1503
rect 4180 1497 4252 1503
rect 4500 1497 4508 1503
rect 4532 1497 4556 1503
rect 4692 1497 4876 1503
rect 5012 1497 5036 1503
rect 5044 1497 5164 1503
rect 5524 1497 5555 1503
rect 404 1477 412 1483
rect 596 1477 620 1483
rect 660 1477 908 1483
rect 1620 1477 1932 1483
rect 1972 1477 2060 1483
rect 2068 1477 2156 1483
rect 2356 1477 2620 1483
rect 2676 1477 2876 1483
rect 3156 1477 3292 1483
rect 3492 1477 3644 1483
rect 3876 1477 4012 1483
rect 4020 1477 4188 1483
rect 4532 1477 5100 1483
rect 5124 1477 5180 1483
rect 324 1457 396 1463
rect 404 1457 508 1463
rect 676 1457 732 1463
rect 740 1457 876 1463
rect 1172 1457 1180 1463
rect 1732 1457 1948 1463
rect 2036 1457 2076 1463
rect 2084 1457 2108 1463
rect 2628 1457 2636 1463
rect 2644 1457 2668 1463
rect 2676 1457 3308 1463
rect 3764 1457 3836 1463
rect 3940 1457 4124 1463
rect 4132 1457 4540 1463
rect 4548 1457 4620 1463
rect 4868 1457 4892 1463
rect 4916 1457 4972 1463
rect 5156 1457 5244 1463
rect 980 1437 1164 1443
rect 1444 1437 1468 1443
rect 1620 1437 1804 1443
rect 3220 1437 3436 1443
rect 3972 1437 4012 1443
rect 4020 1437 4156 1443
rect 4180 1437 4204 1443
rect 4516 1437 5308 1443
rect 132 1417 284 1423
rect 292 1417 716 1423
rect 900 1417 988 1423
rect 996 1417 1052 1423
rect 2340 1417 2492 1423
rect 3108 1417 3324 1423
rect 3332 1417 3388 1423
rect 3716 1417 4540 1423
rect 4644 1417 4748 1423
rect 4788 1417 4828 1423
rect 5044 1417 5356 1423
rect 2722 1414 2782 1416
rect 2722 1406 2723 1414
rect 2732 1406 2733 1414
rect 2771 1406 2772 1414
rect 2781 1406 2782 1414
rect 2722 1404 2782 1406
rect 212 1397 236 1403
rect 1012 1397 1020 1403
rect 2292 1397 2508 1403
rect 3188 1397 3452 1403
rect 3748 1397 4428 1403
rect 4820 1397 4892 1403
rect 5332 1397 5340 1403
rect 36 1377 76 1383
rect 84 1377 332 1383
rect 3149 1377 4412 1383
rect 3149 1364 3155 1377
rect 84 1357 156 1363
rect 164 1357 364 1363
rect 788 1357 844 1363
rect 852 1357 924 1363
rect 932 1357 1116 1363
rect 1156 1357 1340 1363
rect 1428 1357 1452 1363
rect 2420 1357 2428 1363
rect 2468 1357 2524 1363
rect 2580 1357 2732 1363
rect 2740 1357 3148 1363
rect 3204 1357 3484 1363
rect 3572 1357 3612 1363
rect 3636 1357 3708 1363
rect 3732 1357 3852 1363
rect 4132 1357 4268 1363
rect 4276 1357 4812 1363
rect 68 1337 188 1343
rect 196 1337 332 1343
rect 420 1337 700 1343
rect 1236 1337 1516 1343
rect 1620 1337 1660 1343
rect 1684 1337 1724 1343
rect 2036 1337 2188 1343
rect 2276 1337 2316 1343
rect 2388 1337 2492 1343
rect 2500 1337 2524 1343
rect 2532 1337 2604 1343
rect 2932 1337 3068 1343
rect 3620 1337 3644 1343
rect 3668 1337 3756 1343
rect 3764 1337 3948 1343
rect 4132 1337 4220 1343
rect 4436 1337 4700 1343
rect 52 1317 92 1323
rect 180 1317 268 1323
rect 292 1317 348 1323
rect 356 1317 483 1323
rect 477 1304 483 1317
rect 980 1317 1116 1323
rect 1604 1317 1628 1323
rect 1636 1317 1836 1323
rect 1844 1317 2172 1323
rect 2308 1317 2332 1323
rect 2548 1317 2636 1323
rect 3108 1317 3148 1323
rect 3364 1317 3676 1323
rect 3828 1317 4396 1323
rect 4404 1317 4556 1323
rect 5012 1317 5068 1323
rect 388 1297 444 1303
rect 484 1297 588 1303
rect 596 1297 860 1303
rect 1572 1297 1692 1303
rect 1732 1297 1788 1303
rect 1796 1297 1932 1303
rect 1940 1297 2204 1303
rect 2212 1297 2220 1303
rect 2228 1297 2332 1303
rect 2500 1297 2604 1303
rect 3076 1297 3164 1303
rect 3364 1297 3596 1303
rect 3604 1297 3980 1303
rect 4116 1297 4364 1303
rect 4500 1297 4812 1303
rect 4980 1297 5132 1303
rect 5140 1297 5196 1303
rect 228 1277 252 1283
rect 260 1277 316 1283
rect 340 1277 412 1283
rect 1604 1277 1644 1283
rect 1860 1277 1900 1283
rect 2324 1277 2748 1283
rect 3892 1277 4476 1283
rect 4548 1277 4700 1283
rect 228 1257 268 1263
rect 1165 1257 2956 1263
rect 1165 1244 1171 1257
rect 4260 1257 4540 1263
rect 5060 1257 5068 1263
rect 3188 1237 3372 1243
rect 4036 1237 4620 1243
rect 52 1217 204 1223
rect 868 1217 940 1223
rect 948 1217 1196 1223
rect 1652 1217 1964 1223
rect 1972 1217 1996 1223
rect 3796 1217 3820 1223
rect 3956 1217 4076 1223
rect 1218 1214 1278 1216
rect 1218 1206 1219 1214
rect 1228 1206 1229 1214
rect 1267 1206 1268 1214
rect 1277 1206 1278 1214
rect 1218 1204 1278 1206
rect 4226 1214 4286 1216
rect 4226 1206 4227 1214
rect 4236 1206 4237 1214
rect 4275 1206 4276 1214
rect 4285 1206 4286 1214
rect 4226 1204 4286 1206
rect 468 1197 572 1203
rect 612 1197 668 1203
rect 2148 1197 2668 1203
rect 3540 1197 3580 1203
rect 3908 1197 4204 1203
rect 4324 1197 4556 1203
rect 5156 1197 5420 1203
rect 1012 1177 1020 1183
rect 2228 1177 2508 1183
rect 3780 1177 4428 1183
rect 164 1157 204 1163
rect 212 1157 684 1163
rect 1604 1157 1804 1163
rect 1812 1157 2140 1163
rect 3652 1157 3932 1163
rect 4164 1157 4924 1163
rect 148 1137 188 1143
rect 196 1137 284 1143
rect 1652 1137 1788 1143
rect 1796 1137 1964 1143
rect 2468 1137 2524 1143
rect 3732 1137 4604 1143
rect 4852 1137 4876 1143
rect 4884 1137 5004 1143
rect 5060 1137 5132 1143
rect 68 1117 108 1123
rect 180 1117 252 1123
rect 276 1117 316 1123
rect 836 1117 908 1123
rect 916 1117 1308 1123
rect 1348 1117 1676 1123
rect 2132 1117 2396 1123
rect 3140 1117 3180 1123
rect 3213 1117 3852 1123
rect 3213 1104 3219 1117
rect 4052 1117 4140 1123
rect 4212 1117 4396 1123
rect 4564 1117 4716 1123
rect 4740 1117 4956 1123
rect 4980 1117 5036 1123
rect 5044 1117 5052 1123
rect 148 1097 220 1103
rect 708 1097 876 1103
rect 1172 1097 1276 1103
rect 1492 1097 1548 1103
rect 1684 1097 1708 1103
rect 2212 1097 2252 1103
rect 2372 1097 2556 1103
rect 2564 1097 2588 1103
rect 2756 1097 3212 1103
rect 3700 1097 3788 1103
rect 3796 1097 4124 1103
rect 4180 1097 4316 1103
rect 4372 1097 4476 1103
rect 4580 1097 4620 1103
rect 4644 1097 4668 1103
rect 4772 1097 4780 1103
rect 4788 1097 4796 1103
rect 4836 1097 4908 1103
rect 52 1077 76 1083
rect 420 1077 524 1083
rect 532 1077 588 1083
rect 804 1077 844 1083
rect 1460 1077 1484 1083
rect 1492 1077 1548 1083
rect 1748 1077 1836 1083
rect 1940 1077 2156 1083
rect 2468 1077 2492 1083
rect 2500 1077 2508 1083
rect 2948 1077 3164 1083
rect 3524 1077 3772 1083
rect 4004 1077 4060 1083
rect 4244 1077 4332 1083
rect 4468 1077 4492 1083
rect 4596 1077 4732 1083
rect 4836 1077 4860 1083
rect 4868 1077 4924 1083
rect 4996 1077 5148 1083
rect 340 1057 636 1063
rect 1012 1057 1148 1063
rect 1412 1057 1468 1063
rect 1476 1057 1484 1063
rect 1748 1057 1772 1063
rect 1780 1057 2076 1063
rect 2132 1057 2252 1063
rect 2340 1057 2364 1063
rect 2404 1057 2444 1063
rect 2452 1057 2572 1063
rect 2916 1057 3116 1063
rect 3124 1057 3244 1063
rect 3252 1057 3388 1063
rect 3396 1057 3548 1063
rect 3636 1057 3916 1063
rect 3972 1057 4044 1063
rect 4084 1057 4524 1063
rect 4724 1057 4812 1063
rect 4820 1057 4892 1063
rect 4916 1057 5004 1063
rect 5124 1057 5372 1063
rect 820 1037 972 1043
rect 1412 1037 1612 1043
rect 1620 1037 1756 1043
rect 2260 1037 2540 1043
rect 2548 1037 3036 1043
rect 3140 1037 3724 1043
rect 3860 1037 3948 1043
rect 4324 1037 4460 1043
rect 324 1017 444 1023
rect 1444 1017 1452 1023
rect 1460 1017 1500 1023
rect 2356 1017 2508 1023
rect 3700 1017 3740 1023
rect 3956 1017 4220 1023
rect 4420 1017 4684 1023
rect 2722 1014 2782 1016
rect 2722 1006 2723 1014
rect 2732 1006 2733 1014
rect 2771 1006 2772 1014
rect 2781 1006 2782 1014
rect 2722 1004 2782 1006
rect 1044 997 1084 1003
rect 1396 997 1884 1003
rect 1892 997 2220 1003
rect 2468 997 2620 1003
rect 2868 997 2908 1003
rect 3204 997 3212 1003
rect 3380 997 3420 1003
rect 3716 997 3836 1003
rect 3940 997 4460 1003
rect 4532 997 4668 1003
rect 5044 997 5372 1003
rect 292 977 332 983
rect 340 977 428 983
rect 436 977 444 983
rect 468 977 492 983
rect 1540 977 1740 983
rect 1748 977 1836 983
rect 2100 977 2188 983
rect 2260 977 2284 983
rect 2628 977 3084 983
rect 3684 977 4092 983
rect 4164 977 4556 983
rect 4596 977 4748 983
rect 4788 977 5020 983
rect 5028 977 5084 983
rect 5092 977 5180 983
rect 148 957 236 963
rect 404 957 460 963
rect 804 957 876 963
rect 1380 957 1420 963
rect 2084 957 2220 963
rect 2276 957 2348 963
rect 2436 957 2492 963
rect 2500 957 2604 963
rect 3044 957 3068 963
rect 3556 957 3708 963
rect 3908 957 4099 963
rect 164 937 300 943
rect 516 937 524 943
rect 596 937 908 943
rect 1124 937 1356 943
rect 2052 937 2124 943
rect 2196 937 2236 943
rect 2260 937 2284 943
rect 2324 937 2364 943
rect 2644 937 2892 943
rect 3284 937 3452 943
rect 3540 937 3964 943
rect 3988 937 4028 943
rect 4036 937 4044 943
rect 4093 943 4099 957
rect 4116 957 4380 963
rect 4388 957 4524 963
rect 4660 957 4684 963
rect 4996 957 5340 963
rect 4093 937 4380 943
rect 4420 937 4588 943
rect 4660 937 4796 943
rect 212 917 236 923
rect 276 917 396 923
rect 836 917 876 923
rect 884 917 908 923
rect 916 917 956 923
rect 980 917 1004 923
rect 1508 917 1532 923
rect 1716 917 1756 923
rect 1764 917 1804 923
rect 2125 917 2412 923
rect 2125 904 2131 917
rect 2420 917 2476 923
rect 2484 917 2572 923
rect 3156 917 3436 923
rect 3444 917 3484 923
rect 3508 917 3516 923
rect 3524 917 3532 923
rect 3908 917 4156 923
rect 4228 917 4492 923
rect 4644 917 4876 923
rect 5124 917 5260 923
rect 20 897 156 903
rect 164 897 172 903
rect 180 897 220 903
rect 244 897 412 903
rect 1540 897 1612 903
rect 2004 897 2124 903
rect 2228 897 2268 903
rect 3876 897 3900 903
rect 3908 897 3932 903
rect 3972 897 4044 903
rect 4084 897 4124 903
rect 4132 897 4492 903
rect 4500 897 4556 903
rect 4564 897 4684 903
rect 4740 897 4780 903
rect 52 877 124 883
rect 132 877 188 883
rect 212 877 252 883
rect 308 877 380 883
rect 1556 877 1612 883
rect 2052 877 2380 883
rect 3860 877 4396 883
rect 1860 857 2636 863
rect 4036 857 4172 863
rect 4180 857 4300 863
rect 4372 857 4428 863
rect 3268 837 3420 843
rect 3796 837 4188 843
rect 4340 837 4412 843
rect 4436 837 4444 843
rect 164 817 300 823
rect 628 817 652 823
rect 2612 817 3100 823
rect 3108 817 3164 823
rect 4372 817 4460 823
rect 5428 817 5452 823
rect 1218 814 1278 816
rect 1218 806 1219 814
rect 1228 806 1229 814
rect 1267 806 1268 814
rect 1277 806 1278 814
rect 1218 804 1278 806
rect 4226 814 4286 816
rect 4226 806 4227 814
rect 4236 806 4237 814
rect 4275 806 4276 814
rect 4285 806 4286 814
rect 4226 804 4286 806
rect 1348 797 1452 803
rect 1860 797 1932 803
rect 2292 797 2316 803
rect 2868 797 2908 803
rect 3092 797 3788 803
rect 3220 777 3276 783
rect 4676 777 4844 783
rect 3060 757 3260 763
rect 3348 757 3724 763
rect 4980 757 4988 763
rect 5044 757 5068 763
rect 5076 757 5148 763
rect 84 737 524 743
rect 532 737 844 743
rect 2292 737 2476 743
rect 2484 737 3132 743
rect 3588 737 3756 743
rect 3780 737 3916 743
rect 4484 737 4508 743
rect 4852 737 5100 743
rect 372 717 396 723
rect 1636 717 1676 723
rect 1684 717 1772 723
rect 2532 717 2572 723
rect 2580 717 3107 723
rect 3101 704 3107 717
rect 3316 717 3852 723
rect 3924 717 3964 723
rect 4260 717 4700 723
rect 4916 717 5036 723
rect 5044 717 5052 723
rect 5060 717 5084 723
rect 100 697 124 703
rect 228 697 268 703
rect 292 697 460 703
rect 500 697 540 703
rect 788 697 876 703
rect 884 697 1164 703
rect 1172 697 1308 703
rect 1972 697 2108 703
rect 2116 697 2172 703
rect 2740 697 3084 703
rect 3108 697 3148 703
rect 3188 697 3228 703
rect 3236 697 3356 703
rect 3700 697 3740 703
rect 3748 697 3884 703
rect 4468 697 4540 703
rect 4612 697 4908 703
rect 4932 697 4972 703
rect 5012 697 5100 703
rect 68 677 300 683
rect 324 677 428 683
rect 628 677 748 683
rect 772 677 780 683
rect 1124 677 1340 683
rect 1540 677 1596 683
rect 2468 677 2700 683
rect 2708 677 2828 683
rect 2836 677 3212 683
rect 3284 677 3804 683
rect 3876 677 3932 683
rect 4004 677 4588 683
rect 4660 677 4748 683
rect 4836 677 5020 683
rect 5108 677 5164 683
rect 36 657 188 663
rect 356 657 396 663
rect 884 657 1084 663
rect 1092 657 1500 663
rect 1508 657 1644 663
rect 1652 657 1884 663
rect 1892 657 1980 663
rect 1988 657 2252 663
rect 2436 657 2620 663
rect 2644 657 2668 663
rect 2948 657 3116 663
rect 3204 657 3244 663
rect 3396 657 3708 663
rect 4500 657 4588 663
rect 5044 657 5356 663
rect 260 637 364 643
rect 388 637 444 643
rect 2564 637 2940 643
rect 3044 637 3212 643
rect 3364 637 3548 643
rect 3956 637 4044 643
rect 4484 637 4508 643
rect 4564 637 4796 643
rect 308 617 348 623
rect 3380 617 3436 623
rect 3444 617 3676 623
rect 3684 617 3772 623
rect 3812 617 4499 623
rect 2722 614 2782 616
rect 2722 606 2723 614
rect 2732 606 2733 614
rect 2771 606 2772 614
rect 2781 606 2782 614
rect 2722 604 2782 606
rect 500 597 556 603
rect 1332 597 1715 603
rect 1709 584 1715 597
rect 2148 597 2188 603
rect 2196 597 2300 603
rect 2308 597 2492 603
rect 2916 597 2972 603
rect 3284 597 3843 603
rect 116 577 220 583
rect 820 577 1388 583
rect 1396 577 1692 583
rect 1716 577 2428 583
rect 3332 577 3676 583
rect 3837 583 3843 597
rect 3860 597 3916 603
rect 4493 603 4499 617
rect 4516 617 4540 623
rect 4493 597 4604 603
rect 4676 597 4876 603
rect 3837 577 4716 583
rect 4948 577 5004 583
rect 5012 577 5068 583
rect 52 557 92 563
rect 100 557 124 563
rect 212 557 300 563
rect 1044 557 1356 563
rect 1380 557 1436 563
rect 1460 557 1596 563
rect 2356 557 2556 563
rect 3252 557 3532 563
rect 3540 557 3548 563
rect 3588 557 3724 563
rect 3732 557 4188 563
rect 4212 557 4332 563
rect 4349 557 4620 563
rect 20 537 28 543
rect 36 537 44 543
rect 116 537 172 543
rect 244 537 316 543
rect 324 537 460 543
rect 1316 537 1628 543
rect 1636 537 1740 543
rect 1748 537 2028 543
rect 2036 537 2476 543
rect 2484 537 3084 543
rect 3188 537 3580 543
rect 3588 537 3692 543
rect 3876 537 4076 543
rect 4116 537 4252 543
rect 4349 543 4355 557
rect 4772 557 4924 563
rect 4932 557 5148 563
rect 4308 537 4355 543
rect 4413 537 4764 543
rect 196 517 268 523
rect 1236 517 1452 523
rect 1460 517 1548 523
rect 1588 517 1612 523
rect 1620 517 1628 523
rect 1908 517 2156 523
rect 2228 517 2268 523
rect 2276 517 2364 523
rect 3556 517 3596 523
rect 3604 517 3628 523
rect 3652 517 3692 523
rect 4132 517 4172 523
rect 4413 523 4419 537
rect 4980 537 5020 543
rect 5124 537 5340 543
rect 4196 517 4419 523
rect 4500 517 4828 523
rect 4852 517 5084 523
rect 5108 517 5340 523
rect 52 497 156 503
rect 164 497 252 503
rect 1348 497 1484 503
rect 1780 497 1804 503
rect 2260 497 2332 503
rect 2404 497 2620 503
rect 2628 497 2796 503
rect 2804 497 2844 503
rect 2852 497 3148 503
rect 3700 497 4364 503
rect 5220 497 5308 503
rect 5316 497 5468 503
rect 4164 477 4188 483
rect 4308 477 4476 483
rect 4340 457 4780 463
rect 5044 457 5068 463
rect 548 437 572 443
rect 1668 417 1692 423
rect 1860 417 1932 423
rect 2484 417 2524 423
rect 4660 417 4684 423
rect 1218 414 1278 416
rect 1218 406 1219 414
rect 1228 406 1229 414
rect 1267 406 1268 414
rect 1277 406 1278 414
rect 1218 404 1278 406
rect 4226 414 4286 416
rect 4226 406 4227 414
rect 4236 406 4237 414
rect 4275 406 4276 414
rect 4285 406 4286 414
rect 4226 404 4286 406
rect 228 397 268 403
rect 1636 397 1660 403
rect 1668 397 1788 403
rect 1812 397 1948 403
rect 4836 377 4876 383
rect 5316 377 5324 383
rect 1364 337 4076 343
rect 4772 337 4796 343
rect 5284 337 5420 343
rect 2084 317 2188 323
rect 2228 317 2268 323
rect 4884 317 5180 323
rect 5236 317 5324 323
rect 324 297 460 303
rect 756 297 796 303
rect 1156 297 1196 303
rect 1204 297 1628 303
rect 2132 297 2220 303
rect 2708 297 2812 303
rect 2884 297 3244 303
rect 4772 297 5244 303
rect 564 277 572 283
rect 1892 277 2044 283
rect 2708 277 2796 283
rect 2804 277 2860 283
rect 2884 277 3084 283
rect 4036 277 5180 283
rect 2244 257 2268 263
rect 2484 257 3052 263
rect 4500 257 4684 263
rect 4692 257 4828 263
rect 4836 257 4988 263
rect 4996 257 5212 263
rect 932 237 1196 243
rect 1236 237 1356 243
rect 1540 237 2348 243
rect 2516 237 2716 243
rect 4724 237 4972 243
rect 4980 237 4988 243
rect 5012 237 5020 243
rect 612 217 668 223
rect 676 217 908 223
rect 916 217 940 223
rect 1012 217 1068 223
rect 1076 217 1500 223
rect 1508 217 1548 223
rect 1556 217 1852 223
rect 1860 217 1980 223
rect 2036 217 2332 223
rect 2452 217 2700 223
rect 3364 217 3436 223
rect 3684 217 3772 223
rect 3908 217 3980 223
rect 4292 217 4332 223
rect 2722 214 2782 216
rect 2722 206 2723 214
rect 2732 206 2733 214
rect 2771 206 2772 214
rect 2781 206 2782 214
rect 2722 204 2782 206
rect 36 197 92 203
rect 1044 197 1212 203
rect 2628 197 2668 203
rect 3076 197 3404 203
rect 3412 197 3548 203
rect 3556 197 3596 203
rect 3604 197 3868 203
rect 2324 177 2380 183
rect 2388 177 2460 183
rect 2468 177 2652 183
rect 2676 177 2892 183
rect 196 157 524 163
rect 532 157 876 163
rect 884 157 1004 163
rect 2404 157 2668 163
rect 3876 157 4124 163
rect 4132 157 4332 163
rect 212 137 220 143
rect 500 137 700 143
rect 836 137 972 143
rect 1428 137 1580 143
rect 1956 137 2236 143
rect 2276 137 2444 143
rect 2564 137 2572 143
rect 2580 137 2636 143
rect 2692 137 2796 143
rect 3092 137 3244 143
rect 3252 137 3308 143
rect 692 117 796 123
rect 1172 117 2252 123
rect 2436 117 2556 123
rect 2660 117 2716 123
rect 2724 117 2908 123
rect 3300 117 3580 123
rect 3972 117 3996 123
rect 4596 117 4620 123
rect 1668 97 1852 103
rect 2228 97 2300 103
rect 2308 97 2492 103
rect 2500 97 2540 103
rect 2548 97 2748 103
rect 2788 97 2876 103
rect 3332 97 3388 103
rect 5524 97 5555 103
rect 2260 77 2284 83
rect 2372 77 2396 83
rect 2548 77 3100 83
rect 3268 37 3292 43
rect 3716 37 5164 43
rect 5172 37 5356 43
rect 3220 17 3260 23
rect 3508 17 3516 23
rect 4532 17 4700 23
rect 1218 14 1278 16
rect 1218 6 1219 14
rect 1228 6 1229 14
rect 1267 6 1268 14
rect 1277 6 1278 14
rect 1218 4 1278 6
rect 4226 14 4286 16
rect 4226 6 4227 14
rect 4236 6 4237 14
rect 4275 6 4276 14
rect 4285 6 4286 14
rect 4226 4 4286 6
<< m4contact >>
rect 2092 3816 2100 3824
rect 2724 3806 2731 3814
rect 2731 3806 2732 3814
rect 2736 3806 2741 3814
rect 2741 3806 2743 3814
rect 2743 3806 2744 3814
rect 2748 3806 2751 3814
rect 2751 3806 2753 3814
rect 2753 3806 2756 3814
rect 2760 3806 2761 3814
rect 2761 3806 2763 3814
rect 2763 3806 2768 3814
rect 2772 3806 2773 3814
rect 2773 3806 2780 3814
rect 268 3736 276 3744
rect 3596 3736 3604 3744
rect 3916 3716 3924 3724
rect 3660 3676 3668 3684
rect 5260 3676 5268 3684
rect 716 3636 724 3644
rect 3244 3636 3252 3644
rect 1220 3606 1227 3614
rect 1227 3606 1228 3614
rect 1232 3606 1237 3614
rect 1237 3606 1239 3614
rect 1239 3606 1240 3614
rect 1244 3606 1247 3614
rect 1247 3606 1249 3614
rect 1249 3606 1252 3614
rect 1256 3606 1257 3614
rect 1257 3606 1259 3614
rect 1259 3606 1264 3614
rect 1268 3606 1269 3614
rect 1269 3606 1276 3614
rect 4228 3606 4235 3614
rect 4235 3606 4236 3614
rect 4240 3606 4245 3614
rect 4245 3606 4247 3614
rect 4247 3606 4248 3614
rect 4252 3606 4255 3614
rect 4255 3606 4257 3614
rect 4257 3606 4260 3614
rect 4264 3606 4265 3614
rect 4265 3606 4267 3614
rect 4267 3606 4272 3614
rect 4276 3606 4277 3614
rect 4277 3606 4284 3614
rect 3980 3576 3988 3584
rect 4428 3576 4436 3584
rect 4428 3536 4436 3544
rect 3724 3496 3732 3504
rect 4108 3496 4116 3504
rect 4492 3496 4500 3504
rect 2860 3456 2868 3464
rect 4652 3456 4660 3464
rect 748 3436 756 3444
rect 2380 3436 2388 3444
rect 4108 3436 4116 3444
rect 5228 3436 5236 3444
rect 5388 3436 5396 3444
rect 2724 3406 2731 3414
rect 2731 3406 2732 3414
rect 2736 3406 2741 3414
rect 2741 3406 2743 3414
rect 2743 3406 2744 3414
rect 2748 3406 2751 3414
rect 2751 3406 2753 3414
rect 2753 3406 2756 3414
rect 2760 3406 2761 3414
rect 2761 3406 2763 3414
rect 2763 3406 2768 3414
rect 2772 3406 2773 3414
rect 2773 3406 2780 3414
rect 812 3396 820 3404
rect 3660 3396 3668 3404
rect 4684 3396 4692 3404
rect 3244 3376 3252 3384
rect 4588 3376 4596 3384
rect 4748 3356 4756 3364
rect 4012 3336 4020 3344
rect 4364 3336 4372 3344
rect 2092 3316 2100 3324
rect 3372 3316 3380 3324
rect 4492 3316 4500 3324
rect 1804 3296 1812 3304
rect 3724 3296 3732 3304
rect 4076 3296 4084 3304
rect 4364 3296 4372 3304
rect 3596 3276 3604 3284
rect 3980 3276 3988 3284
rect 4044 3276 4052 3284
rect 2860 3236 2868 3244
rect 268 3216 276 3224
rect 2380 3216 2388 3224
rect 3756 3216 3764 3224
rect 3916 3216 3924 3224
rect 1220 3206 1227 3214
rect 1227 3206 1228 3214
rect 1232 3206 1237 3214
rect 1237 3206 1239 3214
rect 1239 3206 1240 3214
rect 1244 3206 1247 3214
rect 1247 3206 1249 3214
rect 1249 3206 1252 3214
rect 1256 3206 1257 3214
rect 1257 3206 1259 3214
rect 1259 3206 1264 3214
rect 1268 3206 1269 3214
rect 1269 3206 1276 3214
rect 4228 3206 4235 3214
rect 4235 3206 4236 3214
rect 4240 3206 4245 3214
rect 4245 3206 4247 3214
rect 4247 3206 4248 3214
rect 4252 3206 4255 3214
rect 4255 3206 4257 3214
rect 4257 3206 4260 3214
rect 4264 3206 4265 3214
rect 4265 3206 4267 3214
rect 4267 3206 4272 3214
rect 4276 3206 4277 3214
rect 4277 3206 4284 3214
rect 4748 3176 4756 3184
rect 556 3156 564 3164
rect 3756 3136 3764 3144
rect 780 3076 788 3084
rect 4044 3076 4052 3084
rect 332 3056 340 3064
rect 1772 3056 1780 3064
rect 460 3036 468 3044
rect 684 3036 692 3044
rect 716 3036 724 3044
rect 3660 3036 3668 3044
rect 5036 3036 5044 3044
rect 4940 3016 4948 3024
rect 2724 3006 2731 3014
rect 2731 3006 2732 3014
rect 2736 3006 2741 3014
rect 2741 3006 2743 3014
rect 2743 3006 2744 3014
rect 2748 3006 2751 3014
rect 2751 3006 2753 3014
rect 2753 3006 2756 3014
rect 2760 3006 2761 3014
rect 2761 3006 2763 3014
rect 2763 3006 2768 3014
rect 2772 3006 2773 3014
rect 2773 3006 2780 3014
rect 524 2996 532 3004
rect 1324 2996 1332 3004
rect 1804 2996 1812 3004
rect 5324 2996 5332 3004
rect 3340 2976 3348 2984
rect 3468 2976 3476 2984
rect 140 2956 148 2964
rect 748 2956 756 2964
rect 3852 2956 3860 2964
rect 5356 2956 5364 2964
rect 4780 2936 4788 2944
rect 2412 2916 2420 2924
rect 3212 2916 3220 2924
rect 3372 2916 3380 2924
rect 1900 2896 1908 2904
rect 2348 2896 2356 2904
rect 3852 2916 3860 2924
rect 4428 2916 4436 2924
rect 5004 2916 5012 2924
rect 3756 2896 3764 2904
rect 4012 2896 4020 2904
rect 4076 2896 4084 2904
rect 396 2856 404 2864
rect 1100 2856 1108 2864
rect 748 2836 756 2844
rect 2060 2836 2068 2844
rect 1220 2806 1227 2814
rect 1227 2806 1228 2814
rect 1232 2806 1237 2814
rect 1237 2806 1239 2814
rect 1239 2806 1240 2814
rect 1244 2806 1247 2814
rect 1247 2806 1249 2814
rect 1249 2806 1252 2814
rect 1256 2806 1257 2814
rect 1257 2806 1259 2814
rect 1259 2806 1264 2814
rect 1268 2806 1269 2814
rect 1269 2806 1276 2814
rect 4228 2806 4235 2814
rect 4235 2806 4236 2814
rect 4240 2806 4245 2814
rect 4245 2806 4247 2814
rect 4247 2806 4248 2814
rect 4252 2806 4255 2814
rect 4255 2806 4257 2814
rect 4257 2806 4260 2814
rect 4264 2806 4265 2814
rect 4265 2806 4267 2814
rect 4267 2806 4272 2814
rect 4276 2806 4277 2814
rect 4277 2806 4284 2814
rect 2252 2796 2260 2804
rect 2828 2796 2836 2804
rect 5260 2796 5268 2804
rect 236 2776 244 2784
rect 1580 2776 1588 2784
rect 1740 2756 1748 2764
rect 2156 2756 2164 2764
rect 2956 2756 2964 2764
rect 2476 2736 2484 2744
rect 3532 2736 3540 2744
rect 300 2716 308 2724
rect 4076 2716 4084 2724
rect 396 2696 404 2704
rect 1356 2696 1364 2704
rect 1420 2696 1428 2704
rect 300 2676 308 2684
rect 1324 2676 1332 2684
rect 1548 2676 1556 2684
rect 1772 2676 1780 2684
rect 2892 2676 2900 2684
rect 460 2656 468 2664
rect 556 2656 564 2664
rect 716 2656 724 2664
rect 748 2656 756 2664
rect 3020 2656 3028 2664
rect 1404 2636 1412 2644
rect 1452 2616 1460 2624
rect 4684 2616 4692 2624
rect 2724 2606 2731 2614
rect 2731 2606 2732 2614
rect 2736 2606 2741 2614
rect 2741 2606 2743 2614
rect 2743 2606 2744 2614
rect 2748 2606 2751 2614
rect 2751 2606 2753 2614
rect 2753 2606 2756 2614
rect 2760 2606 2761 2614
rect 2761 2606 2763 2614
rect 2763 2606 2768 2614
rect 2772 2606 2773 2614
rect 2773 2606 2780 2614
rect 1676 2596 1684 2604
rect 1740 2596 1748 2604
rect 4460 2596 4468 2604
rect 236 2576 244 2584
rect 2412 2576 2420 2584
rect 3820 2576 3828 2584
rect 4556 2576 4564 2584
rect 4812 2576 4820 2584
rect 5420 2576 5428 2584
rect 332 2556 340 2564
rect 460 2556 468 2564
rect 2892 2556 2900 2564
rect 4940 2556 4948 2564
rect 1580 2536 1588 2544
rect 140 2516 148 2524
rect 5100 2516 5108 2524
rect 524 2496 532 2504
rect 620 2496 628 2504
rect 684 2496 692 2504
rect 2828 2496 2836 2504
rect 3468 2476 3476 2484
rect 3660 2476 3668 2484
rect 4428 2476 4436 2484
rect 204 2456 212 2464
rect 300 2456 308 2464
rect 3180 2456 3188 2464
rect 3212 2456 3220 2464
rect 1548 2416 1556 2424
rect 1220 2406 1227 2414
rect 1227 2406 1228 2414
rect 1232 2406 1237 2414
rect 1237 2406 1239 2414
rect 1239 2406 1240 2414
rect 1244 2406 1247 2414
rect 1247 2406 1249 2414
rect 1249 2406 1252 2414
rect 1256 2406 1257 2414
rect 1257 2406 1259 2414
rect 1259 2406 1264 2414
rect 1268 2406 1269 2414
rect 1269 2406 1276 2414
rect 4228 2406 4235 2414
rect 4235 2406 4236 2414
rect 4240 2406 4245 2414
rect 4245 2406 4247 2414
rect 4247 2406 4248 2414
rect 4252 2406 4255 2414
rect 4255 2406 4257 2414
rect 4257 2406 4260 2414
rect 4264 2406 4265 2414
rect 4265 2406 4267 2414
rect 4267 2406 4272 2414
rect 4276 2406 4277 2414
rect 4277 2406 4284 2414
rect 1708 2396 1716 2404
rect 2092 2396 2100 2404
rect 2060 2376 2068 2384
rect 3596 2396 3604 2404
rect 3660 2376 3668 2384
rect 1836 2356 1844 2364
rect 5516 2356 5524 2364
rect 1676 2316 1684 2324
rect 1772 2316 1780 2324
rect 460 2296 468 2304
rect 620 2276 628 2284
rect 1324 2276 1332 2284
rect 2604 2276 2612 2284
rect 204 2256 212 2264
rect 332 2256 340 2264
rect 4588 2276 4596 2284
rect 4716 2276 4724 2284
rect 4748 2276 4756 2284
rect 5516 2276 5524 2284
rect 4428 2256 4436 2264
rect 5260 2256 5268 2264
rect 1644 2236 1652 2244
rect 4588 2216 4596 2224
rect 5228 2216 5236 2224
rect 2724 2206 2731 2214
rect 2731 2206 2732 2214
rect 2736 2206 2741 2214
rect 2741 2206 2743 2214
rect 2743 2206 2744 2214
rect 2748 2206 2751 2214
rect 2751 2206 2753 2214
rect 2753 2206 2756 2214
rect 2760 2206 2761 2214
rect 2761 2206 2763 2214
rect 2763 2206 2768 2214
rect 2772 2206 2773 2214
rect 2773 2206 2780 2214
rect 3372 2196 3380 2204
rect 1356 2176 1364 2184
rect 3756 2176 3764 2184
rect 5004 2176 5012 2184
rect 3372 2156 3380 2164
rect 4076 2156 4084 2164
rect 4108 2156 4116 2164
rect 4460 2156 4468 2164
rect 4556 2136 4564 2144
rect 396 2116 404 2124
rect 3980 2116 3988 2124
rect 4652 2116 4660 2124
rect 4876 2116 4884 2124
rect 5356 2116 5364 2124
rect 3500 2096 3508 2104
rect 3756 2096 3764 2104
rect 428 2076 436 2084
rect 684 2076 692 2084
rect 3820 2076 3828 2084
rect 4140 2076 4148 2084
rect 236 2056 244 2064
rect 2252 2056 2260 2064
rect 2316 2056 2324 2064
rect 2348 2056 2356 2064
rect 4556 2056 4564 2064
rect 2508 2036 2516 2044
rect 4588 2036 4596 2044
rect 5228 2036 5236 2044
rect 2604 2016 2612 2024
rect 4140 2016 4148 2024
rect 4620 2016 4628 2024
rect 1220 2006 1227 2014
rect 1227 2006 1228 2014
rect 1232 2006 1237 2014
rect 1237 2006 1239 2014
rect 1239 2006 1240 2014
rect 1244 2006 1247 2014
rect 1247 2006 1249 2014
rect 1249 2006 1252 2014
rect 1256 2006 1257 2014
rect 1257 2006 1259 2014
rect 1259 2006 1264 2014
rect 1268 2006 1269 2014
rect 1269 2006 1276 2014
rect 4228 2006 4235 2014
rect 4235 2006 4236 2014
rect 4240 2006 4245 2014
rect 4245 2006 4247 2014
rect 4247 2006 4248 2014
rect 4252 2006 4255 2014
rect 4255 2006 4257 2014
rect 4257 2006 4260 2014
rect 4264 2006 4265 2014
rect 4265 2006 4267 2014
rect 4267 2006 4272 2014
rect 4276 2006 4277 2014
rect 4277 2006 4284 2014
rect 940 1996 948 2004
rect 1004 1996 1012 2004
rect 3948 1996 3956 2004
rect 5004 1996 5012 2004
rect 492 1976 500 1984
rect 1100 1976 1108 1984
rect 332 1936 340 1944
rect 460 1936 468 1944
rect 2252 1936 2260 1944
rect 2284 1936 2292 1944
rect 3532 1936 3540 1944
rect 4364 1936 4372 1944
rect 2828 1916 2836 1924
rect 5324 1916 5332 1924
rect 812 1896 820 1904
rect 3756 1896 3764 1904
rect 4652 1896 4660 1904
rect 4812 1896 4820 1904
rect 5036 1896 5044 1904
rect 1324 1876 1332 1884
rect 300 1856 308 1864
rect 4076 1856 4084 1864
rect 5388 1876 5396 1884
rect 524 1836 532 1844
rect 268 1816 276 1824
rect 2124 1816 2132 1824
rect 2724 1806 2731 1814
rect 2731 1806 2732 1814
rect 2736 1806 2741 1814
rect 2741 1806 2743 1814
rect 2743 1806 2744 1814
rect 2748 1806 2751 1814
rect 2751 1806 2753 1814
rect 2753 1806 2756 1814
rect 2760 1806 2761 1814
rect 2761 1806 2763 1814
rect 2763 1806 2768 1814
rect 2772 1806 2773 1814
rect 2773 1806 2780 1814
rect 4172 1796 4180 1804
rect 4684 1796 4692 1804
rect 4780 1796 4788 1804
rect 4812 1796 4820 1804
rect 3500 1776 3508 1784
rect 3596 1776 3604 1784
rect 5452 1796 5460 1804
rect 2284 1756 2292 1764
rect 2476 1756 2484 1764
rect 4972 1756 4980 1764
rect 5324 1756 5332 1764
rect 940 1736 948 1744
rect 2828 1736 2836 1744
rect 3020 1736 3028 1744
rect 4012 1736 4020 1744
rect 4716 1736 4724 1744
rect 4780 1736 4788 1744
rect 5260 1716 5268 1724
rect 3084 1696 3092 1704
rect 4076 1696 4084 1704
rect 5324 1696 5332 1704
rect 428 1676 436 1684
rect 876 1676 884 1684
rect 3276 1676 3284 1684
rect 300 1656 308 1664
rect 3340 1656 3348 1664
rect 3980 1656 3988 1664
rect 4972 1656 4980 1664
rect 1220 1606 1227 1614
rect 1227 1606 1228 1614
rect 1232 1606 1237 1614
rect 1237 1606 1239 1614
rect 1239 1606 1240 1614
rect 1244 1606 1247 1614
rect 1247 1606 1249 1614
rect 1249 1606 1252 1614
rect 1256 1606 1257 1614
rect 1257 1606 1259 1614
rect 1259 1606 1264 1614
rect 1268 1606 1269 1614
rect 1269 1606 1276 1614
rect 4228 1606 4235 1614
rect 4235 1606 4236 1614
rect 4240 1606 4245 1614
rect 4245 1606 4247 1614
rect 4247 1606 4248 1614
rect 4252 1606 4255 1614
rect 4255 1606 4257 1614
rect 4257 1606 4260 1614
rect 4264 1606 4265 1614
rect 4265 1606 4267 1614
rect 4267 1606 4272 1614
rect 4276 1606 4277 1614
rect 4277 1606 4284 1614
rect 492 1596 500 1604
rect 4652 1596 4660 1604
rect 2412 1576 2420 1584
rect 3724 1576 3732 1584
rect 3980 1576 3988 1584
rect 428 1536 436 1544
rect 812 1536 820 1544
rect 5196 1536 5204 1544
rect 44 1516 52 1524
rect 2156 1516 2164 1524
rect 4172 1496 4180 1504
rect 4492 1496 4500 1504
rect 4684 1496 4692 1504
rect 5036 1496 5044 1504
rect 396 1476 404 1484
rect 1964 1476 1972 1484
rect 4012 1476 4020 1484
rect 204 1456 212 1464
rect 1164 1456 1172 1464
rect 3756 1456 3764 1464
rect 4620 1456 4628 1464
rect 4748 1416 4756 1424
rect 2724 1406 2731 1414
rect 2731 1406 2732 1414
rect 2736 1406 2741 1414
rect 2741 1406 2743 1414
rect 2743 1406 2744 1414
rect 2748 1406 2751 1414
rect 2751 1406 2753 1414
rect 2753 1406 2756 1414
rect 2760 1406 2761 1414
rect 2761 1406 2763 1414
rect 2763 1406 2768 1414
rect 2772 1406 2773 1414
rect 2773 1406 2780 1414
rect 236 1396 244 1404
rect 1004 1396 1012 1404
rect 2508 1396 2516 1404
rect 4812 1396 4820 1404
rect 5324 1396 5332 1404
rect 1452 1356 1460 1364
rect 2412 1356 2420 1364
rect 3852 1356 3860 1364
rect 2316 1336 2324 1344
rect 3948 1336 3956 1344
rect 5004 1316 5012 1324
rect 1932 1296 1940 1304
rect 4108 1296 4116 1304
rect 1644 1276 1652 1284
rect 1900 1276 1908 1284
rect 2316 1276 2324 1284
rect 268 1256 276 1264
rect 2956 1256 2964 1264
rect 5068 1256 5076 1264
rect 3180 1236 3188 1244
rect 204 1216 212 1224
rect 300 1216 308 1224
rect 3948 1216 3956 1224
rect 1220 1206 1227 1214
rect 1227 1206 1228 1214
rect 1232 1206 1237 1214
rect 1237 1206 1239 1214
rect 1239 1206 1240 1214
rect 1244 1206 1247 1214
rect 1247 1206 1249 1214
rect 1249 1206 1252 1214
rect 1256 1206 1257 1214
rect 1257 1206 1259 1214
rect 1259 1206 1264 1214
rect 1268 1206 1269 1214
rect 1269 1206 1276 1214
rect 4228 1206 4235 1214
rect 4235 1206 4236 1214
rect 4240 1206 4245 1214
rect 4245 1206 4247 1214
rect 4247 1206 4248 1214
rect 4252 1206 4255 1214
rect 4255 1206 4257 1214
rect 4257 1206 4260 1214
rect 4264 1206 4265 1214
rect 4265 1206 4267 1214
rect 4267 1206 4272 1214
rect 4276 1206 4277 1214
rect 4277 1206 4284 1214
rect 460 1196 468 1204
rect 3532 1196 3540 1204
rect 1004 1176 1012 1184
rect 684 1156 692 1164
rect 1964 1136 1972 1144
rect 3724 1136 3732 1144
rect 44 1116 52 1124
rect 2476 1116 2484 1124
rect 4556 1116 4564 1124
rect 5036 1116 5044 1124
rect 4364 1096 4372 1104
rect 4780 1096 4788 1104
rect 588 1076 596 1084
rect 4460 1076 4468 1084
rect 4556 1076 4564 1084
rect 1484 1056 1492 1064
rect 2124 1056 2132 1064
rect 3628 1056 3636 1064
rect 4076 1056 4084 1064
rect 4524 1056 4532 1064
rect 2252 1036 2260 1044
rect 1452 1016 1460 1024
rect 3692 1016 3700 1024
rect 2724 1006 2731 1014
rect 2731 1006 2732 1014
rect 2736 1006 2741 1014
rect 2741 1006 2743 1014
rect 2743 1006 2744 1014
rect 2748 1006 2751 1014
rect 2751 1006 2753 1014
rect 2753 1006 2756 1014
rect 2760 1006 2761 1014
rect 2761 1006 2763 1014
rect 2763 1006 2768 1014
rect 2772 1006 2773 1014
rect 2773 1006 2780 1014
rect 3212 996 3220 1004
rect 4524 996 4532 1004
rect 4972 996 4980 1004
rect 428 976 436 984
rect 1836 976 1844 984
rect 2284 976 2292 984
rect 300 936 308 944
rect 524 936 532 944
rect 1932 936 1940 944
rect 4076 936 4084 944
rect 396 916 404 924
rect 876 916 884 924
rect 1004 916 1012 924
rect 1708 916 1716 924
rect 3500 916 3508 924
rect 3532 916 3540 924
rect 4492 916 4500 924
rect 4684 896 4692 904
rect 1612 876 1620 884
rect 3852 876 3860 884
rect 4428 836 4436 844
rect 300 816 308 824
rect 3532 816 3540 824
rect 4460 816 4468 824
rect 1220 806 1227 814
rect 1227 806 1228 814
rect 1232 806 1237 814
rect 1237 806 1239 814
rect 1239 806 1240 814
rect 1244 806 1247 814
rect 1247 806 1249 814
rect 1249 806 1252 814
rect 1256 806 1257 814
rect 1257 806 1259 814
rect 1259 806 1264 814
rect 1268 806 1269 814
rect 1269 806 1276 814
rect 4228 806 4235 814
rect 4235 806 4236 814
rect 4240 806 4245 814
rect 4245 806 4247 814
rect 4247 806 4248 814
rect 4252 806 4255 814
rect 4255 806 4257 814
rect 4257 806 4260 814
rect 4264 806 4265 814
rect 4265 806 4267 814
rect 4267 806 4272 814
rect 4276 806 4277 814
rect 4277 806 4284 814
rect 3276 776 3284 784
rect 4972 756 4980 764
rect 2284 736 2292 744
rect 4716 736 4724 744
rect 588 716 596 724
rect 5036 716 5044 724
rect 1164 696 1172 704
rect 5004 696 5012 704
rect 5100 696 5108 704
rect 780 676 788 684
rect 1484 616 1492 624
rect 2724 606 2731 614
rect 2731 606 2732 614
rect 2736 606 2741 614
rect 2741 606 2743 614
rect 2743 606 2744 614
rect 2748 606 2751 614
rect 2751 606 2753 614
rect 2753 606 2756 614
rect 2760 606 2761 614
rect 2761 606 2763 614
rect 2763 606 2768 614
rect 2772 606 2773 614
rect 2773 606 2780 614
rect 556 596 564 604
rect 3852 596 3860 604
rect 4684 616 4692 624
rect 1452 556 1460 564
rect 3532 556 3540 564
rect 4332 556 4340 564
rect 460 536 468 544
rect 2476 536 2484 544
rect 3084 536 3092 544
rect 3692 536 3700 544
rect 4076 536 4084 544
rect 1612 516 1620 524
rect 3628 516 3636 524
rect 4428 516 4436 524
rect 1484 496 1492 504
rect 4332 456 4340 464
rect 5036 456 5044 464
rect 5068 456 5076 464
rect 4972 436 4980 444
rect 4684 416 4692 424
rect 1220 406 1227 414
rect 1227 406 1228 414
rect 1232 406 1237 414
rect 1237 406 1239 414
rect 1239 406 1240 414
rect 1244 406 1247 414
rect 1247 406 1249 414
rect 1249 406 1252 414
rect 1256 406 1257 414
rect 1257 406 1259 414
rect 1259 406 1264 414
rect 1268 406 1269 414
rect 1269 406 1276 414
rect 4228 406 4235 414
rect 4235 406 4236 414
rect 4240 406 4245 414
rect 4245 406 4247 414
rect 4247 406 4248 414
rect 4252 406 4255 414
rect 4255 406 4257 414
rect 4257 406 4260 414
rect 4264 406 4265 414
rect 4265 406 4267 414
rect 4267 406 4272 414
rect 4276 406 4277 414
rect 4277 406 4284 414
rect 204 376 212 384
rect 5196 376 5204 384
rect 5324 376 5332 384
rect 5420 336 5428 344
rect 4876 316 4884 324
rect 5228 316 5236 324
rect 556 276 564 284
rect 3852 276 3860 284
rect 4716 236 4724 244
rect 4972 236 4980 244
rect 5004 236 5012 244
rect 4332 216 4340 224
rect 5036 216 5044 224
rect 2724 206 2731 214
rect 2731 206 2732 214
rect 2736 206 2741 214
rect 2741 206 2743 214
rect 2743 206 2744 214
rect 2748 206 2751 214
rect 2751 206 2753 214
rect 2753 206 2756 214
rect 2760 206 2761 214
rect 2761 206 2763 214
rect 2763 206 2768 214
rect 2772 206 2773 214
rect 2773 206 2780 214
rect 204 136 212 144
rect 3084 136 3092 144
rect 5452 116 5460 124
rect 3212 16 3220 24
rect 3500 16 3508 24
rect 4524 16 4532 24
rect 1220 6 1227 14
rect 1227 6 1228 14
rect 1232 6 1237 14
rect 1237 6 1239 14
rect 1239 6 1240 14
rect 1244 6 1247 14
rect 1247 6 1249 14
rect 1249 6 1252 14
rect 1256 6 1257 14
rect 1257 6 1259 14
rect 1259 6 1264 14
rect 1268 6 1269 14
rect 1269 6 1276 14
rect 4228 6 4235 14
rect 4235 6 4236 14
rect 4240 6 4245 14
rect 4245 6 4247 14
rect 4247 6 4248 14
rect 4252 6 4255 14
rect 4255 6 4257 14
rect 4257 6 4260 14
rect 4264 6 4265 14
rect 4265 6 4267 14
rect 4267 6 4272 14
rect 4276 6 4277 14
rect 4277 6 4284 14
<< metal4 >>
rect 2090 3824 2102 3826
rect 2090 3816 2092 3824
rect 2100 3816 2102 3824
rect 266 3744 278 3746
rect 266 3736 268 3744
rect 276 3736 278 3744
rect 266 3224 278 3736
rect 266 3216 268 3224
rect 276 3216 278 3224
rect 266 3214 278 3216
rect 714 3644 726 3646
rect 714 3636 716 3644
rect 724 3636 726 3644
rect 554 3164 566 3166
rect 554 3156 556 3164
rect 564 3156 566 3164
rect 330 3064 342 3066
rect 330 3056 332 3064
rect 340 3056 342 3064
rect 138 2964 150 2966
rect 138 2956 140 2964
rect 148 2956 150 2964
rect 138 2524 150 2956
rect 234 2784 246 2786
rect 234 2776 236 2784
rect 244 2776 246 2784
rect 234 2584 246 2776
rect 298 2724 310 2726
rect 298 2716 300 2724
rect 308 2716 310 2724
rect 298 2684 310 2716
rect 298 2676 300 2684
rect 308 2676 310 2684
rect 298 2674 310 2676
rect 234 2576 236 2584
rect 244 2576 246 2584
rect 234 2574 246 2576
rect 330 2564 342 3056
rect 458 3044 470 3046
rect 458 3036 460 3044
rect 468 3036 470 3044
rect 330 2556 332 2564
rect 340 2556 342 2564
rect 330 2554 342 2556
rect 394 2864 406 2866
rect 394 2856 396 2864
rect 404 2856 406 2864
rect 394 2704 406 2856
rect 394 2696 396 2704
rect 404 2696 406 2704
rect 138 2516 140 2524
rect 148 2516 150 2524
rect 138 2514 150 2516
rect 202 2464 214 2466
rect 202 2456 204 2464
rect 212 2456 214 2464
rect 202 2264 214 2456
rect 202 2256 204 2264
rect 212 2256 214 2264
rect 202 2254 214 2256
rect 298 2464 310 2466
rect 298 2456 300 2464
rect 308 2456 310 2464
rect 234 2064 246 2066
rect 234 2056 236 2064
rect 244 2056 246 2064
rect 42 1524 54 1526
rect 42 1516 44 1524
rect 52 1516 54 1524
rect 42 1124 54 1516
rect 202 1464 214 1466
rect 202 1456 204 1464
rect 212 1456 214 1464
rect 202 1224 214 1456
rect 234 1404 246 2056
rect 298 1864 310 2456
rect 330 2264 342 2266
rect 330 2256 332 2264
rect 340 2256 342 2264
rect 330 1944 342 2256
rect 394 2124 406 2696
rect 458 2664 470 3036
rect 458 2656 460 2664
rect 468 2656 470 2664
rect 458 2654 470 2656
rect 522 3004 534 3006
rect 522 2996 524 3004
rect 532 2996 534 3004
rect 394 2116 396 2124
rect 404 2116 406 2124
rect 394 2114 406 2116
rect 458 2564 470 2566
rect 458 2556 460 2564
rect 468 2556 470 2564
rect 458 2304 470 2556
rect 522 2504 534 2996
rect 554 2664 566 3156
rect 554 2656 556 2664
rect 564 2656 566 2664
rect 554 2654 566 2656
rect 682 3044 694 3046
rect 682 3036 684 3044
rect 692 3036 694 3044
rect 522 2496 524 2504
rect 532 2496 534 2504
rect 522 2494 534 2496
rect 618 2504 630 2506
rect 618 2496 620 2504
rect 628 2496 630 2504
rect 458 2296 460 2304
rect 468 2296 470 2304
rect 330 1936 332 1944
rect 340 1936 342 1944
rect 330 1934 342 1936
rect 426 2084 438 2086
rect 426 2076 428 2084
rect 436 2076 438 2084
rect 298 1856 300 1864
rect 308 1856 310 1864
rect 298 1854 310 1856
rect 234 1396 236 1404
rect 244 1396 246 1404
rect 234 1394 246 1396
rect 266 1824 278 1826
rect 266 1816 268 1824
rect 276 1816 278 1824
rect 266 1264 278 1816
rect 426 1684 438 2076
rect 458 1944 470 2296
rect 618 2284 630 2496
rect 682 2504 694 3036
rect 714 3044 726 3636
rect 1216 3614 1280 3816
rect 1216 3606 1220 3614
rect 1228 3606 1232 3614
rect 1240 3606 1244 3614
rect 1252 3606 1256 3614
rect 1264 3606 1268 3614
rect 1276 3606 1280 3614
rect 714 3036 716 3044
rect 724 3036 726 3044
rect 714 2664 726 3036
rect 746 3444 758 3446
rect 746 3436 748 3444
rect 756 3436 758 3444
rect 746 2964 758 3436
rect 810 3404 822 3406
rect 810 3396 812 3404
rect 820 3396 822 3404
rect 746 2956 748 2964
rect 756 2956 758 2964
rect 746 2954 758 2956
rect 778 3084 790 3086
rect 778 3076 780 3084
rect 788 3076 790 3084
rect 714 2656 716 2664
rect 724 2656 726 2664
rect 714 2654 726 2656
rect 746 2844 758 2846
rect 746 2836 748 2844
rect 756 2836 758 2844
rect 746 2664 758 2836
rect 746 2656 748 2664
rect 756 2656 758 2664
rect 746 2654 758 2656
rect 682 2496 684 2504
rect 692 2496 694 2504
rect 682 2494 694 2496
rect 618 2276 620 2284
rect 628 2276 630 2284
rect 618 2274 630 2276
rect 682 2084 694 2086
rect 682 2076 684 2084
rect 692 2076 694 2084
rect 458 1936 460 1944
rect 468 1936 470 1944
rect 458 1934 470 1936
rect 490 1984 502 1986
rect 490 1976 492 1984
rect 500 1976 502 1984
rect 426 1676 428 1684
rect 436 1676 438 1684
rect 426 1674 438 1676
rect 266 1256 268 1264
rect 276 1256 278 1264
rect 266 1254 278 1256
rect 298 1664 310 1666
rect 298 1656 300 1664
rect 308 1656 310 1664
rect 202 1216 204 1224
rect 212 1216 214 1224
rect 202 1214 214 1216
rect 298 1224 310 1656
rect 490 1604 502 1976
rect 490 1596 492 1604
rect 500 1596 502 1604
rect 490 1594 502 1596
rect 522 1844 534 1846
rect 522 1836 524 1844
rect 532 1836 534 1844
rect 426 1544 438 1546
rect 426 1536 428 1544
rect 436 1536 438 1544
rect 298 1216 300 1224
rect 308 1216 310 1224
rect 298 1214 310 1216
rect 394 1484 406 1486
rect 394 1476 396 1484
rect 404 1476 406 1484
rect 42 1116 44 1124
rect 52 1116 54 1124
rect 42 1114 54 1116
rect 298 944 310 946
rect 298 936 300 944
rect 308 936 310 944
rect 298 824 310 936
rect 394 924 406 1476
rect 426 984 438 1536
rect 426 976 428 984
rect 436 976 438 984
rect 426 974 438 976
rect 458 1204 470 1206
rect 458 1196 460 1204
rect 468 1196 470 1204
rect 394 916 396 924
rect 404 916 406 924
rect 394 914 406 916
rect 298 816 300 824
rect 308 816 310 824
rect 298 814 310 816
rect 458 544 470 1196
rect 522 944 534 1836
rect 682 1164 694 2076
rect 682 1156 684 1164
rect 692 1156 694 1164
rect 682 1154 694 1156
rect 522 936 524 944
rect 532 936 534 944
rect 522 934 534 936
rect 586 1084 598 1086
rect 586 1076 588 1084
rect 596 1076 598 1084
rect 586 724 598 1076
rect 586 716 588 724
rect 596 716 598 724
rect 586 714 598 716
rect 778 684 790 3076
rect 810 1904 822 3396
rect 1216 3214 1280 3606
rect 2090 3324 2102 3816
rect 2720 3814 2784 3816
rect 2720 3806 2724 3814
rect 2732 3806 2736 3814
rect 2744 3806 2748 3814
rect 2756 3806 2760 3814
rect 2768 3806 2772 3814
rect 2780 3806 2784 3814
rect 2090 3316 2092 3324
rect 2100 3316 2102 3324
rect 1216 3206 1220 3214
rect 1228 3206 1232 3214
rect 1240 3206 1244 3214
rect 1252 3206 1256 3214
rect 1264 3206 1268 3214
rect 1276 3206 1280 3214
rect 1098 2864 1110 2866
rect 1098 2856 1100 2864
rect 1108 2856 1110 2864
rect 810 1896 812 1904
rect 820 1896 822 1904
rect 810 1544 822 1896
rect 938 2004 950 2006
rect 938 1996 940 2004
rect 948 1996 950 2004
rect 938 1744 950 1996
rect 938 1736 940 1744
rect 948 1736 950 1744
rect 938 1734 950 1736
rect 1002 2004 1014 2006
rect 1002 1996 1004 2004
rect 1012 1996 1014 2004
rect 810 1536 812 1544
rect 820 1536 822 1544
rect 810 1534 822 1536
rect 874 1684 886 1686
rect 874 1676 876 1684
rect 884 1676 886 1684
rect 874 924 886 1676
rect 1002 1404 1014 1996
rect 1098 1984 1110 2856
rect 1098 1976 1100 1984
rect 1108 1976 1110 1984
rect 1098 1974 1110 1976
rect 1216 2814 1280 3206
rect 1802 3304 1814 3306
rect 1802 3296 1804 3304
rect 1812 3296 1814 3304
rect 1770 3064 1782 3066
rect 1770 3056 1772 3064
rect 1780 3056 1782 3064
rect 1216 2806 1220 2814
rect 1228 2806 1232 2814
rect 1240 2806 1244 2814
rect 1252 2806 1256 2814
rect 1264 2806 1268 2814
rect 1276 2806 1280 2814
rect 1216 2414 1280 2806
rect 1322 3004 1334 3006
rect 1322 2996 1324 3004
rect 1332 2996 1334 3004
rect 1322 2684 1334 2996
rect 1578 2784 1590 2786
rect 1578 2776 1580 2784
rect 1588 2776 1590 2784
rect 1322 2676 1324 2684
rect 1332 2676 1334 2684
rect 1322 2674 1334 2676
rect 1354 2704 1366 2706
rect 1354 2696 1356 2704
rect 1364 2696 1366 2704
rect 1216 2406 1220 2414
rect 1228 2406 1232 2414
rect 1240 2406 1244 2414
rect 1252 2406 1256 2414
rect 1264 2406 1268 2414
rect 1276 2406 1280 2414
rect 1216 2014 1280 2406
rect 1216 2006 1220 2014
rect 1228 2006 1232 2014
rect 1240 2006 1244 2014
rect 1252 2006 1256 2014
rect 1264 2006 1268 2014
rect 1276 2006 1280 2014
rect 1216 1614 1280 2006
rect 1322 2284 1334 2286
rect 1322 2276 1324 2284
rect 1332 2276 1334 2284
rect 1322 1884 1334 2276
rect 1354 2184 1366 2696
rect 1418 2704 1430 2706
rect 1418 2696 1420 2704
rect 1428 2696 1430 2704
rect 1418 2646 1430 2696
rect 1402 2644 1430 2646
rect 1402 2636 1404 2644
rect 1412 2636 1430 2644
rect 1402 2634 1430 2636
rect 1546 2684 1558 2686
rect 1546 2676 1548 2684
rect 1556 2676 1558 2684
rect 1354 2176 1356 2184
rect 1364 2176 1366 2184
rect 1354 2174 1366 2176
rect 1450 2624 1462 2626
rect 1450 2616 1452 2624
rect 1460 2616 1462 2624
rect 1322 1876 1324 1884
rect 1332 1876 1334 1884
rect 1322 1874 1334 1876
rect 1216 1606 1220 1614
rect 1228 1606 1232 1614
rect 1240 1606 1244 1614
rect 1252 1606 1256 1614
rect 1264 1606 1268 1614
rect 1276 1606 1280 1614
rect 1002 1396 1004 1404
rect 1012 1396 1014 1404
rect 1002 1394 1014 1396
rect 1162 1464 1174 1466
rect 1162 1456 1164 1464
rect 1172 1456 1174 1464
rect 874 916 876 924
rect 884 916 886 924
rect 874 914 886 916
rect 1002 1184 1014 1186
rect 1002 1176 1004 1184
rect 1012 1176 1014 1184
rect 1002 924 1014 1176
rect 1002 916 1004 924
rect 1012 916 1014 924
rect 1002 914 1014 916
rect 1162 704 1174 1456
rect 1162 696 1164 704
rect 1172 696 1174 704
rect 1162 694 1174 696
rect 1216 1214 1280 1606
rect 1450 1364 1462 2616
rect 1546 2424 1558 2676
rect 1578 2544 1590 2776
rect 1738 2764 1750 2766
rect 1738 2756 1740 2764
rect 1748 2756 1750 2764
rect 1578 2536 1580 2544
rect 1588 2536 1590 2544
rect 1578 2534 1590 2536
rect 1674 2604 1686 2606
rect 1674 2596 1676 2604
rect 1684 2596 1686 2604
rect 1546 2416 1548 2424
rect 1556 2416 1558 2424
rect 1546 2414 1558 2416
rect 1674 2324 1686 2596
rect 1738 2604 1750 2756
rect 1738 2596 1740 2604
rect 1748 2596 1750 2604
rect 1738 2594 1750 2596
rect 1770 2684 1782 3056
rect 1802 3004 1814 3296
rect 1802 2996 1804 3004
rect 1812 2996 1814 3004
rect 1802 2994 1814 2996
rect 1770 2676 1772 2684
rect 1780 2676 1782 2684
rect 1674 2316 1676 2324
rect 1684 2316 1686 2324
rect 1674 2314 1686 2316
rect 1706 2404 1718 2406
rect 1706 2396 1708 2404
rect 1716 2396 1718 2404
rect 1450 1356 1452 1364
rect 1460 1356 1462 1364
rect 1450 1354 1462 1356
rect 1642 2244 1654 2246
rect 1642 2236 1644 2244
rect 1652 2236 1654 2244
rect 1642 1284 1654 2236
rect 1642 1276 1644 1284
rect 1652 1276 1654 1284
rect 1642 1274 1654 1276
rect 1216 1206 1220 1214
rect 1228 1206 1232 1214
rect 1240 1206 1244 1214
rect 1252 1206 1256 1214
rect 1264 1206 1268 1214
rect 1276 1206 1280 1214
rect 1216 814 1280 1206
rect 1482 1064 1494 1066
rect 1482 1056 1484 1064
rect 1492 1056 1494 1064
rect 1216 806 1220 814
rect 1228 806 1232 814
rect 1240 806 1244 814
rect 1252 806 1256 814
rect 1264 806 1268 814
rect 1276 806 1280 814
rect 778 676 780 684
rect 788 676 790 684
rect 778 674 790 676
rect 458 536 460 544
rect 468 536 470 544
rect 458 534 470 536
rect 554 604 566 606
rect 554 596 556 604
rect 564 596 566 604
rect 202 384 214 386
rect 202 376 204 384
rect 212 376 214 384
rect 202 144 214 376
rect 554 284 566 596
rect 554 276 556 284
rect 564 276 566 284
rect 554 274 566 276
rect 1216 414 1280 806
rect 1450 1024 1462 1026
rect 1450 1016 1452 1024
rect 1460 1016 1462 1024
rect 1450 564 1462 1016
rect 1450 556 1452 564
rect 1460 556 1462 564
rect 1450 554 1462 556
rect 1482 624 1494 1056
rect 1706 924 1718 2396
rect 1770 2324 1782 2676
rect 1898 2904 1910 2906
rect 1898 2896 1900 2904
rect 1908 2896 1910 2904
rect 1770 2316 1772 2324
rect 1780 2316 1782 2324
rect 1770 2314 1782 2316
rect 1834 2364 1846 2366
rect 1834 2356 1836 2364
rect 1844 2356 1846 2364
rect 1834 984 1846 2356
rect 1898 1284 1910 2896
rect 2058 2844 2070 2846
rect 2058 2836 2060 2844
rect 2068 2836 2070 2844
rect 2058 2384 2070 2836
rect 2090 2404 2102 3316
rect 2378 3444 2390 3446
rect 2378 3436 2380 3444
rect 2388 3436 2390 3444
rect 2378 3224 2390 3436
rect 2378 3216 2380 3224
rect 2388 3216 2390 3224
rect 2378 3214 2390 3216
rect 2720 3414 2784 3806
rect 3594 3744 3606 3746
rect 3594 3736 3596 3744
rect 3604 3736 3606 3744
rect 3242 3644 3254 3646
rect 3242 3636 3244 3644
rect 3252 3636 3254 3644
rect 2720 3406 2724 3414
rect 2732 3406 2736 3414
rect 2744 3406 2748 3414
rect 2756 3406 2760 3414
rect 2768 3406 2772 3414
rect 2780 3406 2784 3414
rect 2720 3014 2784 3406
rect 2858 3464 2870 3466
rect 2858 3456 2860 3464
rect 2868 3456 2870 3464
rect 2858 3244 2870 3456
rect 3242 3384 3254 3636
rect 3242 3376 3244 3384
rect 3252 3376 3254 3384
rect 3242 3374 3254 3376
rect 2858 3236 2860 3244
rect 2868 3236 2870 3244
rect 2858 3234 2870 3236
rect 3370 3324 3382 3326
rect 3370 3316 3372 3324
rect 3380 3316 3382 3324
rect 2720 3006 2724 3014
rect 2732 3006 2736 3014
rect 2744 3006 2748 3014
rect 2756 3006 2760 3014
rect 2768 3006 2772 3014
rect 2780 3006 2784 3014
rect 2410 2924 2422 2926
rect 2410 2916 2412 2924
rect 2420 2916 2422 2924
rect 2346 2904 2358 2906
rect 2346 2896 2348 2904
rect 2356 2896 2358 2904
rect 2250 2804 2262 2806
rect 2250 2796 2252 2804
rect 2260 2796 2262 2804
rect 2090 2396 2092 2404
rect 2100 2396 2102 2404
rect 2090 2394 2102 2396
rect 2154 2764 2166 2766
rect 2154 2756 2156 2764
rect 2164 2756 2166 2764
rect 2058 2376 2060 2384
rect 2068 2376 2070 2384
rect 2058 2374 2070 2376
rect 2122 1824 2134 1826
rect 2122 1816 2124 1824
rect 2132 1816 2134 1824
rect 1962 1484 1974 1486
rect 1962 1476 1964 1484
rect 1972 1476 1974 1484
rect 1898 1276 1900 1284
rect 1908 1276 1910 1284
rect 1898 1274 1910 1276
rect 1930 1304 1942 1306
rect 1930 1296 1932 1304
rect 1940 1296 1942 1304
rect 1834 976 1836 984
rect 1844 976 1846 984
rect 1834 974 1846 976
rect 1930 944 1942 1296
rect 1962 1144 1974 1476
rect 1962 1136 1964 1144
rect 1972 1136 1974 1144
rect 1962 1134 1974 1136
rect 2122 1064 2134 1816
rect 2154 1524 2166 2756
rect 2250 2064 2262 2796
rect 2250 2056 2252 2064
rect 2260 2056 2262 2064
rect 2250 2054 2262 2056
rect 2314 2064 2326 2066
rect 2314 2056 2316 2064
rect 2324 2056 2326 2064
rect 2154 1516 2156 1524
rect 2164 1516 2166 1524
rect 2154 1514 2166 1516
rect 2250 1944 2262 1946
rect 2250 1936 2252 1944
rect 2260 1936 2262 1944
rect 2122 1056 2124 1064
rect 2132 1056 2134 1064
rect 2122 1054 2134 1056
rect 2250 1044 2262 1936
rect 2282 1944 2294 1946
rect 2282 1936 2284 1944
rect 2292 1936 2294 1944
rect 2282 1764 2294 1936
rect 2282 1756 2284 1764
rect 2292 1756 2294 1764
rect 2282 1754 2294 1756
rect 2314 1344 2326 2056
rect 2346 2064 2358 2896
rect 2410 2584 2422 2916
rect 2410 2576 2412 2584
rect 2420 2576 2422 2584
rect 2410 2574 2422 2576
rect 2474 2744 2486 2746
rect 2474 2736 2476 2744
rect 2484 2736 2486 2744
rect 2346 2056 2348 2064
rect 2356 2056 2358 2064
rect 2346 2054 2358 2056
rect 2474 1764 2486 2736
rect 2720 2614 2784 3006
rect 3338 2984 3350 2986
rect 3338 2976 3340 2984
rect 3348 2976 3350 2984
rect 3210 2924 3222 2926
rect 3210 2916 3212 2924
rect 3220 2916 3222 2924
rect 2720 2606 2724 2614
rect 2732 2606 2736 2614
rect 2744 2606 2748 2614
rect 2756 2606 2760 2614
rect 2768 2606 2772 2614
rect 2780 2606 2784 2614
rect 2602 2284 2614 2286
rect 2602 2276 2604 2284
rect 2612 2276 2614 2284
rect 2474 1756 2476 1764
rect 2484 1756 2486 1764
rect 2474 1754 2486 1756
rect 2506 2044 2518 2046
rect 2506 2036 2508 2044
rect 2516 2036 2518 2044
rect 2410 1584 2422 1586
rect 2410 1576 2412 1584
rect 2420 1576 2422 1584
rect 2410 1364 2422 1576
rect 2506 1404 2518 2036
rect 2602 2024 2614 2276
rect 2602 2016 2604 2024
rect 2612 2016 2614 2024
rect 2602 2014 2614 2016
rect 2720 2214 2784 2606
rect 2826 2804 2838 2806
rect 2826 2796 2828 2804
rect 2836 2796 2838 2804
rect 2826 2504 2838 2796
rect 2954 2764 2966 2766
rect 2954 2756 2956 2764
rect 2964 2756 2966 2764
rect 2890 2684 2902 2686
rect 2890 2676 2892 2684
rect 2900 2676 2902 2684
rect 2890 2564 2902 2676
rect 2890 2556 2892 2564
rect 2900 2556 2902 2564
rect 2890 2554 2902 2556
rect 2826 2496 2828 2504
rect 2836 2496 2838 2504
rect 2826 2494 2838 2496
rect 2720 2206 2724 2214
rect 2732 2206 2736 2214
rect 2744 2206 2748 2214
rect 2756 2206 2760 2214
rect 2768 2206 2772 2214
rect 2780 2206 2784 2214
rect 2506 1396 2508 1404
rect 2516 1396 2518 1404
rect 2506 1394 2518 1396
rect 2720 1814 2784 2206
rect 2720 1806 2724 1814
rect 2732 1806 2736 1814
rect 2744 1806 2748 1814
rect 2756 1806 2760 1814
rect 2768 1806 2772 1814
rect 2780 1806 2784 1814
rect 2720 1414 2784 1806
rect 2826 1924 2838 1926
rect 2826 1916 2828 1924
rect 2836 1916 2838 1924
rect 2826 1744 2838 1916
rect 2826 1736 2828 1744
rect 2836 1736 2838 1744
rect 2826 1734 2838 1736
rect 2720 1406 2724 1414
rect 2732 1406 2736 1414
rect 2744 1406 2748 1414
rect 2756 1406 2760 1414
rect 2768 1406 2772 1414
rect 2780 1406 2784 1414
rect 2410 1356 2412 1364
rect 2420 1356 2422 1364
rect 2410 1354 2422 1356
rect 2314 1336 2316 1344
rect 2324 1336 2326 1344
rect 2314 1284 2326 1336
rect 2314 1276 2316 1284
rect 2324 1276 2326 1284
rect 2314 1274 2326 1276
rect 2250 1036 2252 1044
rect 2260 1036 2262 1044
rect 2250 1034 2262 1036
rect 2474 1124 2486 1126
rect 2474 1116 2476 1124
rect 2484 1116 2486 1124
rect 1930 936 1932 944
rect 1940 936 1942 944
rect 1930 934 1942 936
rect 2282 984 2294 986
rect 2282 976 2284 984
rect 2292 976 2294 984
rect 1706 916 1708 924
rect 1716 916 1718 924
rect 1706 914 1718 916
rect 1482 616 1484 624
rect 1492 616 1494 624
rect 1482 504 1494 616
rect 1610 884 1622 886
rect 1610 876 1612 884
rect 1620 876 1622 884
rect 1610 524 1622 876
rect 2282 744 2294 976
rect 2282 736 2284 744
rect 2292 736 2294 744
rect 2282 734 2294 736
rect 2474 544 2486 1116
rect 2474 536 2476 544
rect 2484 536 2486 544
rect 2474 534 2486 536
rect 2720 1014 2784 1406
rect 2954 1264 2966 2756
rect 3018 2664 3030 2666
rect 3018 2656 3020 2664
rect 3028 2656 3030 2664
rect 3018 1744 3030 2656
rect 3018 1736 3020 1744
rect 3028 1736 3030 1744
rect 3018 1734 3030 1736
rect 3178 2464 3190 2466
rect 3178 2456 3180 2464
rect 3188 2456 3190 2464
rect 2954 1256 2956 1264
rect 2964 1256 2966 1264
rect 2954 1254 2966 1256
rect 3082 1704 3094 1706
rect 3082 1696 3084 1704
rect 3092 1696 3094 1704
rect 2720 1006 2724 1014
rect 2732 1006 2736 1014
rect 2744 1006 2748 1014
rect 2756 1006 2760 1014
rect 2768 1006 2772 1014
rect 2780 1006 2784 1014
rect 2720 614 2784 1006
rect 2720 606 2724 614
rect 2732 606 2736 614
rect 2744 606 2748 614
rect 2756 606 2760 614
rect 2768 606 2772 614
rect 2780 606 2784 614
rect 1610 516 1612 524
rect 1620 516 1622 524
rect 1610 514 1622 516
rect 1482 496 1484 504
rect 1492 496 1494 504
rect 1482 494 1494 496
rect 1216 406 1220 414
rect 1228 406 1232 414
rect 1240 406 1244 414
rect 1252 406 1256 414
rect 1264 406 1268 414
rect 1276 406 1280 414
rect 202 136 204 144
rect 212 136 214 144
rect 202 134 214 136
rect 1216 14 1280 406
rect 1216 6 1220 14
rect 1228 6 1232 14
rect 1240 6 1244 14
rect 1252 6 1256 14
rect 1264 6 1268 14
rect 1276 6 1280 14
rect 1216 -10 1280 6
rect 2720 214 2784 606
rect 2720 206 2724 214
rect 2732 206 2736 214
rect 2744 206 2748 214
rect 2756 206 2760 214
rect 2768 206 2772 214
rect 2780 206 2784 214
rect 2720 -10 2784 206
rect 3082 544 3094 1696
rect 3178 1244 3190 2456
rect 3210 2464 3222 2916
rect 3210 2456 3212 2464
rect 3220 2456 3222 2464
rect 3210 2454 3222 2456
rect 3178 1236 3180 1244
rect 3188 1236 3190 1244
rect 3178 1234 3190 1236
rect 3274 1684 3286 1686
rect 3274 1676 3276 1684
rect 3284 1676 3286 1684
rect 3082 536 3084 544
rect 3092 536 3094 544
rect 3082 144 3094 536
rect 3082 136 3084 144
rect 3092 136 3094 144
rect 3082 134 3094 136
rect 3210 1004 3222 1006
rect 3210 996 3212 1004
rect 3220 996 3222 1004
rect 3210 24 3222 996
rect 3274 784 3286 1676
rect 3338 1664 3350 2976
rect 3370 2924 3382 3316
rect 3594 3284 3606 3736
rect 3914 3724 3926 3726
rect 3914 3716 3916 3724
rect 3924 3716 3926 3724
rect 3594 3276 3596 3284
rect 3604 3276 3606 3284
rect 3594 3274 3606 3276
rect 3658 3684 3670 3686
rect 3658 3676 3660 3684
rect 3668 3676 3670 3684
rect 3658 3404 3670 3676
rect 3658 3396 3660 3404
rect 3668 3396 3670 3404
rect 3658 3044 3670 3396
rect 3722 3504 3734 3506
rect 3722 3496 3724 3504
rect 3732 3496 3734 3504
rect 3722 3304 3734 3496
rect 3722 3296 3724 3304
rect 3732 3296 3734 3304
rect 3722 3294 3734 3296
rect 3658 3036 3660 3044
rect 3668 3036 3670 3044
rect 3658 3034 3670 3036
rect 3754 3224 3766 3226
rect 3754 3216 3756 3224
rect 3764 3216 3766 3224
rect 3754 3144 3766 3216
rect 3914 3224 3926 3716
rect 4224 3614 4288 3816
rect 4224 3606 4228 3614
rect 4236 3606 4240 3614
rect 4248 3606 4252 3614
rect 4260 3606 4264 3614
rect 4272 3606 4276 3614
rect 4284 3606 4288 3614
rect 3978 3584 3990 3586
rect 3978 3576 3980 3584
rect 3988 3576 3990 3584
rect 3978 3284 3990 3576
rect 4106 3504 4118 3506
rect 4106 3496 4108 3504
rect 4116 3496 4118 3504
rect 4106 3444 4118 3496
rect 4106 3436 4108 3444
rect 4116 3436 4118 3444
rect 4106 3434 4118 3436
rect 3978 3276 3980 3284
rect 3988 3276 3990 3284
rect 3978 3274 3990 3276
rect 4010 3344 4022 3346
rect 4010 3336 4012 3344
rect 4020 3336 4022 3344
rect 3914 3216 3916 3224
rect 3924 3216 3926 3224
rect 3914 3214 3926 3216
rect 3754 3136 3756 3144
rect 3764 3136 3766 3144
rect 3370 2916 3372 2924
rect 3380 2916 3382 2924
rect 3370 2914 3382 2916
rect 3466 2984 3478 2986
rect 3466 2976 3468 2984
rect 3476 2976 3478 2984
rect 3466 2484 3478 2976
rect 3754 2904 3766 3136
rect 3850 2964 3862 2966
rect 3850 2956 3852 2964
rect 3860 2956 3862 2964
rect 3850 2924 3862 2956
rect 3850 2916 3852 2924
rect 3860 2916 3862 2924
rect 3850 2914 3862 2916
rect 3754 2896 3756 2904
rect 3764 2896 3766 2904
rect 3754 2894 3766 2896
rect 4010 2904 4022 3336
rect 4074 3304 4086 3306
rect 4074 3296 4076 3304
rect 4084 3296 4086 3304
rect 4042 3284 4054 3286
rect 4042 3276 4044 3284
rect 4052 3276 4054 3284
rect 4042 3084 4054 3276
rect 4042 3076 4044 3084
rect 4052 3076 4054 3084
rect 4042 3074 4054 3076
rect 4010 2896 4012 2904
rect 4020 2896 4022 2904
rect 4010 2894 4022 2896
rect 4074 2904 4086 3296
rect 4074 2896 4076 2904
rect 4084 2896 4086 2904
rect 4074 2894 4086 2896
rect 4224 3214 4288 3606
rect 5258 3684 5270 3686
rect 5258 3676 5260 3684
rect 5268 3676 5270 3684
rect 4426 3584 4438 3586
rect 4426 3576 4428 3584
rect 4436 3576 4438 3584
rect 4426 3544 4438 3576
rect 4426 3536 4428 3544
rect 4436 3536 4438 3544
rect 4426 3534 4438 3536
rect 4490 3504 4502 3506
rect 4490 3496 4492 3504
rect 4500 3496 4502 3504
rect 4362 3344 4374 3346
rect 4362 3336 4364 3344
rect 4372 3336 4374 3344
rect 4362 3304 4374 3336
rect 4490 3324 4502 3496
rect 4650 3464 4662 3466
rect 4650 3456 4652 3464
rect 4660 3456 4662 3464
rect 4490 3316 4492 3324
rect 4500 3316 4502 3324
rect 4490 3314 4502 3316
rect 4586 3384 4598 3386
rect 4586 3376 4588 3384
rect 4596 3376 4598 3384
rect 4362 3296 4364 3304
rect 4372 3296 4374 3304
rect 4362 3294 4374 3296
rect 4224 3206 4228 3214
rect 4236 3206 4240 3214
rect 4248 3206 4252 3214
rect 4260 3206 4264 3214
rect 4272 3206 4276 3214
rect 4284 3206 4288 3214
rect 4224 2814 4288 3206
rect 4224 2806 4228 2814
rect 4236 2806 4240 2814
rect 4248 2806 4252 2814
rect 4260 2806 4264 2814
rect 4272 2806 4276 2814
rect 4284 2806 4288 2814
rect 3466 2476 3468 2484
rect 3476 2476 3478 2484
rect 3466 2474 3478 2476
rect 3530 2744 3542 2746
rect 3530 2736 3532 2744
rect 3540 2736 3542 2744
rect 3370 2204 3382 2206
rect 3370 2196 3372 2204
rect 3380 2196 3382 2204
rect 3370 2164 3382 2196
rect 3370 2156 3372 2164
rect 3380 2156 3382 2164
rect 3370 2154 3382 2156
rect 3498 2104 3510 2106
rect 3498 2096 3500 2104
rect 3508 2096 3510 2104
rect 3498 1784 3510 2096
rect 3530 1944 3542 2736
rect 4074 2724 4086 2726
rect 4074 2716 4076 2724
rect 4084 2716 4086 2724
rect 3818 2584 3830 2586
rect 3818 2576 3820 2584
rect 3828 2576 3830 2584
rect 3658 2484 3670 2486
rect 3658 2476 3660 2484
rect 3668 2476 3670 2484
rect 3530 1936 3532 1944
rect 3540 1936 3542 1944
rect 3530 1934 3542 1936
rect 3594 2404 3606 2406
rect 3594 2396 3596 2404
rect 3604 2396 3606 2404
rect 3498 1776 3500 1784
rect 3508 1776 3510 1784
rect 3498 1774 3510 1776
rect 3594 1784 3606 2396
rect 3658 2384 3670 2476
rect 3658 2376 3660 2384
rect 3668 2376 3670 2384
rect 3658 2374 3670 2376
rect 3754 2184 3766 2186
rect 3754 2176 3756 2184
rect 3764 2176 3766 2184
rect 3754 2104 3766 2176
rect 3754 2096 3756 2104
rect 3764 2096 3766 2104
rect 3754 2094 3766 2096
rect 3818 2084 3830 2576
rect 4074 2164 4086 2716
rect 4224 2414 4288 2806
rect 4224 2406 4228 2414
rect 4236 2406 4240 2414
rect 4248 2406 4252 2414
rect 4260 2406 4264 2414
rect 4272 2406 4276 2414
rect 4284 2406 4288 2414
rect 4074 2156 4076 2164
rect 4084 2156 4086 2164
rect 4074 2154 4086 2156
rect 4106 2164 4118 2166
rect 4106 2156 4108 2164
rect 4116 2156 4118 2164
rect 3818 2076 3820 2084
rect 3828 2076 3830 2084
rect 3818 2074 3830 2076
rect 3978 2124 3990 2126
rect 3978 2116 3980 2124
rect 3988 2116 3990 2124
rect 3946 2004 3958 2006
rect 3946 1996 3948 2004
rect 3956 1996 3958 2004
rect 3594 1776 3596 1784
rect 3604 1776 3606 1784
rect 3594 1774 3606 1776
rect 3754 1904 3766 1906
rect 3754 1896 3756 1904
rect 3764 1896 3766 1904
rect 3338 1656 3340 1664
rect 3348 1656 3350 1664
rect 3338 1654 3350 1656
rect 3722 1584 3734 1586
rect 3722 1576 3724 1584
rect 3732 1576 3734 1584
rect 3530 1204 3542 1206
rect 3530 1196 3532 1204
rect 3540 1196 3542 1204
rect 3274 776 3276 784
rect 3284 776 3286 784
rect 3274 774 3286 776
rect 3498 924 3510 926
rect 3498 916 3500 924
rect 3508 916 3510 924
rect 3210 16 3212 24
rect 3220 16 3222 24
rect 3210 14 3222 16
rect 3498 24 3510 916
rect 3530 924 3542 1196
rect 3722 1144 3734 1576
rect 3754 1464 3766 1896
rect 3754 1456 3756 1464
rect 3764 1456 3766 1464
rect 3754 1454 3766 1456
rect 3722 1136 3724 1144
rect 3732 1136 3734 1144
rect 3722 1134 3734 1136
rect 3850 1364 3862 1366
rect 3850 1356 3852 1364
rect 3860 1356 3862 1364
rect 3530 916 3532 924
rect 3540 916 3542 924
rect 3530 914 3542 916
rect 3626 1064 3638 1066
rect 3626 1056 3628 1064
rect 3636 1056 3638 1064
rect 3530 824 3542 826
rect 3530 816 3532 824
rect 3540 816 3542 824
rect 3530 564 3542 816
rect 3530 556 3532 564
rect 3540 556 3542 564
rect 3530 554 3542 556
rect 3626 524 3638 1056
rect 3690 1024 3702 1026
rect 3690 1016 3692 1024
rect 3700 1016 3702 1024
rect 3690 544 3702 1016
rect 3850 884 3862 1356
rect 3946 1344 3958 1996
rect 3978 1664 3990 2116
rect 4074 1864 4086 1866
rect 4074 1856 4076 1864
rect 4084 1856 4086 1864
rect 3978 1656 3980 1664
rect 3988 1656 3990 1664
rect 3978 1584 3990 1656
rect 3978 1576 3980 1584
rect 3988 1576 3990 1584
rect 3978 1574 3990 1576
rect 4010 1744 4022 1746
rect 4010 1736 4012 1744
rect 4020 1736 4022 1744
rect 4010 1484 4022 1736
rect 4010 1476 4012 1484
rect 4020 1476 4022 1484
rect 4010 1474 4022 1476
rect 4074 1704 4086 1856
rect 4074 1696 4076 1704
rect 4084 1696 4086 1704
rect 3946 1336 3948 1344
rect 3956 1336 3958 1344
rect 3946 1224 3958 1336
rect 3946 1216 3948 1224
rect 3956 1216 3958 1224
rect 3946 1214 3958 1216
rect 4074 1064 4086 1696
rect 4106 1304 4118 2156
rect 4138 2084 4150 2086
rect 4138 2076 4140 2084
rect 4148 2076 4150 2084
rect 4138 2024 4150 2076
rect 4138 2016 4140 2024
rect 4148 2016 4150 2024
rect 4138 2014 4150 2016
rect 4224 2014 4288 2406
rect 4426 2924 4438 2926
rect 4426 2916 4428 2924
rect 4436 2916 4438 2924
rect 4426 2484 4438 2916
rect 4426 2476 4428 2484
rect 4436 2476 4438 2484
rect 4426 2264 4438 2476
rect 4426 2256 4428 2264
rect 4436 2256 4438 2264
rect 4426 2254 4438 2256
rect 4458 2604 4470 2606
rect 4458 2596 4460 2604
rect 4468 2596 4470 2604
rect 4458 2164 4470 2596
rect 4458 2156 4460 2164
rect 4468 2156 4470 2164
rect 4458 2154 4470 2156
rect 4554 2584 4566 2586
rect 4554 2576 4556 2584
rect 4564 2576 4566 2584
rect 4554 2144 4566 2576
rect 4586 2284 4598 3376
rect 4586 2276 4588 2284
rect 4596 2276 4598 2284
rect 4586 2274 4598 2276
rect 4554 2136 4556 2144
rect 4564 2136 4566 2144
rect 4554 2134 4566 2136
rect 4586 2224 4598 2226
rect 4586 2216 4588 2224
rect 4596 2216 4598 2224
rect 4224 2006 4228 2014
rect 4236 2006 4240 2014
rect 4248 2006 4252 2014
rect 4260 2006 4264 2014
rect 4272 2006 4276 2014
rect 4284 2006 4288 2014
rect 4170 1804 4182 1806
rect 4170 1796 4172 1804
rect 4180 1796 4182 1804
rect 4170 1504 4182 1796
rect 4170 1496 4172 1504
rect 4180 1496 4182 1504
rect 4170 1494 4182 1496
rect 4224 1614 4288 2006
rect 4554 2064 4566 2066
rect 4554 2056 4556 2064
rect 4564 2056 4566 2064
rect 4224 1606 4228 1614
rect 4236 1606 4240 1614
rect 4248 1606 4252 1614
rect 4260 1606 4264 1614
rect 4272 1606 4276 1614
rect 4284 1606 4288 1614
rect 4106 1296 4108 1304
rect 4116 1296 4118 1304
rect 4106 1294 4118 1296
rect 4074 1056 4076 1064
rect 4084 1056 4086 1064
rect 4074 1054 4086 1056
rect 4224 1214 4288 1606
rect 4224 1206 4228 1214
rect 4236 1206 4240 1214
rect 4248 1206 4252 1214
rect 4260 1206 4264 1214
rect 4272 1206 4276 1214
rect 4284 1206 4288 1214
rect 3850 876 3852 884
rect 3860 876 3862 884
rect 3850 874 3862 876
rect 4074 944 4086 946
rect 4074 936 4076 944
rect 4084 936 4086 944
rect 3690 536 3692 544
rect 3700 536 3702 544
rect 3690 534 3702 536
rect 3850 604 3862 606
rect 3850 596 3852 604
rect 3860 596 3862 604
rect 3626 516 3628 524
rect 3636 516 3638 524
rect 3626 514 3638 516
rect 3850 284 3862 596
rect 4074 544 4086 936
rect 4074 536 4076 544
rect 4084 536 4086 544
rect 4074 534 4086 536
rect 4224 814 4288 1206
rect 4362 1944 4374 1946
rect 4362 1936 4364 1944
rect 4372 1936 4374 1944
rect 4362 1104 4374 1936
rect 4362 1096 4364 1104
rect 4372 1096 4374 1104
rect 4362 1094 4374 1096
rect 4490 1504 4502 1506
rect 4490 1496 4492 1504
rect 4500 1496 4502 1504
rect 4458 1084 4470 1086
rect 4458 1076 4460 1084
rect 4468 1076 4470 1084
rect 4224 806 4228 814
rect 4236 806 4240 814
rect 4248 806 4252 814
rect 4260 806 4264 814
rect 4272 806 4276 814
rect 4284 806 4288 814
rect 3850 276 3852 284
rect 3860 276 3862 284
rect 3850 274 3862 276
rect 4224 414 4288 806
rect 4426 844 4438 846
rect 4426 836 4428 844
rect 4436 836 4438 844
rect 4224 406 4228 414
rect 4236 406 4240 414
rect 4248 406 4252 414
rect 4260 406 4264 414
rect 4272 406 4276 414
rect 4284 406 4288 414
rect 3498 16 3500 24
rect 3508 16 3510 24
rect 3498 14 3510 16
rect 4224 14 4288 406
rect 4330 564 4342 566
rect 4330 556 4332 564
rect 4340 556 4342 564
rect 4330 464 4342 556
rect 4426 524 4438 836
rect 4458 824 4470 1076
rect 4490 924 4502 1496
rect 4554 1124 4566 2056
rect 4586 2044 4598 2216
rect 4650 2124 4662 3456
rect 5226 3444 5238 3446
rect 5226 3436 5228 3444
rect 5236 3436 5238 3444
rect 4682 3404 4694 3406
rect 4682 3396 4684 3404
rect 4692 3396 4694 3404
rect 4682 2624 4694 3396
rect 4746 3364 4758 3366
rect 4746 3356 4748 3364
rect 4756 3356 4758 3364
rect 4746 3184 4758 3356
rect 4746 3176 4748 3184
rect 4756 3176 4758 3184
rect 4746 3174 4758 3176
rect 5034 3044 5046 3046
rect 5034 3036 5036 3044
rect 5044 3036 5046 3044
rect 4938 3024 4950 3026
rect 4938 3016 4940 3024
rect 4948 3016 4950 3024
rect 4682 2616 4684 2624
rect 4692 2616 4694 2624
rect 4682 2614 4694 2616
rect 4778 2944 4790 2946
rect 4778 2936 4780 2944
rect 4788 2936 4790 2944
rect 4650 2116 4652 2124
rect 4660 2116 4662 2124
rect 4650 2114 4662 2116
rect 4714 2284 4726 2286
rect 4714 2276 4716 2284
rect 4724 2276 4726 2284
rect 4586 2036 4588 2044
rect 4596 2036 4598 2044
rect 4586 2034 4598 2036
rect 4618 2024 4630 2026
rect 4618 2016 4620 2024
rect 4628 2016 4630 2024
rect 4618 1464 4630 2016
rect 4650 1904 4662 1906
rect 4650 1896 4652 1904
rect 4660 1896 4662 1904
rect 4650 1604 4662 1896
rect 4650 1596 4652 1604
rect 4660 1596 4662 1604
rect 4650 1594 4662 1596
rect 4682 1804 4694 1806
rect 4682 1796 4684 1804
rect 4692 1796 4694 1804
rect 4618 1456 4620 1464
rect 4628 1456 4630 1464
rect 4618 1454 4630 1456
rect 4682 1504 4694 1796
rect 4714 1744 4726 2276
rect 4714 1736 4716 1744
rect 4724 1736 4726 1744
rect 4714 1734 4726 1736
rect 4746 2284 4758 2286
rect 4746 2276 4748 2284
rect 4756 2276 4758 2284
rect 4682 1496 4684 1504
rect 4692 1496 4694 1504
rect 4554 1116 4556 1124
rect 4564 1116 4566 1124
rect 4554 1084 4566 1116
rect 4554 1076 4556 1084
rect 4564 1076 4566 1084
rect 4554 1074 4566 1076
rect 4490 916 4492 924
rect 4500 916 4502 924
rect 4490 914 4502 916
rect 4522 1064 4534 1066
rect 4522 1056 4524 1064
rect 4532 1056 4534 1064
rect 4522 1004 4534 1056
rect 4522 996 4524 1004
rect 4532 996 4534 1004
rect 4458 816 4460 824
rect 4468 816 4470 824
rect 4458 814 4470 816
rect 4426 516 4428 524
rect 4436 516 4438 524
rect 4426 514 4438 516
rect 4330 456 4332 464
rect 4340 456 4342 464
rect 4330 224 4342 456
rect 4330 216 4332 224
rect 4340 216 4342 224
rect 4330 214 4342 216
rect 4522 24 4534 996
rect 4682 904 4694 1496
rect 4746 1424 4758 2276
rect 4778 1804 4790 2936
rect 4810 2584 4822 2586
rect 4810 2576 4812 2584
rect 4820 2576 4822 2584
rect 4810 1904 4822 2576
rect 4938 2564 4950 3016
rect 4938 2556 4940 2564
rect 4948 2556 4950 2564
rect 4938 2554 4950 2556
rect 5002 2924 5014 2926
rect 5002 2916 5004 2924
rect 5012 2916 5014 2924
rect 5002 2184 5014 2916
rect 5002 2176 5004 2184
rect 5012 2176 5014 2184
rect 5002 2174 5014 2176
rect 4810 1896 4812 1904
rect 4820 1896 4822 1904
rect 4810 1894 4822 1896
rect 4874 2124 4886 2126
rect 4874 2116 4876 2124
rect 4884 2116 4886 2124
rect 4778 1796 4780 1804
rect 4788 1796 4790 1804
rect 4778 1794 4790 1796
rect 4810 1804 4822 1806
rect 4810 1796 4812 1804
rect 4820 1796 4822 1804
rect 4746 1416 4748 1424
rect 4756 1416 4758 1424
rect 4746 1414 4758 1416
rect 4778 1744 4790 1746
rect 4778 1736 4780 1744
rect 4788 1736 4790 1744
rect 4778 1104 4790 1736
rect 4810 1404 4822 1796
rect 4810 1396 4812 1404
rect 4820 1396 4822 1404
rect 4810 1394 4822 1396
rect 4778 1096 4780 1104
rect 4788 1096 4790 1104
rect 4778 1094 4790 1096
rect 4682 896 4684 904
rect 4692 896 4694 904
rect 4682 894 4694 896
rect 4714 744 4726 746
rect 4714 736 4716 744
rect 4724 736 4726 744
rect 4682 624 4694 626
rect 4682 616 4684 624
rect 4692 616 4694 624
rect 4682 424 4694 616
rect 4682 416 4684 424
rect 4692 416 4694 424
rect 4682 414 4694 416
rect 4714 244 4726 736
rect 4874 324 4886 2116
rect 5002 2004 5014 2006
rect 5002 1996 5004 2004
rect 5012 1996 5014 2004
rect 4970 1764 4982 1766
rect 4970 1756 4972 1764
rect 4980 1756 4982 1764
rect 4970 1664 4982 1756
rect 4970 1656 4972 1664
rect 4980 1656 4982 1664
rect 4970 1654 4982 1656
rect 5002 1324 5014 1996
rect 5034 1904 5046 3036
rect 5034 1896 5036 1904
rect 5044 1896 5046 1904
rect 5034 1504 5046 1896
rect 5034 1496 5036 1504
rect 5044 1496 5046 1504
rect 5034 1494 5046 1496
rect 5098 2524 5110 2526
rect 5098 2516 5100 2524
rect 5108 2516 5110 2524
rect 5002 1316 5004 1324
rect 5012 1316 5014 1324
rect 5002 1314 5014 1316
rect 5066 1264 5078 1266
rect 5066 1256 5068 1264
rect 5076 1256 5078 1264
rect 5034 1124 5046 1126
rect 5034 1116 5036 1124
rect 5044 1116 5046 1124
rect 4970 1004 4982 1006
rect 4970 996 4972 1004
rect 4980 996 4982 1004
rect 4970 764 4982 996
rect 4970 756 4972 764
rect 4980 756 4982 764
rect 4970 754 4982 756
rect 5034 724 5046 1116
rect 5034 716 5036 724
rect 5044 716 5046 724
rect 5034 714 5046 716
rect 5002 704 5014 706
rect 5002 696 5004 704
rect 5012 696 5014 704
rect 4874 316 4876 324
rect 4884 316 4886 324
rect 4874 314 4886 316
rect 4970 444 4982 446
rect 4970 436 4972 444
rect 4980 436 4982 444
rect 4714 236 4716 244
rect 4724 236 4726 244
rect 4714 234 4726 236
rect 4970 244 4982 436
rect 4970 236 4972 244
rect 4980 236 4982 244
rect 4970 234 4982 236
rect 5002 244 5014 696
rect 5002 236 5004 244
rect 5012 236 5014 244
rect 5002 234 5014 236
rect 5034 464 5046 466
rect 5034 456 5036 464
rect 5044 456 5046 464
rect 5034 224 5046 456
rect 5066 464 5078 1256
rect 5098 704 5110 2516
rect 5226 2224 5238 3436
rect 5258 2804 5270 3676
rect 5386 3444 5398 3446
rect 5386 3436 5388 3444
rect 5396 3436 5398 3444
rect 5258 2796 5260 2804
rect 5268 2796 5270 2804
rect 5258 2794 5270 2796
rect 5322 3004 5334 3006
rect 5322 2996 5324 3004
rect 5332 2996 5334 3004
rect 5226 2216 5228 2224
rect 5236 2216 5238 2224
rect 5226 2214 5238 2216
rect 5258 2264 5270 2266
rect 5258 2256 5260 2264
rect 5268 2256 5270 2264
rect 5226 2044 5238 2046
rect 5226 2036 5228 2044
rect 5236 2036 5238 2044
rect 5098 696 5100 704
rect 5108 696 5110 704
rect 5098 694 5110 696
rect 5194 1544 5206 1546
rect 5194 1536 5196 1544
rect 5204 1536 5206 1544
rect 5066 456 5068 464
rect 5076 456 5078 464
rect 5066 454 5078 456
rect 5194 384 5206 1536
rect 5194 376 5196 384
rect 5204 376 5206 384
rect 5194 374 5206 376
rect 5226 324 5238 2036
rect 5258 1724 5270 2256
rect 5322 1924 5334 2996
rect 5354 2964 5366 2966
rect 5354 2956 5356 2964
rect 5364 2956 5366 2964
rect 5354 2124 5366 2956
rect 5354 2116 5356 2124
rect 5364 2116 5366 2124
rect 5354 2114 5366 2116
rect 5322 1916 5324 1924
rect 5332 1916 5334 1924
rect 5322 1914 5334 1916
rect 5386 1884 5398 3436
rect 5386 1876 5388 1884
rect 5396 1876 5398 1884
rect 5386 1874 5398 1876
rect 5418 2584 5430 2586
rect 5418 2576 5420 2584
rect 5428 2576 5430 2584
rect 5258 1716 5260 1724
rect 5268 1716 5270 1724
rect 5258 1714 5270 1716
rect 5322 1764 5334 1766
rect 5322 1756 5324 1764
rect 5332 1756 5334 1764
rect 5322 1704 5334 1756
rect 5322 1696 5324 1704
rect 5332 1696 5334 1704
rect 5322 1694 5334 1696
rect 5322 1404 5334 1406
rect 5322 1396 5324 1404
rect 5332 1396 5334 1404
rect 5322 384 5334 1396
rect 5322 376 5324 384
rect 5332 376 5334 384
rect 5322 374 5334 376
rect 5418 344 5430 2576
rect 5514 2364 5526 2366
rect 5514 2356 5516 2364
rect 5524 2356 5526 2364
rect 5514 2284 5526 2356
rect 5514 2276 5516 2284
rect 5524 2276 5526 2284
rect 5514 2274 5526 2276
rect 5418 336 5420 344
rect 5428 336 5430 344
rect 5418 334 5430 336
rect 5450 1804 5462 1806
rect 5450 1796 5452 1804
rect 5460 1796 5462 1804
rect 5226 316 5228 324
rect 5236 316 5238 324
rect 5226 314 5238 316
rect 5034 216 5036 224
rect 5044 216 5046 224
rect 5034 214 5046 216
rect 5450 124 5462 1796
rect 5450 116 5452 124
rect 5460 116 5462 124
rect 5450 114 5462 116
rect 4522 16 4524 24
rect 4532 16 4534 24
rect 4522 14 4534 16
rect 4224 6 4228 14
rect 4236 6 4240 14
rect 4248 6 4252 14
rect 4260 6 4264 14
rect 4272 6 4276 14
rect 4284 6 4288 14
rect 4224 -10 4288 6
use DFFSR  _1723_
timestamp 1618002947
transform -1 0 360 0 -1 210
box -4 -6 356 206
use DFFSR  _1704_
timestamp 1618002947
transform 1 0 360 0 -1 210
box -4 -6 356 206
use DFFSR  _1722_
timestamp 1618002947
transform -1 0 360 0 1 210
box -4 -6 356 206
use DFFSR  _1721_
timestamp 1618002947
transform -1 0 712 0 1 210
box -4 -6 356 206
use AND2X2  _1408_
timestamp 1618002947
transform -1 0 776 0 -1 210
box -4 -6 68 206
use BUFX2  _1754_
timestamp 1618002947
transform -1 0 760 0 1 210
box -4 -6 52 206
use AND2X2  _1409_
timestamp 1618002947
transform 1 0 776 0 -1 210
box -4 -6 68 206
use DFFSR  _1705_
timestamp 1618002947
transform 1 0 840 0 -1 210
box -4 -6 356 206
use CLKBUF1  CLKBUF1_insert14
timestamp 1618002947
transform 1 0 760 0 1 210
box -4 -6 148 206
use DFFSR  _1681_
timestamp 1618002947
transform 1 0 904 0 1 210
box -4 -6 356 206
use FILL  SFILL12560x2100
timestamp 1618002947
transform 1 0 1256 0 1 210
box -4 -6 20 206
use FILL  SFILL12560x100
timestamp 1618002947
transform -1 0 1272 0 -1 210
box -4 -6 20 206
use FILL  SFILL12400x100
timestamp 1618002947
transform -1 0 1256 0 -1 210
box -4 -6 20 206
use NOR2X1  _1319_
timestamp 1618002947
transform 1 0 1192 0 -1 210
box -4 -6 52 206
use FILL  SFILL13040x2100
timestamp 1618002947
transform 1 0 1304 0 1 210
box -4 -6 20 206
use FILL  SFILL12880x2100
timestamp 1618002947
transform 1 0 1288 0 1 210
box -4 -6 20 206
use FILL  SFILL12720x2100
timestamp 1618002947
transform 1 0 1272 0 1 210
box -4 -6 20 206
use FILL  SFILL12880x100
timestamp 1618002947
transform -1 0 1304 0 -1 210
box -4 -6 20 206
use FILL  SFILL12720x100
timestamp 1618002947
transform -1 0 1288 0 -1 210
box -4 -6 20 206
use OAI21X1  _1318_
timestamp 1618002947
transform -1 0 1368 0 -1 210
box -4 -6 68 206
use DFFSR  _1684_
timestamp 1618002947
transform -1 0 1672 0 1 210
box -4 -6 356 206
use DFFSR  _1682_
timestamp 1618002947
transform -1 0 1720 0 -1 210
box -4 -6 356 206
use BUFX2  _1751_
timestamp 1618002947
transform -1 0 1768 0 -1 210
box -4 -6 52 206
use BUFX2  _1753_
timestamp 1618002947
transform 1 0 1768 0 -1 210
box -4 -6 52 206
use DFFSR  _1685_
timestamp 1618002947
transform -1 0 2024 0 1 210
box -4 -6 356 206
use DFFSR  _1711_
timestamp 1618002947
transform 1 0 1816 0 -1 210
box -4 -6 356 206
use INVX1  _1417_
timestamp 1618002947
transform 1 0 2168 0 -1 210
box -4 -6 36 206
use NAND2X1  _1422_
timestamp 1618002947
transform 1 0 2024 0 1 210
box -4 -6 52 206
use OAI21X1  _1421_
timestamp 1618002947
transform -1 0 2136 0 1 210
box -4 -6 68 206
use INVX1  _1419_
timestamp 1618002947
transform 1 0 2136 0 1 210
box -4 -6 36 206
use OAI21X1  _1420_
timestamp 1618002947
transform 1 0 2168 0 1 210
box -4 -6 68 206
use OAI21X1  _1440_
timestamp 1618002947
transform 1 0 2200 0 -1 210
box -4 -6 68 206
use OAI21X1  _1439_
timestamp 1618002947
transform 1 0 2264 0 -1 210
box -4 -6 68 206
use NAND2X1  _1428_
timestamp 1618002947
transform 1 0 2328 0 -1 210
box -4 -6 52 206
use OAI21X1  _1427_
timestamp 1618002947
transform 1 0 2376 0 -1 210
box -4 -6 68 206
use OAI21X1  _1435_
timestamp 1618002947
transform 1 0 2440 0 -1 210
box -4 -6 68 206
use OAI21X1  _1436_
timestamp 1618002947
transform -1 0 2568 0 -1 210
box -4 -6 68 206
use OAI21X1  _1441_
timestamp 1618002947
transform 1 0 2232 0 1 210
box -4 -6 68 206
use DFFSR  _1708_
timestamp 1618002947
transform -1 0 2648 0 1 210
box -4 -6 356 206
use OAI21X1  _1434_
timestamp 1618002947
transform 1 0 2680 0 1 210
box -4 -6 68 206
use INVX1  _1423_
timestamp 1618002947
transform 1 0 2648 0 1 210
box -4 -6 36 206
use OAI21X1  _1437_
timestamp 1618002947
transform 1 0 2696 0 -1 210
box -4 -6 68 206
use INVX1  _1425_
timestamp 1618002947
transform 1 0 2664 0 -1 210
box -4 -6 36 206
use INVX1  _1424_
timestamp 1618002947
transform -1 0 2664 0 -1 210
box -4 -6 36 206
use OAI21X1  _1426_
timestamp 1618002947
transform -1 0 2632 0 -1 210
box -4 -6 68 206
use FILL  SFILL27600x100
timestamp 1618002947
transform -1 0 2776 0 -1 210
box -4 -6 20 206
use FILL  SFILL27760x100
timestamp 1618002947
transform -1 0 2792 0 -1 210
box -4 -6 20 206
use FILL  SFILL27440x2100
timestamp 1618002947
transform 1 0 2744 0 1 210
box -4 -6 20 206
use FILL  SFILL27600x2100
timestamp 1618002947
transform 1 0 2760 0 1 210
box -4 -6 20 206
use FILL  SFILL27760x2100
timestamp 1618002947
transform 1 0 2776 0 1 210
box -4 -6 20 206
use OAI21X1  _1438_
timestamp 1618002947
transform 1 0 2824 0 -1 210
box -4 -6 68 206
use OAI21X1  _1433_
timestamp 1618002947
transform -1 0 2872 0 1 210
box -4 -6 68 206
use FILL  SFILL27920x100
timestamp 1618002947
transform -1 0 2808 0 -1 210
box -4 -6 20 206
use FILL  SFILL28080x100
timestamp 1618002947
transform -1 0 2824 0 -1 210
box -4 -6 20 206
use FILL  SFILL27920x2100
timestamp 1618002947
transform 1 0 2792 0 1 210
box -4 -6 20 206
use DFFSR  _1710_
timestamp 1618002947
transform -1 0 3224 0 1 210
box -4 -6 356 206
use DFFSR  _1709_
timestamp 1618002947
transform -1 0 3240 0 -1 210
box -4 -6 356 206
use AND2X2  _1410_
timestamp 1618002947
transform 1 0 3240 0 -1 210
box -4 -6 68 206
use DFFSR  _1703_
timestamp 1618002947
transform -1 0 3576 0 1 210
box -4 -6 356 206
use AND2X2  _1411_
timestamp 1618002947
transform 1 0 3304 0 -1 210
box -4 -6 68 206
use DFFSR  _1702_
timestamp 1618002947
transform -1 0 3720 0 -1 210
box -4 -6 356 206
use CLKBUF1  CLKBUF1_insert16
timestamp 1618002947
transform -1 0 3720 0 1 210
box -4 -6 148 206
use BUFX2  _1756_
timestamp 1618002947
transform -1 0 3768 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _1010_
timestamp 1618002947
transform -1 0 3960 0 -1 210
box -4 -6 196 206
use DFFSR  _1034_
timestamp 1618002947
transform 1 0 3960 0 -1 210
box -4 -6 356 206
use DFFSR  _1063_
timestamp 1618002947
transform 1 0 3720 0 1 210
box -4 -6 356 206
use INVX1  _871_
timestamp 1618002947
transform 1 0 4072 0 1 210
box -4 -6 36 206
use DFFSR  _1032_
timestamp 1618002947
transform 1 0 4168 0 1 210
box -4 -6 356 206
use FILL  SFILL43120x100
timestamp 1618002947
transform -1 0 4328 0 -1 210
box -4 -6 20 206
use FILL  SFILL43280x100
timestamp 1618002947
transform -1 0 4344 0 -1 210
box -4 -6 20 206
use FILL  SFILL41040x2100
timestamp 1618002947
transform 1 0 4104 0 1 210
box -4 -6 20 206
use FILL  SFILL41200x2100
timestamp 1618002947
transform 1 0 4120 0 1 210
box -4 -6 20 206
use FILL  SFILL41360x2100
timestamp 1618002947
transform 1 0 4136 0 1 210
box -4 -6 20 206
use FILL  SFILL41520x2100
timestamp 1618002947
transform 1 0 4152 0 1 210
box -4 -6 20 206
use DFFPOSX1  _1013_
timestamp 1618002947
transform 1 0 4376 0 -1 210
box -4 -6 196 206
use BUFX2  _1759_
timestamp 1618002947
transform 1 0 4568 0 -1 210
box -4 -6 52 206
use BUFX2  _1757_
timestamp 1618002947
transform 1 0 4616 0 -1 210
box -4 -6 52 206
use DFFSR  _1033_
timestamp 1618002947
transform 1 0 4664 0 -1 210
box -4 -6 356 206
use DFFPOSX1  _1011_
timestamp 1618002947
transform -1 0 4712 0 1 210
box -4 -6 196 206
use FILL  SFILL43440x100
timestamp 1618002947
transform -1 0 4360 0 -1 210
box -4 -6 20 206
use FILL  SFILL43600x100
timestamp 1618002947
transform -1 0 4376 0 -1 210
box -4 -6 20 206
use INVX1  _863_
timestamp 1618002947
transform 1 0 5016 0 -1 210
box -4 -6 36 206
use DFFSR  _1019_
timestamp 1618002947
transform 1 0 5048 0 -1 210
box -4 -6 356 206
use INVX1  _926_
timestamp 1618002947
transform 1 0 4712 0 1 210
box -4 -6 36 206
use OAI21X1  _928_
timestamp 1618002947
transform 1 0 4744 0 1 210
box -4 -6 68 206
use DFFSR  _1229_
timestamp 1618002947
transform -1 0 5160 0 1 210
box -4 -6 356 206
use BUFX2  _1764_
timestamp 1618002947
transform 1 0 5400 0 -1 210
box -4 -6 52 206
use MUX2X1  _934_
timestamp 1618002947
transform -1 0 5256 0 1 210
box -4 -6 100 206
use MUX2X1  _936_
timestamp 1618002947
transform 1 0 5256 0 1 210
box -4 -6 100 206
use CLKBUF1  CLKBUF1_insert9
timestamp 1618002947
transform 1 0 5352 0 1 210
box -4 -6 148 206
use BUFX2  _1762_
timestamp 1618002947
transform 1 0 5448 0 -1 210
box -4 -6 52 206
use FILL  FILL53040x100
timestamp 1618002947
transform -1 0 5512 0 -1 210
box -4 -6 20 206
use FILL  FILL53040x2100
timestamp 1618002947
transform 1 0 5496 0 1 210
box -4 -6 20 206
use INVX1  _1490_
timestamp 1618002947
transform 1 0 8 0 -1 610
box -4 -6 36 206
use NAND2X1  _1495_
timestamp 1618002947
transform 1 0 40 0 -1 610
box -4 -6 52 206
use INVX1  _1494_
timestamp 1618002947
transform 1 0 88 0 -1 610
box -4 -6 36 206
use NAND2X1  _1491_
timestamp 1618002947
transform 1 0 120 0 -1 610
box -4 -6 52 206
use OAI22X1  _1545_
timestamp 1618002947
transform 1 0 168 0 -1 610
box -4 -6 84 206
use OAI22X1  _1544_
timestamp 1618002947
transform 1 0 248 0 -1 610
box -4 -6 84 206
use NAND2X1  _1292_
timestamp 1618002947
transform 1 0 328 0 -1 610
box -4 -6 52 206
use INVX1  _1291_
timestamp 1618002947
transform -1 0 408 0 -1 610
box -4 -6 36 206
use DFFSR  _1715_
timestamp 1618002947
transform 1 0 408 0 -1 610
box -4 -6 356 206
use CLKBUF1  CLKBUF1_insert15
timestamp 1618002947
transform 1 0 760 0 -1 610
box -4 -6 148 206
use DFFSR  _1687_
timestamp 1618002947
transform 1 0 904 0 -1 610
box -4 -6 356 206
use NOR2X1  _1323_
timestamp 1618002947
transform 1 0 1320 0 -1 610
box -4 -6 52 206
use INVX1  _1324_
timestamp 1618002947
transform -1 0 1400 0 -1 610
box -4 -6 36 206
use NOR2X1  _1326_
timestamp 1618002947
transform -1 0 1448 0 -1 610
box -4 -6 52 206
use NAND2X1  _1325_
timestamp 1618002947
transform -1 0 1496 0 -1 610
box -4 -6 52 206
use FILL  SFILL12560x4100
timestamp 1618002947
transform -1 0 1272 0 -1 610
box -4 -6 20 206
use FILL  SFILL12720x4100
timestamp 1618002947
transform -1 0 1288 0 -1 610
box -4 -6 20 206
use FILL  SFILL12880x4100
timestamp 1618002947
transform -1 0 1304 0 -1 610
box -4 -6 20 206
use FILL  SFILL13040x4100
timestamp 1618002947
transform -1 0 1320 0 -1 610
box -4 -6 20 206
use NAND2X1  _1322_
timestamp 1618002947
transform 1 0 1496 0 -1 610
box -4 -6 52 206
use NOR2X1  _1321_
timestamp 1618002947
transform 1 0 1544 0 -1 610
box -4 -6 52 206
use NAND2X1  _1416_
timestamp 1618002947
transform -1 0 1640 0 -1 610
box -4 -6 52 206
use INVX1  _1320_
timestamp 1618002947
transform -1 0 1672 0 -1 610
box -4 -6 36 206
use NOR2X1  _1315_
timestamp 1618002947
transform -1 0 1720 0 -1 610
box -4 -6 52 206
use INVX4  _1262_
timestamp 1618002947
transform 1 0 1720 0 -1 610
box -4 -6 52 206
use DFFSR  _1713_
timestamp 1618002947
transform 1 0 1768 0 -1 610
box -4 -6 356 206
use OAI21X1  _1444_
timestamp 1618002947
transform 1 0 2120 0 -1 610
box -4 -6 68 206
use OAI21X1  _1443_
timestamp 1618002947
transform -1 0 2248 0 -1 610
box -4 -6 68 206
use INVX1  _1418_
timestamp 1618002947
transform -1 0 2280 0 -1 610
box -4 -6 36 206
use OAI21X1  _1442_
timestamp 1618002947
transform 1 0 2280 0 -1 610
box -4 -6 68 206
use DFFSR  _1712_
timestamp 1618002947
transform -1 0 2696 0 -1 610
box -4 -6 356 206
use BUFX2  BUFX2_insert4
timestamp 1618002947
transform 1 0 2696 0 -1 610
box -4 -6 52 206
use DFFSR  _1057_
timestamp 1618002947
transform 1 0 2808 0 -1 610
box -4 -6 356 206
use FILL  SFILL27440x4100
timestamp 1618002947
transform -1 0 2760 0 -1 610
box -4 -6 20 206
use FILL  SFILL27600x4100
timestamp 1618002947
transform -1 0 2776 0 -1 610
box -4 -6 20 206
use FILL  SFILL27760x4100
timestamp 1618002947
transform -1 0 2792 0 -1 610
box -4 -6 20 206
use FILL  SFILL27920x4100
timestamp 1618002947
transform -1 0 2808 0 -1 610
box -4 -6 20 206
use INVX1  _903_
timestamp 1618002947
transform 1 0 3160 0 -1 610
box -4 -6 36 206
use DFFSR  _1025_
timestamp 1618002947
transform 1 0 3192 0 -1 610
box -4 -6 356 206
use NOR2X1  _904_
timestamp 1618002947
transform 1 0 3544 0 -1 610
box -4 -6 52 206
use INVX1  _902_
timestamp 1618002947
transform 1 0 3592 0 -1 610
box -4 -6 36 206
use OAI21X1  _906_
timestamp 1618002947
transform 1 0 3624 0 -1 610
box -4 -6 68 206
use NAND2X1  _905_
timestamp 1618002947
transform -1 0 3736 0 -1 610
box -4 -6 52 206
use DFFSR  _1039_
timestamp 1618002947
transform 1 0 3736 0 -1 610
box -4 -6 356 206
use MUX2X1  _930_
timestamp 1618002947
transform -1 0 4184 0 -1 610
box -4 -6 100 206
use INVX1  _929_
timestamp 1618002947
transform -1 0 4216 0 -1 610
box -4 -6 36 206
use MUX2X1  _909_
timestamp 1618002947
transform -1 0 4376 0 -1 610
box -4 -6 100 206
use FILL  SFILL42160x4100
timestamp 1618002947
transform -1 0 4232 0 -1 610
box -4 -6 20 206
use FILL  SFILL42320x4100
timestamp 1618002947
transform -1 0 4248 0 -1 610
box -4 -6 20 206
use FILL  SFILL42480x4100
timestamp 1618002947
transform -1 0 4264 0 -1 610
box -4 -6 20 206
use FILL  SFILL42640x4100
timestamp 1618002947
transform -1 0 4280 0 -1 610
box -4 -6 20 206
use INVX1  _907_
timestamp 1618002947
transform -1 0 4408 0 -1 610
box -4 -6 36 206
use DFFSR  _1026_
timestamp 1618002947
transform -1 0 4760 0 -1 610
box -4 -6 356 206
use NAND2X1  _927_
timestamp 1618002947
transform 1 0 4760 0 -1 610
box -4 -6 52 206
use MUX2X1  _1140_
timestamp 1618002947
transform -1 0 4904 0 -1 610
box -4 -6 100 206
use MUX2X1  _1143_
timestamp 1618002947
transform 1 0 4904 0 -1 610
box -4 -6 100 206
use OAI21X1  _1144_
timestamp 1618002947
transform 1 0 5000 0 -1 610
box -4 -6 68 206
use OAI21X1  _1141_
timestamp 1618002947
transform 1 0 5064 0 -1 610
box -4 -6 68 206
use DFFSR  _1230_
timestamp 1618002947
transform -1 0 5480 0 -1 610
box -4 -6 356 206
use FILL  FILL52880x4100
timestamp 1618002947
transform -1 0 5496 0 -1 610
box -4 -6 20 206
use FILL  FILL53040x4100
timestamp 1618002947
transform -1 0 5512 0 -1 610
box -4 -6 20 206
use NOR2X1  _1269_
timestamp 1618002947
transform 1 0 8 0 1 610
box -4 -6 52 206
use INVX1  _1489_
timestamp 1618002947
transform 1 0 56 0 1 610
box -4 -6 36 206
use NOR2X1  _1496_
timestamp 1618002947
transform 1 0 88 0 1 610
box -4 -6 52 206
use NOR2X1  _1492_
timestamp 1618002947
transform -1 0 184 0 1 610
box -4 -6 52 206
use INVX1  _1290_
timestamp 1618002947
transform 1 0 184 0 1 610
box -4 -6 36 206
use NOR2X1  _1499_
timestamp 1618002947
transform -1 0 264 0 1 610
box -4 -6 52 206
use NOR2X1  _1293_
timestamp 1618002947
transform -1 0 312 0 1 610
box -4 -6 52 206
use NOR2X1  _1270_
timestamp 1618002947
transform -1 0 360 0 1 610
box -4 -6 52 206
use NAND2X1  _1498_
timestamp 1618002947
transform -1 0 408 0 1 610
box -4 -6 52 206
use INVX1  _1497_
timestamp 1618002947
transform -1 0 440 0 1 610
box -4 -6 36 206
use OAI22X1  _1543_
timestamp 1618002947
transform 1 0 440 0 1 610
box -4 -6 84 206
use OAI21X1  _1504_
timestamp 1618002947
transform 1 0 520 0 1 610
box -4 -6 68 206
use NAND2X1  _1451_
timestamp 1618002947
transform -1 0 632 0 1 610
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert6
timestamp 1618002947
transform -1 0 776 0 1 610
box -4 -6 148 206
use NAND3X1  _1316_
timestamp 1618002947
transform 1 0 776 0 1 610
box -4 -6 68 206
use NAND3X1  _1314_
timestamp 1618002947
transform -1 0 904 0 1 610
box -4 -6 68 206
use DFFSR  _1683_
timestamp 1618002947
transform -1 0 1256 0 1 610
box -4 -6 356 206
use DFFSR  _1686_
timestamp 1618002947
transform -1 0 1672 0 1 610
box -4 -6 356 206
use FILL  SFILL12560x6100
timestamp 1618002947
transform 1 0 1256 0 1 610
box -4 -6 20 206
use FILL  SFILL12720x6100
timestamp 1618002947
transform 1 0 1272 0 1 610
box -4 -6 20 206
use FILL  SFILL12880x6100
timestamp 1618002947
transform 1 0 1288 0 1 610
box -4 -6 20 206
use FILL  SFILL13040x6100
timestamp 1618002947
transform 1 0 1304 0 1 610
box -4 -6 20 206
use BUFX2  BUFX2_insert19
timestamp 1618002947
transform -1 0 1720 0 1 610
box -4 -6 52 206
use DFFSR  _1694_
timestamp 1618002947
transform 1 0 1720 0 1 610
box -4 -6 356 206
use DFFSR  _1693_
timestamp 1618002947
transform -1 0 2424 0 1 610
box -4 -6 356 206
use BUFX2  BUFX2_insert3
timestamp 1618002947
transform -1 0 2472 0 1 610
box -4 -6 52 206
use INVX1  _993_
timestamp 1618002947
transform 1 0 2472 0 1 610
box -4 -6 36 206
use OAI21X1  _995_
timestamp 1618002947
transform 1 0 2504 0 1 610
box -4 -6 68 206
use OAI21X1  _994_
timestamp 1618002947
transform -1 0 2632 0 1 610
box -4 -6 68 206
use INVX1  _809_
timestamp 1618002947
transform 1 0 2632 0 1 610
box -4 -6 36 206
use DFFSR  _1055_
timestamp 1618002947
transform -1 0 3080 0 1 610
box -4 -6 356 206
use FILL  SFILL26640x6100
timestamp 1618002947
transform 1 0 2664 0 1 610
box -4 -6 20 206
use FILL  SFILL26800x6100
timestamp 1618002947
transform 1 0 2680 0 1 610
box -4 -6 20 206
use FILL  SFILL26960x6100
timestamp 1618002947
transform 1 0 2696 0 1 610
box -4 -6 20 206
use FILL  SFILL27120x6100
timestamp 1618002947
transform 1 0 2712 0 1 610
box -4 -6 20 206
use OAI21X1  _990_
timestamp 1618002947
transform 1 0 3080 0 1 610
box -4 -6 68 206
use OAI21X1  _989_
timestamp 1618002947
transform -1 0 3208 0 1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert5
timestamp 1618002947
transform 1 0 3208 0 1 610
box -4 -6 52 206
use OAI22X1  _828_
timestamp 1618002947
transform -1 0 3336 0 1 610
box -4 -6 84 206
use INVX1  _826_
timestamp 1618002947
transform -1 0 3368 0 1 610
box -4 -6 36 206
use DFFSR  _1024_
timestamp 1618002947
transform -1 0 3720 0 1 610
box -4 -6 356 206
use OAI21X1  _901_
timestamp 1618002947
transform 1 0 3720 0 1 610
box -4 -6 68 206
use OAI22X1  _814_
timestamp 1618002947
transform -1 0 3864 0 1 610
box -4 -6 84 206
use OAI21X1  _1009_
timestamp 1618002947
transform 1 0 3864 0 1 610
box -4 -6 68 206
use INVX1  _808_
timestamp 1618002947
transform -1 0 3960 0 1 610
box -4 -6 36 206
use NAND2X1  _825_
timestamp 1618002947
transform -1 0 4008 0 1 610
box -4 -6 52 206
use NOR2X1  _791_
timestamp 1618002947
transform -1 0 4056 0 1 610
box -4 -6 52 206
use INVX1  _795_
timestamp 1618002947
transform 1 0 4056 0 1 610
box -4 -6 36 206
use DFFSR  _1022_
timestamp 1618002947
transform -1 0 4504 0 1 610
box -4 -6 356 206
use FILL  SFILL40880x6100
timestamp 1618002947
transform 1 0 4088 0 1 610
box -4 -6 20 206
use FILL  SFILL41040x6100
timestamp 1618002947
transform 1 0 4104 0 1 610
box -4 -6 20 206
use FILL  SFILL41200x6100
timestamp 1618002947
transform 1 0 4120 0 1 610
box -4 -6 20 206
use FILL  SFILL41360x6100
timestamp 1618002947
transform 1 0 4136 0 1 610
box -4 -6 20 206
use OAI21X1  _925_
timestamp 1618002947
transform -1 0 4568 0 1 610
box -4 -6 68 206
use INVX1  _830_
timestamp 1618002947
transform -1 0 4600 0 1 610
box -4 -6 36 206
use AOI21X1  _815_
timestamp 1618002947
transform -1 0 4664 0 1 610
box -4 -6 68 206
use NAND2X1  _837_
timestamp 1618002947
transform -1 0 4712 0 1 610
box -4 -6 52 206
use AOI21X1  _829_
timestamp 1618002947
transform -1 0 4776 0 1 610
box -4 -6 68 206
use MUX2X1  _1146_
timestamp 1618002947
transform -1 0 4872 0 1 610
box -4 -6 100 206
use NAND2X1  _1134_
timestamp 1618002947
transform 1 0 4872 0 1 610
box -4 -6 52 206
use OAI21X1  _1138_
timestamp 1618002947
transform 1 0 4920 0 1 610
box -4 -6 68 206
use OAI21X1  _1147_
timestamp 1618002947
transform -1 0 5048 0 1 610
box -4 -6 68 206
use NAND2X1  _1142_
timestamp 1618002947
transform -1 0 5096 0 1 610
box -4 -6 52 206
use NAND2X1  _1139_
timestamp 1618002947
transform -1 0 5144 0 1 610
box -4 -6 52 206
use DFFSR  _1231_
timestamp 1618002947
transform -1 0 5496 0 1 610
box -4 -6 356 206
use FILL  FILL53040x6100
timestamp 1618002947
transform 1 0 5496 0 1 610
box -4 -6 20 206
use NAND2X1  _1311_
timestamp 1618002947
transform 1 0 8 0 -1 1010
box -4 -6 52 206
use NOR2X1  _1312_
timestamp 1618002947
transform -1 0 104 0 -1 1010
box -4 -6 52 206
use NAND3X1  _1517_
timestamp 1618002947
transform -1 0 168 0 -1 1010
box -4 -6 68 206
use NAND3X1  _1516_
timestamp 1618002947
transform -1 0 232 0 -1 1010
box -4 -6 68 206
use OAI21X1  _1500_
timestamp 1618002947
transform 1 0 232 0 -1 1010
box -4 -6 68 206
use NAND2X1  _1493_
timestamp 1618002947
transform 1 0 296 0 -1 1010
box -4 -6 52 206
use NAND2X1  _1501_
timestamp 1618002947
transform 1 0 344 0 -1 1010
box -4 -6 52 206
use OAI21X1  _1580_
timestamp 1618002947
transform 1 0 392 0 -1 1010
box -4 -6 68 206
use DFFSR  _1733_
timestamp 1618002947
transform 1 0 456 0 -1 1010
box -4 -6 356 206
use OAI21X1  _1317_
timestamp 1618002947
transform -1 0 872 0 -1 1010
box -4 -6 68 206
use NOR2X1  _1576_
timestamp 1618002947
transform 1 0 872 0 -1 1010
box -4 -6 52 206
use AOI21X1  _1577_
timestamp 1618002947
transform -1 0 984 0 -1 1010
box -4 -6 68 206
use DFFSR  _1692_
timestamp 1618002947
transform 1 0 984 0 -1 1010
box -4 -6 356 206
use INVX1  _1333_
timestamp 1618002947
transform -1 0 1432 0 -1 1010
box -4 -6 36 206
use OR2X2  _1429_
timestamp 1618002947
transform 1 0 1432 0 -1 1010
box -4 -6 68 206
use FILL  SFILL13360x8100
timestamp 1618002947
transform -1 0 1352 0 -1 1010
box -4 -6 20 206
use FILL  SFILL13520x8100
timestamp 1618002947
transform -1 0 1368 0 -1 1010
box -4 -6 20 206
use FILL  SFILL13680x8100
timestamp 1618002947
transform -1 0 1384 0 -1 1010
box -4 -6 20 206
use FILL  SFILL13840x8100
timestamp 1618002947
transform -1 0 1400 0 -1 1010
box -4 -6 20 206
use OAI21X1  _1431_
timestamp 1618002947
transform -1 0 1560 0 -1 1010
box -4 -6 68 206
use DFFPOSX1  _1678_
timestamp 1618002947
transform 1 0 1560 0 -1 1010
box -4 -6 196 206
use BUFX2  BUFX2_insert27
timestamp 1618002947
transform 1 0 1752 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert25
timestamp 1618002947
transform 1 0 1800 0 -1 1010
box -4 -6 52 206
use INVX1  _1371_
timestamp 1618002947
transform 1 0 1848 0 -1 1010
box -4 -6 36 206
use AOI21X1  _1375_
timestamp 1618002947
transform 1 0 1880 0 -1 1010
box -4 -6 68 206
use NAND2X1  _1374_
timestamp 1618002947
transform 1 0 1944 0 -1 1010
box -4 -6 52 206
use NAND2X1  _1373_
timestamp 1618002947
transform -1 0 2040 0 -1 1010
box -4 -6 52 206
use OAI21X1  _1372_
timestamp 1618002947
transform -1 0 2104 0 -1 1010
box -4 -6 68 206
use INVX1  _1332_
timestamp 1618002947
transform -1 0 2136 0 -1 1010
box -4 -6 36 206
use NAND2X1  _1340_
timestamp 1618002947
transform 1 0 2136 0 -1 1010
box -4 -6 52 206
use NOR2X1  _1339_
timestamp 1618002947
transform 1 0 2184 0 -1 1010
box -4 -6 52 206
use NAND2X1  _1368_
timestamp 1618002947
transform 1 0 2232 0 -1 1010
box -4 -6 52 206
use INVX1  _1367_
timestamp 1618002947
transform 1 0 2280 0 -1 1010
box -4 -6 36 206
use AOI21X1  _1370_
timestamp 1618002947
transform -1 0 2376 0 -1 1010
box -4 -6 68 206
use OAI21X1  _1376_
timestamp 1618002947
transform 1 0 2376 0 -1 1010
box -4 -6 68 206
use NOR3X1  _1379_
timestamp 1618002947
transform 1 0 2440 0 -1 1010
box -4 -6 132 206
use NOR2X1  _1341_
timestamp 1618002947
transform -1 0 2616 0 -1 1010
box -4 -6 52 206
use DFFSR  _1695_
timestamp 1618002947
transform -1 0 3032 0 -1 1010
box -4 -6 356 206
use FILL  SFILL26160x8100
timestamp 1618002947
transform -1 0 2632 0 -1 1010
box -4 -6 20 206
use FILL  SFILL26320x8100
timestamp 1618002947
transform -1 0 2648 0 -1 1010
box -4 -6 20 206
use FILL  SFILL26480x8100
timestamp 1618002947
transform -1 0 2664 0 -1 1010
box -4 -6 20 206
use FILL  SFILL26640x8100
timestamp 1618002947
transform -1 0 2680 0 -1 1010
box -4 -6 20 206
use INVX1  _827_
timestamp 1618002947
transform 1 0 3032 0 -1 1010
box -4 -6 36 206
use DFFSR  _1056_
timestamp 1618002947
transform -1 0 3416 0 -1 1010
box -4 -6 356 206
use OAI21X1  _992_
timestamp 1618002947
transform 1 0 3416 0 -1 1010
box -4 -6 68 206
use OAI21X1  _991_
timestamp 1618002947
transform -1 0 3544 0 -1 1010
box -4 -6 68 206
use DFFSR  _1031_
timestamp 1618002947
transform 1 0 3544 0 -1 1010
box -4 -6 356 206
use NAND2X1  _900_
timestamp 1618002947
transform -1 0 3944 0 -1 1010
box -4 -6 52 206
use NAND2X1  _1008_
timestamp 1618002947
transform -1 0 3992 0 -1 1010
box -4 -6 52 206
use NAND2X1  _922_
timestamp 1618002947
transform 1 0 4040 0 -1 1010
box -4 -6 52 206
use NAND2X1  _790_
timestamp 1618002947
transform 1 0 3992 0 -1 1010
box -4 -6 52 206
use OAI21X1  _923_
timestamp 1618002947
transform -1 0 4152 0 -1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert18
timestamp 1618002947
transform -1 0 4232 0 -1 1010
box -4 -6 52 206
use INVX1  _816_
timestamp 1618002947
transform 1 0 4152 0 -1 1010
box -4 -6 36 206
use FILL  SFILL42480x8100
timestamp 1618002947
transform -1 0 4264 0 -1 1010
box -4 -6 20 206
use FILL  SFILL42320x8100
timestamp 1618002947
transform -1 0 4248 0 -1 1010
box -4 -6 20 206
use FILL  SFILL42800x8100
timestamp 1618002947
transform -1 0 4296 0 -1 1010
box -4 -6 20 206
use FILL  SFILL42640x8100
timestamp 1618002947
transform -1 0 4280 0 -1 1010
box -4 -6 20 206
use AOI21X1  _852_
timestamp 1618002947
transform -1 0 4392 0 -1 1010
box -4 -6 68 206
use INVX1  _792_
timestamp 1618002947
transform 1 0 4296 0 -1 1010
box -4 -6 36 206
use NAND3X1  _853_
timestamp 1618002947
transform 1 0 4392 0 -1 1010
box -4 -6 68 206
use NAND2X1  _924_
timestamp 1618002947
transform 1 0 4456 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert28
timestamp 1618002947
transform 1 0 4504 0 -1 1010
box -4 -6 52 206
use MUX2X1  _1135_
timestamp 1618002947
transform -1 0 4648 0 -1 1010
box -4 -6 100 206
use AOI22X1  _843_
timestamp 1618002947
transform 1 0 4648 0 -1 1010
box -4 -6 84 206
use AOI22X1  _849_
timestamp 1618002947
transform -1 0 4808 0 -1 1010
box -4 -6 84 206
use DFFSR  _1232_
timestamp 1618002947
transform -1 0 5160 0 -1 1010
box -4 -6 356 206
use DFFSR  _1233_
timestamp 1618002947
transform -1 0 5512 0 -1 1010
box -4 -6 356 206
use NAND3X1  _1470_
timestamp 1618002947
transform -1 0 72 0 1 1010
box -4 -6 68 206
use NAND2X1  _1271_
timestamp 1618002947
transform 1 0 72 0 1 1010
box -4 -6 52 206
use NAND3X1  _1518_
timestamp 1618002947
transform -1 0 184 0 1 1010
box -4 -6 68 206
use NAND3X1  _1519_
timestamp 1618002947
transform -1 0 248 0 1 1010
box -4 -6 68 206
use NAND3X1  _1507_
timestamp 1618002947
transform 1 0 248 0 1 1010
box -4 -6 68 206
use OAI21X1  _1538_
timestamp 1618002947
transform -1 0 376 0 1 1010
box -4 -6 68 206
use INVX4  _1531_
timestamp 1618002947
transform -1 0 424 0 1 1010
box -4 -6 52 206
use DFFSR  _1720_
timestamp 1618002947
transform -1 0 776 0 1 1010
box -4 -6 356 206
use OAI21X1  _1570_
timestamp 1618002947
transform 1 0 776 0 1 1010
box -4 -6 68 206
use DFFSR  _1680_
timestamp 1618002947
transform 1 0 840 0 1 1010
box -4 -6 356 206
use INVX1  _1313_
timestamp 1618002947
transform -1 0 1224 0 1 1010
box -4 -6 36 206
use NOR2X1  _1304_
timestamp 1618002947
transform -1 0 1336 0 1 1010
box -4 -6 52 206
use AOI21X1  _1366_
timestamp 1618002947
transform -1 0 1400 0 1 1010
box -4 -6 68 206
use INVX1  _1412_
timestamp 1618002947
transform 1 0 1400 0 1 1010
box -4 -6 36 206
use NOR2X1  _1261_
timestamp 1618002947
transform -1 0 1480 0 1 1010
box -4 -6 52 206
use FILL  SFILL12240x10100
timestamp 1618002947
transform 1 0 1224 0 1 1010
box -4 -6 20 206
use FILL  SFILL12400x10100
timestamp 1618002947
transform 1 0 1240 0 1 1010
box -4 -6 20 206
use FILL  SFILL12560x10100
timestamp 1618002947
transform 1 0 1256 0 1 1010
box -4 -6 20 206
use FILL  SFILL12720x10100
timestamp 1618002947
transform 1 0 1272 0 1 1010
box -4 -6 20 206
use OAI21X1  _1430_
timestamp 1618002947
transform 1 0 1480 0 1 1010
box -4 -6 68 206
use AOI21X1  _1264_
timestamp 1618002947
transform 1 0 1544 0 1 1010
box -4 -6 68 206
use NOR2X1  _1364_
timestamp 1618002947
transform 1 0 1608 0 1 1010
box -4 -6 52 206
use OAI21X1  _1365_
timestamp 1618002947
transform 1 0 1656 0 1 1010
box -4 -6 68 206
use INVX1  _1363_
timestamp 1618002947
transform -1 0 1752 0 1 1010
box -4 -6 36 206
use NAND2X1  _1338_
timestamp 1618002947
transform 1 0 1752 0 1 1010
box -4 -6 52 206
use DFFSR  _1696_
timestamp 1618002947
transform 1 0 1800 0 1 1010
box -4 -6 356 206
use AOI21X1  _1384_
timestamp 1618002947
transform -1 0 2216 0 1 1010
box -4 -6 68 206
use NAND2X1  _1383_
timestamp 1618002947
transform -1 0 2264 0 1 1010
box -4 -6 52 206
use OAI21X1  _1382_
timestamp 1618002947
transform -1 0 2328 0 1 1010
box -4 -6 68 206
use NOR2X1  _1381_
timestamp 1618002947
transform 1 0 2328 0 1 1010
box -4 -6 52 206
use INVX1  _1380_
timestamp 1618002947
transform -1 0 2408 0 1 1010
box -4 -6 36 206
use OR2X2  _1347_
timestamp 1618002947
transform 1 0 2408 0 1 1010
box -4 -6 68 206
use OAI21X1  _1432_
timestamp 1618002947
transform -1 0 2536 0 1 1010
box -4 -6 68 206
use OAI21X1  _1377_
timestamp 1618002947
transform 1 0 2536 0 1 1010
box -4 -6 68 206
use AOI21X1  _1378_
timestamp 1618002947
transform 1 0 2600 0 1 1010
box -4 -6 68 206
use DFFSR  _1049_
timestamp 1618002947
transform -1 0 3080 0 1 1010
box -4 -6 356 206
use FILL  SFILL26640x10100
timestamp 1618002947
transform 1 0 2664 0 1 1010
box -4 -6 20 206
use FILL  SFILL26800x10100
timestamp 1618002947
transform 1 0 2680 0 1 1010
box -4 -6 20 206
use FILL  SFILL26960x10100
timestamp 1618002947
transform 1 0 2696 0 1 1010
box -4 -6 20 206
use FILL  SFILL27120x10100
timestamp 1618002947
transform 1 0 2712 0 1 1010
box -4 -6 20 206
use OAI21X1  _971_
timestamp 1618002947
transform 1 0 3080 0 1 1010
box -4 -6 68 206
use OAI21X1  _972_
timestamp 1618002947
transform -1 0 3208 0 1 1010
box -4 -6 68 206
use INVX1  _970_
timestamp 1618002947
transform 1 0 3208 0 1 1010
box -4 -6 36 206
use CLKBUF1  CLKBUF1_insert17
timestamp 1618002947
transform -1 0 3384 0 1 1010
box -4 -6 148 206
use DFFSR  _1041_
timestamp 1618002947
transform 1 0 3384 0 1 1010
box -4 -6 356 206
use OAI22X1  _942_
timestamp 1618002947
transform -1 0 3816 0 1 1010
box -4 -6 84 206
use INVX1  _839_
timestamp 1618002947
transform -1 0 3848 0 1 1010
box -4 -6 36 206
use AOI22X1  _846_
timestamp 1618002947
transform 1 0 3848 0 1 1010
box -4 -6 84 206
use NOR2X1  _899_
timestamp 1618002947
transform -1 0 3976 0 1 1010
box -4 -6 52 206
use OAI22X1  _940_
timestamp 1618002947
transform -1 0 4136 0 1 1010
box -4 -6 84 206
use NOR2X1  _921_
timestamp 1618002947
transform -1 0 4056 0 1 1010
box -4 -6 52 206
use INVX1  _920_
timestamp 1618002947
transform 1 0 3976 0 1 1010
box -4 -6 36 206
use OAI21X1  _820_
timestamp 1618002947
transform -1 0 4200 0 1 1010
box -4 -6 68 206
use NOR2X1  _824_
timestamp 1618002947
transform -1 0 4248 0 1 1010
box -4 -6 52 206
use FILL  SFILL42960x10100
timestamp 1618002947
transform 1 0 4296 0 1 1010
box -4 -6 20 206
use FILL  SFILL42800x10100
timestamp 1618002947
transform 1 0 4280 0 1 1010
box -4 -6 20 206
use FILL  SFILL42640x10100
timestamp 1618002947
transform 1 0 4264 0 1 1010
box -4 -6 20 206
use FILL  SFILL42480x10100
timestamp 1618002947
transform 1 0 4248 0 1 1010
box -4 -6 20 206
use OAI22X1  _823_
timestamp 1618002947
transform -1 0 4392 0 1 1010
box -4 -6 84 206
use NAND3X1  _847_
timestamp 1618002947
transform 1 0 4392 0 1 1010
box -4 -6 68 206
use AOI21X1  _797_
timestamp 1618002947
transform 1 0 4456 0 1 1010
box -4 -6 68 206
use NAND2X1  _796_
timestamp 1618002947
transform -1 0 4568 0 1 1010
box -4 -6 52 206
use OAI21X1  _832_
timestamp 1618002947
transform 1 0 4568 0 1 1010
box -4 -6 68 206
use NOR2X1  _836_
timestamp 1618002947
transform 1 0 4632 0 1 1010
box -4 -6 52 206
use NAND2X1  _908_
timestamp 1618002947
transform 1 0 4680 0 1 1010
box -4 -6 52 206
use INVX2  _842_
timestamp 1618002947
transform 1 0 4728 0 1 1010
box -4 -6 36 206
use AOI22X1  _856_
timestamp 1618002947
transform 1 0 4760 0 1 1010
box -4 -6 84 206
use MUX2X1  _1149_
timestamp 1618002947
transform 1 0 4840 0 1 1010
box -4 -6 100 206
use NAND2X1  _1145_
timestamp 1618002947
transform 1 0 4936 0 1 1010
box -4 -6 52 206
use OAI21X1  _1150_
timestamp 1618002947
transform 1 0 4984 0 1 1010
box -4 -6 68 206
use NAND2X1  _1148_
timestamp 1618002947
transform -1 0 5096 0 1 1010
box -4 -6 52 206
use OAI21X1  _1153_
timestamp 1618002947
transform -1 0 5160 0 1 1010
box -4 -6 68 206
use DFFSR  _1234_
timestamp 1618002947
transform -1 0 5512 0 1 1010
box -4 -6 356 206
use INVX2  _1310_
timestamp 1618002947
transform -1 0 40 0 -1 1410
box -4 -6 36 206
use INVX1  _1473_
timestamp 1618002947
transform 1 0 40 0 -1 1410
box -4 -6 36 206
use NAND2X1  _1472_
timestamp 1618002947
transform -1 0 120 0 -1 1410
box -4 -6 52 206
use NOR2X1  _1468_
timestamp 1618002947
transform 1 0 120 0 -1 1410
box -4 -6 52 206
use OAI21X1  _1474_
timestamp 1618002947
transform 1 0 168 0 -1 1410
box -4 -6 68 206
use NAND3X1  _1537_
timestamp 1618002947
transform -1 0 296 0 -1 1410
box -4 -6 68 206
use NAND3X1  _1535_
timestamp 1618002947
transform -1 0 360 0 -1 1410
box -4 -6 68 206
use OAI21X1  _1536_
timestamp 1618002947
transform 1 0 360 0 -1 1410
box -4 -6 68 206
use NAND3X1  _1503_
timestamp 1618002947
transform -1 0 488 0 -1 1410
box -4 -6 68 206
use DFFSR  _1719_
timestamp 1618002947
transform -1 0 840 0 -1 1410
box -4 -6 356 206
use NOR2X1  _1306_
timestamp 1618002947
transform 1 0 840 0 -1 1410
box -4 -6 52 206
use INVX2  _1305_
timestamp 1618002947
transform -1 0 920 0 -1 1410
box -4 -6 36 206
use AOI21X1  _1449_
timestamp 1618002947
transform 1 0 920 0 -1 1410
box -4 -6 68 206
use DFFSR  _1714_
timestamp 1618002947
transform 1 0 984 0 -1 1410
box -4 -6 356 206
use INVX1  _1362_
timestamp 1618002947
transform -1 0 1432 0 -1 1410
box -4 -6 36 206
use OAI21X1  _1414_
timestamp 1618002947
transform 1 0 1432 0 -1 1410
box -4 -6 68 206
use FILL  SFILL13360x12100
timestamp 1618002947
transform -1 0 1352 0 -1 1410
box -4 -6 20 206
use FILL  SFILL13520x12100
timestamp 1618002947
transform -1 0 1368 0 -1 1410
box -4 -6 20 206
use FILL  SFILL13680x12100
timestamp 1618002947
transform -1 0 1384 0 -1 1410
box -4 -6 20 206
use FILL  SFILL13840x12100
timestamp 1618002947
transform -1 0 1400 0 -1 1410
box -4 -6 20 206
use AND2X2  _1415_
timestamp 1618002947
transform 1 0 1496 0 -1 1410
box -4 -6 68 206
use AND2X2  _1350_
timestamp 1618002947
transform -1 0 1624 0 -1 1410
box -4 -6 68 206
use NOR2X1  _1335_
timestamp 1618002947
transform -1 0 1672 0 -1 1410
box -4 -6 52 206
use OAI21X1  _1351_
timestamp 1618002947
transform 1 0 1672 0 -1 1410
box -4 -6 68 206
use NAND2X1  _1336_
timestamp 1618002947
transform -1 0 1784 0 -1 1410
box -4 -6 52 206
use INVX1  _1334_
timestamp 1618002947
transform -1 0 1816 0 -1 1410
box -4 -6 36 206
use DFFSR  _1688_
timestamp 1618002947
transform -1 0 2168 0 -1 1410
box -4 -6 356 206
use NOR2X1  _1345_
timestamp 1618002947
transform 1 0 2168 0 -1 1410
box -4 -6 52 206
use OAI21X1  _1344_
timestamp 1618002947
transform -1 0 2280 0 -1 1410
box -4 -6 68 206
use OAI21X1  _1369_
timestamp 1618002947
transform 1 0 2280 0 -1 1410
box -4 -6 68 206
use NAND3X1  _1343_
timestamp 1618002947
transform -1 0 2408 0 -1 1410
box -4 -6 68 206
use INVX1  _1331_
timestamp 1618002947
transform -1 0 2440 0 -1 1410
box -4 -6 36 206
use NAND2X1  _1348_
timestamp 1618002947
transform -1 0 2488 0 -1 1410
box -4 -6 52 206
use NOR2X1  _1349_
timestamp 1618002947
transform -1 0 2536 0 -1 1410
box -4 -6 52 206
use NOR2X1  _1342_
timestamp 1618002947
transform 1 0 2536 0 -1 1410
box -4 -6 52 206
use OAI21X1  _1385_
timestamp 1618002947
transform 1 0 2584 0 -1 1410
box -4 -6 68 206
use DFFSR  _1059_
timestamp 1618002947
transform -1 0 3064 0 -1 1410
box -4 -6 356 206
use FILL  SFILL26480x12100
timestamp 1618002947
transform -1 0 2664 0 -1 1410
box -4 -6 20 206
use FILL  SFILL26640x12100
timestamp 1618002947
transform -1 0 2680 0 -1 1410
box -4 -6 20 206
use FILL  SFILL26800x12100
timestamp 1618002947
transform -1 0 2696 0 -1 1410
box -4 -6 20 206
use FILL  SFILL26960x12100
timestamp 1618002947
transform -1 0 2712 0 -1 1410
box -4 -6 20 206
use OAI21X1  _1001_
timestamp 1618002947
transform -1 0 3128 0 -1 1410
box -4 -6 68 206
use INVX1  _999_
timestamp 1618002947
transform -1 0 3160 0 -1 1410
box -4 -6 36 206
use OAI21X1  _1000_
timestamp 1618002947
transform -1 0 3224 0 -1 1410
box -4 -6 68 206
use DFFSR  _1040_
timestamp 1618002947
transform 1 0 3224 0 -1 1410
box -4 -6 356 206
use INVX1  _898_
timestamp 1618002947
transform 1 0 3576 0 -1 1410
box -4 -6 36 206
use INVX1  _833_
timestamp 1618002947
transform 1 0 3608 0 -1 1410
box -4 -6 36 206
use OAI22X1  _941_
timestamp 1618002947
transform -1 0 3720 0 -1 1410
box -4 -6 84 206
use AOI21X1  _841_
timestamp 1618002947
transform 1 0 3720 0 -1 1410
box -4 -6 68 206
use NOR2X1  _840_
timestamp 1618002947
transform 1 0 3784 0 -1 1410
box -4 -6 52 206
use AOI22X1  _857_
timestamp 1618002947
transform 1 0 3832 0 -1 1410
box -4 -6 84 206
use INVX1  _844_
timestamp 1618002947
transform -1 0 3944 0 -1 1410
box -4 -6 36 206
use DFFSR  _1029_
timestamp 1618002947
transform -1 0 4296 0 -1 1410
box -4 -6 356 206
use FILL  SFILL42960x12100
timestamp 1618002947
transform -1 0 4312 0 -1 1410
box -4 -6 20 206
use FILL  SFILL43120x12100
timestamp 1618002947
transform -1 0 4328 0 -1 1410
box -4 -6 20 206
use FILL  SFILL43280x12100
timestamp 1618002947
transform -1 0 4344 0 -1 1410
box -4 -6 20 206
use NOR2X1  _851_
timestamp 1618002947
transform 1 0 4360 0 -1 1410
box -4 -6 52 206
use AOI21X1  _855_
timestamp 1618002947
transform 1 0 4408 0 -1 1410
box -4 -6 68 206
use NAND3X1  _858_
timestamp 1618002947
transform 1 0 4472 0 -1 1410
box -4 -6 68 206
use OAI22X1  _835_
timestamp 1618002947
transform 1 0 4536 0 -1 1410
box -4 -6 84 206
use INVX1  _834_
timestamp 1618002947
transform -1 0 4648 0 -1 1410
box -4 -6 36 206
use DFFSR  _1035_
timestamp 1618002947
transform 1 0 4648 0 -1 1410
box -4 -6 356 206
use FILL  SFILL43440x12100
timestamp 1618002947
transform -1 0 4360 0 -1 1410
box -4 -6 20 206
use MUX2X1  _1152_
timestamp 1618002947
transform 1 0 5000 0 -1 1410
box -4 -6 100 206
use NAND2X1  _1151_
timestamp 1618002947
transform 1 0 5096 0 -1 1410
box -4 -6 52 206
use DFFSR  _1037_
timestamp 1618002947
transform -1 0 5496 0 -1 1410
box -4 -6 356 206
use FILL  FILL53040x12100
timestamp 1618002947
transform -1 0 5512 0 -1 1410
box -4 -6 20 206
use BUFX2  _1752_
timestamp 1618002947
transform -1 0 56 0 1 1410
box -4 -6 52 206
use NAND3X1  _1288_
timestamp 1618002947
transform 1 0 56 0 1 1410
box -4 -6 68 206
use NOR3X1  _1471_
timestamp 1618002947
transform -1 0 248 0 1 1410
box -4 -6 132 206
use INVX1  _1469_
timestamp 1618002947
transform 1 0 248 0 1 1410
box -4 -6 36 206
use NOR2X1  _1266_
timestamp 1618002947
transform 1 0 280 0 1 1410
box -4 -6 52 206
use NOR2X1  _1289_
timestamp 1618002947
transform 1 0 328 0 1 1410
box -4 -6 52 206
use INVX1  _1467_
timestamp 1618002947
transform -1 0 408 0 1 1410
box -4 -6 36 206
use NAND2X1  _1294_
timestamp 1618002947
transform 1 0 408 0 1 1410
box -4 -6 52 206
use NOR3X1  _1502_
timestamp 1618002947
transform 1 0 456 0 1 1410
box -4 -6 132 206
use OAI21X1  _1534_
timestamp 1618002947
transform 1 0 584 0 1 1410
box -4 -6 68 206
use NAND2X1  _1533_
timestamp 1618002947
transform -1 0 696 0 1 1410
box -4 -6 52 206
use DFFSR  _1718_
timestamp 1618002947
transform -1 0 1048 0 1 1410
box -4 -6 356 206
use NOR2X1  _1450_
timestamp 1618002947
transform -1 0 1096 0 1 1410
box -4 -6 52 206
use INVX2  _1303_
timestamp 1618002947
transform 1 0 1096 0 1 1410
box -4 -6 36 206
use OAI21X1  _1448_
timestamp 1618002947
transform 1 0 1128 0 1 1410
box -4 -6 68 206
use INVX1  _1260_
timestamp 1618002947
transform 1 0 1192 0 1 1410
box -4 -6 36 206
use DFFPOSX1  _1677_
timestamp 1618002947
transform 1 0 1288 0 1 1410
box -4 -6 196 206
use FILL  SFILL12240x14100
timestamp 1618002947
transform 1 0 1224 0 1 1410
box -4 -6 20 206
use FILL  SFILL12400x14100
timestamp 1618002947
transform 1 0 1240 0 1 1410
box -4 -6 20 206
use FILL  SFILL12560x14100
timestamp 1618002947
transform 1 0 1256 0 1 1410
box -4 -6 20 206
use FILL  SFILL12720x14100
timestamp 1618002947
transform 1 0 1272 0 1 1410
box -4 -6 20 206
use DFFSR  _1689_
timestamp 1618002947
transform 1 0 1480 0 1 1410
box -4 -6 356 206
use OAI21X1  _1354_
timestamp 1618002947
transform 1 0 1832 0 1 1410
box -4 -6 68 206
use NAND2X1  _1355_
timestamp 1618002947
transform 1 0 1896 0 1 1410
box -4 -6 52 206
use AOI21X1  _1352_
timestamp 1618002947
transform -1 0 2008 0 1 1410
box -4 -6 68 206
use INVX1  _1346_
timestamp 1618002947
transform 1 0 2008 0 1 1410
box -4 -6 36 206
use NOR2X1  _1337_
timestamp 1618002947
transform -1 0 2088 0 1 1410
box -4 -6 52 206
use AND2X2  _1359_
timestamp 1618002947
transform 1 0 2088 0 1 1410
box -4 -6 68 206
use OAI21X1  _1360_
timestamp 1618002947
transform 1 0 2152 0 1 1410
box -4 -6 68 206
use DFFSR  _1697_
timestamp 1618002947
transform 1 0 2216 0 1 1410
box -4 -6 356 206
use NAND2X1  _1391_
timestamp 1618002947
transform -1 0 2616 0 1 1410
box -4 -6 52 206
use AOI21X1  _1388_
timestamp 1618002947
transform -1 0 2680 0 1 1410
box -4 -6 68 206
use NAND3X1  _1390_
timestamp 1618002947
transform 1 0 2680 0 1 1410
box -4 -6 68 206
use AND2X2  _1386_
timestamp 1618002947
transform 1 0 2808 0 1 1410
box -4 -6 68 206
use OAI21X1  _1387_
timestamp 1618002947
transform -1 0 2936 0 1 1410
box -4 -6 68 206
use FILL  SFILL27440x14100
timestamp 1618002947
transform 1 0 2744 0 1 1410
box -4 -6 20 206
use FILL  SFILL27600x14100
timestamp 1618002947
transform 1 0 2760 0 1 1410
box -4 -6 20 206
use FILL  SFILL27760x14100
timestamp 1618002947
transform 1 0 2776 0 1 1410
box -4 -6 20 206
use FILL  SFILL27920x14100
timestamp 1618002947
transform 1 0 2792 0 1 1410
box -4 -6 20 206
use DFFSR  _1058_
timestamp 1618002947
transform -1 0 3288 0 1 1410
box -4 -6 356 206
use OAI21X1  _998_
timestamp 1618002947
transform -1 0 3352 0 1 1410
box -4 -6 68 206
use INVX1  _996_
timestamp 1618002947
transform -1 0 3384 0 1 1410
box -4 -6 36 206
use OAI21X1  _997_
timestamp 1618002947
transform -1 0 3448 0 1 1410
box -4 -6 68 206
use OAI21X1  _977_
timestamp 1618002947
transform -1 0 3512 0 1 1410
box -4 -6 68 206
use OAI21X1  _968_
timestamp 1618002947
transform -1 0 3576 0 1 1410
box -4 -6 68 206
use OAI21X1  _965_
timestamp 1618002947
transform 1 0 3576 0 1 1410
box -4 -6 68 206
use NAND2X1  _911_
timestamp 1618002947
transform 1 0 3640 0 1 1410
box -4 -6 52 206
use AOI22X1  _848_
timestamp 1618002947
transform -1 0 3768 0 1 1410
box -4 -6 84 206
use MUX2X1  _912_
timestamp 1618002947
transform -1 0 3864 0 1 1410
box -4 -6 100 206
use INVX1  _910_
timestamp 1618002947
transform -1 0 3896 0 1 1410
box -4 -6 36 206
use AND2X2  _845_
timestamp 1618002947
transform -1 0 3960 0 1 1410
box -4 -6 68 206
use NAND3X1  _878_
timestamp 1618002947
transform -1 0 4024 0 1 1410
box -4 -6 68 206
use NAND3X1  _818_
timestamp 1618002947
transform -1 0 4088 0 1 1410
box -4 -6 68 206
use OAI21X1  _879_
timestamp 1618002947
transform -1 0 4152 0 1 1410
box -4 -6 68 206
use INVX1  _877_
timestamp 1618002947
transform 1 0 4152 0 1 1410
box -4 -6 36 206
use MUX2X1  _916_
timestamp 1618002947
transform 1 0 4184 0 1 1410
box -4 -6 100 206
use FILL  SFILL42800x14100
timestamp 1618002947
transform 1 0 4280 0 1 1410
box -4 -6 20 206
use FILL  SFILL42960x14100
timestamp 1618002947
transform 1 0 4296 0 1 1410
box -4 -6 20 206
use FILL  SFILL43120x14100
timestamp 1618002947
transform 1 0 4312 0 1 1410
box -4 -6 20 206
use FILL  SFILL43280x14100
timestamp 1618002947
transform 1 0 4328 0 1 1410
box -4 -6 20 206
use DFFPOSX1  _1012_
timestamp 1618002947
transform 1 0 4344 0 1 1410
box -4 -6 196 206
use NAND3X1  _813_
timestamp 1618002947
transform -1 0 4600 0 1 1410
box -4 -6 68 206
use NAND3X1  _822_
timestamp 1618002947
transform 1 0 4600 0 1 1410
box -4 -6 68 206
use NOR3X1  _838_
timestamp 1618002947
transform 1 0 4664 0 1 1410
box -4 -6 132 206
use MUX2X1  _932_
timestamp 1618002947
transform -1 0 4888 0 1 1410
box -4 -6 100 206
use INVX1  _931_
timestamp 1618002947
transform -1 0 4920 0 1 1410
box -4 -6 36 206
use OAI22X1  _872_
timestamp 1618002947
transform -1 0 5000 0 1 1410
box -4 -6 84 206
use MUX2X1  _935_
timestamp 1618002947
transform -1 0 5096 0 1 1410
box -4 -6 100 206
use INVX1  _864_
timestamp 1618002947
transform -1 0 5128 0 1 1410
box -4 -6 36 206
use INVX1  _870_
timestamp 1618002947
transform -1 0 5160 0 1 1410
box -4 -6 36 206
use MUX2X1  _1155_
timestamp 1618002947
transform 1 0 5160 0 1 1410
box -4 -6 100 206
use DFFPOSX1  _1014_
timestamp 1618002947
transform 1 0 5256 0 1 1410
box -4 -6 196 206
use BUFX2  _1758_
timestamp 1618002947
transform 1 0 5448 0 1 1410
box -4 -6 52 206
use FILL  FILL53040x14100
timestamp 1618002947
transform 1 0 5496 0 1 1410
box -4 -6 20 206
use INVX1  _1478_
timestamp 1618002947
transform 1 0 8 0 -1 1810
box -4 -6 36 206
use NOR2X1  _1481_
timestamp 1618002947
transform -1 0 88 0 -1 1810
box -4 -6 52 206
use NOR2X1  _1272_
timestamp 1618002947
transform 1 0 88 0 -1 1810
box -4 -6 52 206
use NOR2X1  _1477_
timestamp 1618002947
transform -1 0 184 0 -1 1810
box -4 -6 52 206
use INVX1  _1512_
timestamp 1618002947
transform 1 0 184 0 -1 1810
box -4 -6 36 206
use INVX1  _1479_
timestamp 1618002947
transform -1 0 248 0 -1 1810
box -4 -6 36 206
use NAND3X1  _1513_
timestamp 1618002947
transform -1 0 312 0 -1 1810
box -4 -6 68 206
use NAND3X1  _1514_
timestamp 1618002947
transform 1 0 312 0 -1 1810
box -4 -6 68 206
use OAI22X1  _1532_
timestamp 1618002947
transform 1 0 376 0 -1 1810
box -4 -6 84 206
use NAND2X1  _1482_
timestamp 1618002947
transform 1 0 456 0 -1 1810
box -4 -6 52 206
use NAND2X1  _1487_
timestamp 1618002947
transform -1 0 552 0 -1 1810
box -4 -6 52 206
use DFFSR  _1717_
timestamp 1618002947
transform -1 0 904 0 -1 1810
box -4 -6 356 206
use OAI21X1  _1578_
timestamp 1618002947
transform 1 0 904 0 -1 1810
box -4 -6 68 206
use NOR2X1  _1579_
timestamp 1618002947
transform -1 0 1016 0 -1 1810
box -4 -6 52 206
use AOI22X1  _1583_
timestamp 1618002947
transform -1 0 1096 0 -1 1810
box -4 -6 84 206
use DFFSR  _1734_
timestamp 1618002947
transform -1 0 1512 0 -1 1810
box -4 -6 356 206
use FILL  SFILL10960x16100
timestamp 1618002947
transform -1 0 1112 0 -1 1810
box -4 -6 20 206
use FILL  SFILL11120x16100
timestamp 1618002947
transform -1 0 1128 0 -1 1810
box -4 -6 20 206
use FILL  SFILL11280x16100
timestamp 1618002947
transform -1 0 1144 0 -1 1810
box -4 -6 20 206
use FILL  SFILL11440x16100
timestamp 1618002947
transform -1 0 1160 0 -1 1810
box -4 -6 20 206
use DFFSR  _1690_
timestamp 1618002947
transform 1 0 1512 0 -1 1810
box -4 -6 356 206
use NAND2X1  _1356_
timestamp 1618002947
transform 1 0 1864 0 -1 1810
box -4 -6 52 206
use AOI21X1  _1357_
timestamp 1618002947
transform -1 0 1976 0 -1 1810
box -4 -6 68 206
use INVX1  _1353_
timestamp 1618002947
transform -1 0 2008 0 -1 1810
box -4 -6 36 206
use DFFSR  _1691_
timestamp 1618002947
transform -1 0 2360 0 -1 1810
box -4 -6 356 206
use AOI21X1  _1361_
timestamp 1618002947
transform -1 0 2424 0 -1 1810
box -4 -6 68 206
use INVX1  _1358_
timestamp 1618002947
transform -1 0 2456 0 -1 1810
box -4 -6 36 206
use OAI21X1  _1393_
timestamp 1618002947
transform -1 0 2520 0 -1 1810
box -4 -6 68 206
use NAND2X1  _1406_
timestamp 1618002947
transform -1 0 2568 0 -1 1810
box -4 -6 52 206
use AOI21X1  _1394_
timestamp 1618002947
transform -1 0 2632 0 -1 1810
box -4 -6 68 206
use NAND3X1  _1401_
timestamp 1618002947
transform -1 0 2696 0 -1 1810
box -4 -6 68 206
use AOI21X1  _1403_
timestamp 1618002947
transform -1 0 2760 0 -1 1810
box -4 -6 68 206
use OAI21X1  _1400_
timestamp 1618002947
transform 1 0 2824 0 -1 1810
box -4 -6 68 206
use NOR2X1  _1328_
timestamp 1618002947
transform 1 0 2888 0 -1 1810
box -4 -6 52 206
use FILL  SFILL27600x16100
timestamp 1618002947
transform -1 0 2776 0 -1 1810
box -4 -6 20 206
use FILL  SFILL27760x16100
timestamp 1618002947
transform -1 0 2792 0 -1 1810
box -4 -6 20 206
use FILL  SFILL27920x16100
timestamp 1618002947
transform -1 0 2808 0 -1 1810
box -4 -6 20 206
use FILL  SFILL28080x16100
timestamp 1618002947
transform -1 0 2824 0 -1 1810
box -4 -6 20 206
use DFFSR  _1700_
timestamp 1618002947
transform -1 0 3288 0 -1 1810
box -4 -6 356 206
use NAND2X1  _1263_
timestamp 1618002947
transform -1 0 3336 0 -1 1810
box -4 -6 52 206
use INVX1  _973_
timestamp 1618002947
transform 1 0 3336 0 -1 1810
box -4 -6 36 206
use OAI21X1  _975_
timestamp 1618002947
transform 1 0 3368 0 -1 1810
box -4 -6 68 206
use OAI21X1  _974_
timestamp 1618002947
transform -1 0 3496 0 -1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert1
timestamp 1618002947
transform 1 0 3496 0 -1 1810
box -4 -6 52 206
use INVX1  _962_
timestamp 1618002947
transform -1 0 3576 0 -1 1810
box -4 -6 36 206
use OAI21X1  _966_
timestamp 1618002947
transform 1 0 3576 0 -1 1810
box -4 -6 68 206
use DFFSR  _1027_
timestamp 1618002947
transform 1 0 3640 0 -1 1810
box -4 -6 356 206
use NAND3X1  _831_
timestamp 1618002947
transform -1 0 4056 0 -1 1810
box -4 -6 68 206
use NOR2X1  _880_
timestamp 1618002947
transform -1 0 4104 0 -1 1810
box -4 -6 52 206
use DFFSR  _1030_
timestamp 1618002947
transform -1 0 4520 0 -1 1810
box -4 -6 356 206
use FILL  SFILL41040x16100
timestamp 1618002947
transform -1 0 4120 0 -1 1810
box -4 -6 20 206
use FILL  SFILL41200x16100
timestamp 1618002947
transform -1 0 4136 0 -1 1810
box -4 -6 20 206
use FILL  SFILL41360x16100
timestamp 1618002947
transform -1 0 4152 0 -1 1810
box -4 -6 20 206
use FILL  SFILL41520x16100
timestamp 1618002947
transform -1 0 4168 0 -1 1810
box -4 -6 20 206
use NOR2X1  _854_
timestamp 1618002947
transform -1 0 4568 0 -1 1810
box -4 -6 52 206
use INVX4  _805_
timestamp 1618002947
transform 1 0 4568 0 -1 1810
box -4 -6 52 206
use NOR2X1  _817_
timestamp 1618002947
transform -1 0 4664 0 -1 1810
box -4 -6 52 206
use NAND3X1  _811_
timestamp 1618002947
transform -1 0 4728 0 -1 1810
box -4 -6 68 206
use NAND3X1  _806_
timestamp 1618002947
transform -1 0 4792 0 -1 1810
box -4 -6 68 206
use INVX2  _812_
timestamp 1618002947
transform -1 0 4824 0 -1 1810
box -4 -6 36 206
use NAND3X1  _821_
timestamp 1618002947
transform 1 0 4824 0 -1 1810
box -4 -6 68 206
use INVX1  _810_
timestamp 1618002947
transform -1 0 4920 0 -1 1810
box -4 -6 36 206
use NAND3X1  _819_
timestamp 1618002947
transform -1 0 4984 0 -1 1810
box -4 -6 68 206
use INVX2  _807_
timestamp 1618002947
transform 1 0 4984 0 -1 1810
box -4 -6 36 206
use AOI21X1  _873_
timestamp 1618002947
transform -1 0 5080 0 -1 1810
box -4 -6 68 206
use NAND2X1  _881_
timestamp 1618002947
transform 1 0 5080 0 -1 1810
box -4 -6 52 206
use DFFSR  _1038_
timestamp 1618002947
transform -1 0 5480 0 -1 1810
box -4 -6 356 206
use FILL  FILL52880x16100
timestamp 1618002947
transform -1 0 5496 0 -1 1810
box -4 -6 20 206
use FILL  FILL53040x16100
timestamp 1618002947
transform -1 0 5512 0 -1 1810
box -4 -6 20 206
use NAND2X1  _1268_
timestamp 1618002947
transform 1 0 8 0 1 1810
box -4 -6 52 206
use NAND2X1  _1480_
timestamp 1618002947
transform -1 0 104 0 1 1810
box -4 -6 52 206
use NOR2X1  _1485_
timestamp 1618002947
transform -1 0 152 0 1 1810
box -4 -6 52 206
use AND2X2  _1486_
timestamp 1618002947
transform 1 0 152 0 1 1810
box -4 -6 68 206
use NOR2X1  _1267_
timestamp 1618002947
transform 1 0 216 0 1 1810
box -4 -6 52 206
use OR2X2  _1520_
timestamp 1618002947
transform 1 0 264 0 1 1810
box -4 -6 68 206
use NAND3X1  _1515_
timestamp 1618002947
transform 1 0 328 0 1 1810
box -4 -6 68 206
use NAND3X1  _1511_
timestamp 1618002947
transform -1 0 456 0 1 1810
box -4 -6 68 206
use INVX1  _1476_
timestamp 1618002947
transform 1 0 456 0 1 1810
box -4 -6 36 206
use NAND2X1  _1542_
timestamp 1618002947
transform 1 0 488 0 1 1810
box -4 -6 52 206
use NAND3X1  _1488_
timestamp 1618002947
transform -1 0 600 0 1 1810
box -4 -6 68 206
use AND2X2  _1307_
timestamp 1618002947
transform 1 0 600 0 1 1810
box -4 -6 68 206
use DFFSR  _1679_
timestamp 1618002947
transform 1 0 664 0 1 1810
box -4 -6 356 206
use DFFSR  _1706_
timestamp 1618002947
transform -1 0 1368 0 1 1810
box -4 -6 356 206
use DFFSR  _1707_
timestamp 1618002947
transform 1 0 1432 0 1 1810
box -4 -6 356 206
use FILL  SFILL13680x18100
timestamp 1618002947
transform 1 0 1368 0 1 1810
box -4 -6 20 206
use FILL  SFILL13840x18100
timestamp 1618002947
transform 1 0 1384 0 1 1810
box -4 -6 20 206
use FILL  SFILL14000x18100
timestamp 1618002947
transform 1 0 1400 0 1 1810
box -4 -6 20 206
use FILL  SFILL14160x18100
timestamp 1618002947
transform 1 0 1416 0 1 1810
box -4 -6 20 206
use INVX2  _1327_
timestamp 1618002947
transform -1 0 1816 0 1 1810
box -4 -6 36 206
use DFFSR  _1744_
timestamp 1618002947
transform -1 0 2168 0 1 1810
box -4 -6 356 206
use INVX1  _1389_
timestamp 1618002947
transform -1 0 2200 0 1 1810
box -4 -6 36 206
use NAND3X1  _1397_
timestamp 1618002947
transform -1 0 2264 0 1 1810
box -4 -6 68 206
use INVX1  _1396_
timestamp 1618002947
transform -1 0 2296 0 1 1810
box -4 -6 36 206
use NAND2X1  _1392_
timestamp 1618002947
transform 1 0 2296 0 1 1810
box -4 -6 52 206
use NOR2X1  _1329_
timestamp 1618002947
transform -1 0 2392 0 1 1810
box -4 -6 52 206
use NAND2X1  _1330_
timestamp 1618002947
transform -1 0 2440 0 1 1810
box -4 -6 52 206
use INVX1  _1404_
timestamp 1618002947
transform 1 0 2440 0 1 1810
box -4 -6 36 206
use OAI21X1  _1405_
timestamp 1618002947
transform 1 0 2472 0 1 1810
box -4 -6 68 206
use AOI21X1  _1407_
timestamp 1618002947
transform 1 0 2536 0 1 1810
box -4 -6 68 206
use DFFSR  _1701_
timestamp 1618002947
transform -1 0 3016 0 1 1810
box -4 -6 356 206
use FILL  SFILL26000x18100
timestamp 1618002947
transform 1 0 2600 0 1 1810
box -4 -6 20 206
use FILL  SFILL26160x18100
timestamp 1618002947
transform 1 0 2616 0 1 1810
box -4 -6 20 206
use FILL  SFILL26320x18100
timestamp 1618002947
transform 1 0 2632 0 1 1810
box -4 -6 20 206
use FILL  SFILL26480x18100
timestamp 1618002947
transform 1 0 2648 0 1 1810
box -4 -6 20 206
use DFFSR  _1050_
timestamp 1618002947
transform -1 0 3368 0 1 1810
box -4 -6 356 206
use INVX1  _976_
timestamp 1618002947
transform 1 0 3368 0 1 1810
box -4 -6 36 206
use OAI21X1  _978_
timestamp 1618002947
transform 1 0 3400 0 1 1810
box -4 -6 68 206
use DFFSR  _1051_
timestamp 1618002947
transform 1 0 3464 0 1 1810
box -4 -6 356 206
use OAI21X1  _964_
timestamp 1618002947
transform -1 0 3880 0 1 1810
box -4 -6 68 206
use NAND3X1  _860_
timestamp 1618002947
transform 1 0 3880 0 1 1810
box -4 -6 68 206
use NAND2X1  _963_
timestamp 1618002947
transform -1 0 3992 0 1 1810
box -4 -6 52 206
use OAI21X1  _897_
timestamp 1618002947
transform 1 0 3992 0 1 1810
box -4 -6 68 206
use NAND3X1  _939_
timestamp 1618002947
transform 1 0 4088 0 1 1810
box -4 -6 68 206
use INVX1  _959_
timestamp 1618002947
transform 1 0 4056 0 1 1810
box -4 -6 36 206
use OAI21X1  _938_
timestamp 1618002947
transform 1 0 4184 0 1 1810
box -4 -6 68 206
use INVX1  _882_
timestamp 1618002947
transform -1 0 4184 0 1 1810
box -4 -6 36 206
use FILL  SFILL42480x18100
timestamp 1618002947
transform 1 0 4248 0 1 1810
box -4 -6 20 206
use FILL  SFILL42960x18100
timestamp 1618002947
transform 1 0 4296 0 1 1810
box -4 -6 20 206
use FILL  SFILL42800x18100
timestamp 1618002947
transform 1 0 4280 0 1 1810
box -4 -6 20 206
use FILL  SFILL42640x18100
timestamp 1618002947
transform 1 0 4264 0 1 1810
box -4 -6 20 206
use INVX1  _883_
timestamp 1618002947
transform -1 0 4344 0 1 1810
box -4 -6 36 206
use MUX2X1  _918_
timestamp 1618002947
transform 1 0 4344 0 1 1810
box -4 -6 100 206
use NAND3X1  _944_
timestamp 1618002947
transform -1 0 4504 0 1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert22
timestamp 1618002947
transform 1 0 4504 0 1 1810
box -4 -6 52 206
use NAND3X1  _888_
timestamp 1618002947
transform -1 0 4616 0 1 1810
box -4 -6 68 206
use OAI21X1  _889_
timestamp 1618002947
transform -1 0 4680 0 1 1810
box -4 -6 68 206
use DFFSR  _1028_
timestamp 1618002947
transform -1 0 5032 0 1 1810
box -4 -6 356 206
use OAI22X1  _865_
timestamp 1618002947
transform 1 0 5032 0 1 1810
box -4 -6 84 206
use MUX2X1  _1157_
timestamp 1618002947
transform 1 0 5112 0 1 1810
box -4 -6 100 206
use DFFPOSX1  _1016_
timestamp 1618002947
transform 1 0 5208 0 1 1810
box -4 -6 196 206
use OAI21X1  _1156_
timestamp 1618002947
transform 1 0 5400 0 1 1810
box -4 -6 68 206
use NAND2X1  _1154_
timestamp 1618002947
transform -1 0 5512 0 1 1810
box -4 -6 52 206
use INVX4  _1279_
timestamp 1618002947
transform -1 0 56 0 -1 2210
box -4 -6 52 206
use NOR2X1  _1286_
timestamp 1618002947
transform 1 0 56 0 -1 2210
box -4 -6 52 206
use AOI22X1  _1287_
timestamp 1618002947
transform 1 0 104 0 -1 2210
box -4 -6 84 206
use NAND2X1  _1285_
timestamp 1618002947
transform -1 0 232 0 -1 2210
box -4 -6 52 206
use NAND3X1  _1508_
timestamp 1618002947
transform -1 0 296 0 -1 2210
box -4 -6 68 206
use AND2X2  _1276_
timestamp 1618002947
transform 1 0 296 0 -1 2210
box -4 -6 68 206
use AND2X2  _1510_
timestamp 1618002947
transform 1 0 360 0 -1 2210
box -4 -6 68 206
use NAND3X1  _1475_
timestamp 1618002947
transform -1 0 488 0 -1 2210
box -4 -6 68 206
use NOR3X1  _1521_
timestamp 1618002947
transform 1 0 488 0 -1 2210
box -4 -6 132 206
use NAND3X1  _1302_
timestamp 1618002947
transform 1 0 616 0 -1 2210
box -4 -6 68 206
use NAND3X1  _1582_
timestamp 1618002947
transform 1 0 680 0 -1 2210
box -4 -6 68 206
use NAND3X1  _1573_
timestamp 1618002947
transform 1 0 744 0 -1 2210
box -4 -6 68 206
use OR2X2  _1574_
timestamp 1618002947
transform 1 0 808 0 -1 2210
box -4 -6 68 206
use NAND2X1  _1301_
timestamp 1618002947
transform -1 0 920 0 -1 2210
box -4 -6 52 206
use AOI21X1  _1572_
timestamp 1618002947
transform 1 0 920 0 -1 2210
box -4 -6 68 206
use NAND2X1  _1546_
timestamp 1618002947
transform 1 0 984 0 -1 2210
box -4 -6 52 206
use OAI21X1  _1547_
timestamp 1618002947
transform 1 0 1032 0 -1 2210
box -4 -6 68 206
use DFFSR  _1745_
timestamp 1618002947
transform 1 0 1160 0 -1 2210
box -4 -6 356 206
use FILL  SFILL10960x20100
timestamp 1618002947
transform -1 0 1112 0 -1 2210
box -4 -6 20 206
use FILL  SFILL11120x20100
timestamp 1618002947
transform -1 0 1128 0 -1 2210
box -4 -6 20 206
use FILL  SFILL11280x20100
timestamp 1618002947
transform -1 0 1144 0 -1 2210
box -4 -6 20 206
use FILL  SFILL11440x20100
timestamp 1618002947
transform -1 0 1160 0 -1 2210
box -4 -6 20 206
use NOR2X1  _1254_
timestamp 1618002947
transform -1 0 1560 0 -1 2210
box -4 -6 52 206
use NAND2X1  _1647_
timestamp 1618002947
transform 1 0 1560 0 -1 2210
box -4 -6 52 206
use OAI21X1  _1643_
timestamp 1618002947
transform 1 0 1608 0 -1 2210
box -4 -6 68 206
use AOI22X1  _1646_
timestamp 1618002947
transform -1 0 1752 0 -1 2210
box -4 -6 84 206
use INVX1  _1413_
timestamp 1618002947
transform -1 0 1784 0 -1 2210
box -4 -6 36 206
use AND2X2  _1637_
timestamp 1618002947
transform 1 0 1784 0 -1 2210
box -4 -6 68 206
use NOR2X1  _1636_
timestamp 1618002947
transform -1 0 1896 0 -1 2210
box -4 -6 52 206
use OAI21X1  _1638_
timestamp 1618002947
transform 1 0 1896 0 -1 2210
box -4 -6 68 206
use NAND2X1  _1639_
timestamp 1618002947
transform 1 0 1960 0 -1 2210
box -4 -6 52 206
use NAND3X1  _1641_
timestamp 1618002947
transform -1 0 2072 0 -1 2210
box -4 -6 68 206
use AOI22X1  _1627_
timestamp 1618002947
transform -1 0 2152 0 -1 2210
box -4 -6 84 206
use NAND2X1  _1640_
timestamp 1618002947
transform -1 0 2200 0 -1 2210
box -4 -6 52 206
use OAI21X1  _1402_
timestamp 1618002947
transform 1 0 2200 0 -1 2210
box -4 -6 68 206
use OAI21X1  _1395_
timestamp 1618002947
transform 1 0 2264 0 -1 2210
box -4 -6 68 206
use AOI21X1  _1399_
timestamp 1618002947
transform 1 0 2328 0 -1 2210
box -4 -6 68 206
use OAI21X1  _1398_
timestamp 1618002947
transform -1 0 2456 0 -1 2210
box -4 -6 68 206
use DFFSR  _1699_
timestamp 1618002947
transform -1 0 2808 0 -1 2210
box -4 -6 356 206
use INVX1  _875_
timestamp 1618002947
transform 1 0 2872 0 -1 2210
box -4 -6 36 206
use FILL  SFILL28080x20100
timestamp 1618002947
transform -1 0 2824 0 -1 2210
box -4 -6 20 206
use FILL  SFILL28240x20100
timestamp 1618002947
transform -1 0 2840 0 -1 2210
box -4 -6 20 206
use FILL  SFILL28400x20100
timestamp 1618002947
transform -1 0 2856 0 -1 2210
box -4 -6 20 206
use FILL  SFILL28560x20100
timestamp 1618002947
transform -1 0 2872 0 -1 2210
box -4 -6 20 206
use DFFSR  _1054_
timestamp 1618002947
transform -1 0 3256 0 -1 2210
box -4 -6 356 206
use INVX1  _985_
timestamp 1618002947
transform 1 0 3256 0 -1 2210
box -4 -6 36 206
use OAI21X1  _987_
timestamp 1618002947
transform 1 0 3288 0 -1 2210
box -4 -6 68 206
use OAI21X1  _986_
timestamp 1618002947
transform -1 0 3416 0 -1 2210
box -4 -6 68 206
use INVX1  _884_
timestamp 1618002947
transform 1 0 3416 0 -1 2210
box -4 -6 36 206
use DFFPOSX1  _1017_
timestamp 1618002947
transform -1 0 3640 0 -1 2210
box -4 -6 196 206
use OAI21X1  _988_
timestamp 1618002947
transform -1 0 3704 0 -1 2210
box -4 -6 68 206
use OAI22X1  _885_
timestamp 1618002947
transform -1 0 3784 0 -1 2210
box -4 -6 84 206
use AOI21X1  _886_
timestamp 1618002947
transform -1 0 3848 0 -1 2210
box -4 -6 68 206
use NAND2X1  _893_
timestamp 1618002947
transform 1 0 3848 0 -1 2210
box -4 -6 52 206
use OAI21X1  _861_
timestamp 1618002947
transform 1 0 3896 0 -1 2210
box -4 -6 68 206
use OAI22X1  _876_
timestamp 1618002947
transform -1 0 4040 0 -1 2210
box -4 -6 84 206
use OAI22X1  _961_
timestamp 1618002947
transform -1 0 4120 0 -1 2210
box -4 -6 84 206
use NOR2X1  _937_
timestamp 1618002947
transform -1 0 4168 0 -1 2210
box -4 -6 52 206
use OAI21X1  _960_
timestamp 1618002947
transform -1 0 4232 0 -1 2210
box -4 -6 68 206
use AOI22X1  _945_
timestamp 1618002947
transform -1 0 4376 0 -1 2210
box -4 -6 84 206
use FILL  SFILL42320x20100
timestamp 1618002947
transform -1 0 4248 0 -1 2210
box -4 -6 20 206
use FILL  SFILL42480x20100
timestamp 1618002947
transform -1 0 4264 0 -1 2210
box -4 -6 20 206
use FILL  SFILL42640x20100
timestamp 1618002947
transform -1 0 4280 0 -1 2210
box -4 -6 20 206
use FILL  SFILL42800x20100
timestamp 1618002947
transform -1 0 4296 0 -1 2210
box -4 -6 20 206
use NOR2X1  _956_
timestamp 1618002947
transform 1 0 4376 0 -1 2210
box -4 -6 52 206
use NOR2X1  _892_
timestamp 1618002947
transform -1 0 4472 0 -1 2210
box -4 -6 52 206
use OAI22X1  _891_
timestamp 1618002947
transform -1 0 4552 0 -1 2210
box -4 -6 84 206
use OAI22X1  _867_
timestamp 1618002947
transform 1 0 4552 0 -1 2210
box -4 -6 84 206
use MUX2X1  _914_
timestamp 1618002947
transform 1 0 4632 0 -1 2210
box -4 -6 100 206
use OAI21X1  _919_
timestamp 1618002947
transform 1 0 4728 0 -1 2210
box -4 -6 68 206
use DFFSR  _1036_
timestamp 1618002947
transform -1 0 5144 0 -1 2210
box -4 -6 356 206
use DFFSR  _1235_
timestamp 1618002947
transform 1 0 5144 0 -1 2210
box -4 -6 356 206
use FILL  FILL53040x20100
timestamp 1618002947
transform -1 0 5512 0 -1 2210
box -4 -6 20 206
use DFFSR  _1732_
timestamp 1618002947
transform -1 0 360 0 1 2210
box -4 -6 356 206
use NAND3X1  _1509_
timestamp 1618002947
transform 1 0 360 0 1 2210
box -4 -6 68 206
use OAI22X1  _1569_
timestamp 1618002947
transform 1 0 424 0 1 2210
box -4 -6 84 206
use NOR2X1  _1309_
timestamp 1618002947
transform -1 0 552 0 1 2210
box -4 -6 52 206
use AND2X2  _1275_
timestamp 1618002947
transform -1 0 616 0 1 2210
box -4 -6 68 206
use NAND2X1  _1308_
timestamp 1618002947
transform -1 0 664 0 1 2210
box -4 -6 52 206
use NAND3X1  _1484_
timestamp 1618002947
transform -1 0 728 0 1 2210
box -4 -6 68 206
use AND2X2  _1298_
timestamp 1618002947
transform 1 0 728 0 1 2210
box -4 -6 68 206
use AOI21X1  _1581_
timestamp 1618002947
transform -1 0 856 0 1 2210
box -4 -6 68 206
use NOR2X1  _1483_
timestamp 1618002947
transform 1 0 856 0 1 2210
box -4 -6 52 206
use AND2X2  _1300_
timestamp 1618002947
transform 1 0 904 0 1 2210
box -4 -6 68 206
use AOI21X1  _1575_
timestamp 1618002947
transform -1 0 1032 0 1 2210
box -4 -6 68 206
use DFFSR  _1724_
timestamp 1618002947
transform -1 0 1384 0 1 2210
box -4 -6 356 206
use INVX4  _1587_
timestamp 1618002947
transform 1 0 1448 0 1 2210
box -4 -6 52 206
use FILL  SFILL13840x22100
timestamp 1618002947
transform 1 0 1384 0 1 2210
box -4 -6 20 206
use FILL  SFILL14000x22100
timestamp 1618002947
transform 1 0 1400 0 1 2210
box -4 -6 20 206
use FILL  SFILL14160x22100
timestamp 1618002947
transform 1 0 1416 0 1 2210
box -4 -6 20 206
use FILL  SFILL14320x22100
timestamp 1618002947
transform 1 0 1432 0 1 2210
box -4 -6 20 206
use INVX1  _1642_
timestamp 1618002947
transform -1 0 1528 0 1 2210
box -4 -6 36 206
use OAI21X1  _1645_
timestamp 1618002947
transform -1 0 1592 0 1 2210
box -4 -6 68 206
use OAI21X1  _1644_
timestamp 1618002947
transform 1 0 1592 0 1 2210
box -4 -6 68 206
use NAND2X1  _1265_
timestamp 1618002947
transform -1 0 1704 0 1 2210
box -4 -6 52 206
use AND2X2  _1585_
timestamp 1618002947
transform 1 0 1704 0 1 2210
box -4 -6 68 206
use NAND2X1  _1586_
timestamp 1618002947
transform 1 0 1768 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert26
timestamp 1618002947
transform -1 0 1864 0 1 2210
box -4 -6 52 206
use NAND2X1  _1626_
timestamp 1618002947
transform 1 0 1864 0 1 2210
box -4 -6 52 206
use OAI21X1  _1671_
timestamp 1618002947
transform -1 0 1976 0 1 2210
box -4 -6 68 206
use OAI21X1  _1628_
timestamp 1618002947
transform 1 0 1976 0 1 2210
box -4 -6 68 206
use DFFSR  _1742_
timestamp 1618002947
transform -1 0 2392 0 1 2210
box -4 -6 356 206
use DFFSR  _1698_
timestamp 1618002947
transform -1 0 2744 0 1 2210
box -4 -6 356 206
use INVX1  _859_
timestamp 1618002947
transform 1 0 2808 0 1 2210
box -4 -6 36 206
use DFFSR  _1061_
timestamp 1618002947
transform -1 0 3192 0 1 2210
box -4 -6 356 206
use FILL  SFILL27440x22100
timestamp 1618002947
transform 1 0 2744 0 1 2210
box -4 -6 20 206
use FILL  SFILL27600x22100
timestamp 1618002947
transform 1 0 2760 0 1 2210
box -4 -6 20 206
use FILL  SFILL27760x22100
timestamp 1618002947
transform 1 0 2776 0 1 2210
box -4 -6 20 206
use FILL  SFILL27920x22100
timestamp 1618002947
transform 1 0 2792 0 1 2210
box -4 -6 20 206
use OAI21X1  _1003_
timestamp 1618002947
transform 1 0 3192 0 1 2210
box -4 -6 68 206
use OAI21X1  _1005_
timestamp 1618002947
transform 1 0 3256 0 1 2210
box -4 -6 68 206
use OAI21X1  _1002_
timestamp 1618002947
transform -1 0 3384 0 1 2210
box -4 -6 68 206
use OAI21X1  _1004_
timestamp 1618002947
transform -1 0 3448 0 1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert2
timestamp 1618002947
transform -1 0 3496 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert0
timestamp 1618002947
transform 1 0 3496 0 1 2210
box -4 -6 52 206
use OAI21X1  _1007_
timestamp 1618002947
transform 1 0 3544 0 1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert20
timestamp 1618002947
transform -1 0 3656 0 1 2210
box -4 -6 52 206
use OAI21X1  _1006_
timestamp 1618002947
transform -1 0 3720 0 1 2210
box -4 -6 68 206
use NAND2X1  _915_
timestamp 1618002947
transform 1 0 3720 0 1 2210
box -4 -6 52 206
use DFFSR  _1044_
timestamp 1618002947
transform -1 0 4120 0 1 2210
box -4 -6 356 206
use INVX1  _874_
timestamp 1618002947
transform 1 0 4120 0 1 2210
box -4 -6 36 206
use OAI21X1  _955_
timestamp 1618002947
transform 1 0 4152 0 1 2210
box -4 -6 68 206
use NAND3X1  _954_
timestamp 1618002947
transform 1 0 4280 0 1 2210
box -4 -6 68 206
use FILL  SFILL42160x22100
timestamp 1618002947
transform 1 0 4216 0 1 2210
box -4 -6 20 206
use FILL  SFILL42320x22100
timestamp 1618002947
transform 1 0 4232 0 1 2210
box -4 -6 20 206
use FILL  SFILL42480x22100
timestamp 1618002947
transform 1 0 4248 0 1 2210
box -4 -6 20 206
use FILL  SFILL42640x22100
timestamp 1618002947
transform 1 0 4264 0 1 2210
box -4 -6 20 206
use NOR2X1  _953_
timestamp 1618002947
transform -1 0 4392 0 1 2210
box -4 -6 52 206
use NAND3X1  _957_
timestamp 1618002947
transform 1 0 4392 0 1 2210
box -4 -6 68 206
use NAND2X1  _946_
timestamp 1618002947
transform 1 0 4456 0 1 2210
box -4 -6 52 206
use OAI21X1  _949_
timestamp 1618002947
transform 1 0 4504 0 1 2210
box -4 -6 68 206
use NAND3X1  _948_
timestamp 1618002947
transform 1 0 4568 0 1 2210
box -4 -6 68 206
use NAND3X1  _951_
timestamp 1618002947
transform 1 0 4632 0 1 2210
box -4 -6 68 206
use NOR2X1  _947_
timestamp 1618002947
transform 1 0 4696 0 1 2210
box -4 -6 52 206
use NOR2X1  _950_
timestamp 1618002947
transform 1 0 4744 0 1 2210
box -4 -6 52 206
use AOI21X1  _800_
timestamp 1618002947
transform 1 0 4792 0 1 2210
box -4 -6 68 206
use NAND2X1  _913_
timestamp 1618002947
transform 1 0 4856 0 1 2210
box -4 -6 52 206
use NAND2X1  _917_
timestamp 1618002947
transform -1 0 4952 0 1 2210
box -4 -6 52 206
use DFFSR  _1021_
timestamp 1618002947
transform -1 0 5304 0 1 2210
box -4 -6 356 206
use AOI21X1  _943_
timestamp 1618002947
transform -1 0 5368 0 1 2210
box -4 -6 68 206
use NAND2X1  _896_
timestamp 1618002947
transform -1 0 5416 0 1 2210
box -4 -6 52 206
use NOR2X1  _895_
timestamp 1618002947
transform 1 0 5416 0 1 2210
box -4 -6 52 206
use BUFX2  _1755_
timestamp 1618002947
transform 1 0 5464 0 1 2210
box -4 -6 52 206
use INVX1  _1278_
timestamp 1618002947
transform 1 0 8 0 -1 2610
box -4 -6 36 206
use NOR2X1  _1282_
timestamp 1618002947
transform 1 0 40 0 -1 2610
box -4 -6 52 206
use NAND2X1  _1295_
timestamp 1618002947
transform 1 0 88 0 -1 2610
box -4 -6 52 206
use AND2X2  _1284_
timestamp 1618002947
transform 1 0 136 0 -1 2610
box -4 -6 68 206
use NOR2X1  _1465_
timestamp 1618002947
transform -1 0 248 0 -1 2610
box -4 -6 52 206
use AND2X2  _1564_
timestamp 1618002947
transform 1 0 248 0 -1 2610
box -4 -6 68 206
use OAI21X1  _1466_
timestamp 1618002947
transform 1 0 312 0 -1 2610
box -4 -6 68 206
use NOR2X1  _1297_
timestamp 1618002947
transform -1 0 424 0 -1 2610
box -4 -6 52 206
use NAND2X1  _1296_
timestamp 1618002947
transform 1 0 424 0 -1 2610
box -4 -6 52 206
use NAND3X1  _1571_
timestamp 1618002947
transform 1 0 472 0 -1 2610
box -4 -6 68 206
use NAND2X1  _1454_
timestamp 1618002947
transform 1 0 536 0 -1 2610
box -4 -6 52 206
use NAND2X1  _1554_
timestamp 1618002947
transform -1 0 632 0 -1 2610
box -4 -6 52 206
use NOR2X1  _1273_
timestamp 1618002947
transform 1 0 632 0 -1 2610
box -4 -6 52 206
use OAI21X1  _1555_
timestamp 1618002947
transform -1 0 744 0 -1 2610
box -4 -6 68 206
use NOR2X1  _1274_
timestamp 1618002947
transform 1 0 744 0 -1 2610
box -4 -6 52 206
use DFFSR  _1726_
timestamp 1618002947
transform -1 0 1144 0 -1 2610
box -4 -6 356 206
use NOR3X1  _1650_
timestamp 1618002947
transform -1 0 1272 0 -1 2610
box -4 -6 132 206
use AOI22X1  _1652_
timestamp 1618002947
transform -1 0 1416 0 -1 2610
box -4 -6 84 206
use INVX1  _1648_
timestamp 1618002947
transform -1 0 1448 0 -1 2610
box -4 -6 36 206
use DFFSR  _1741_
timestamp 1618002947
transform 1 0 1448 0 -1 2610
box -4 -6 356 206
use FILL  SFILL12720x24100
timestamp 1618002947
transform -1 0 1288 0 -1 2610
box -4 -6 20 206
use FILL  SFILL12880x24100
timestamp 1618002947
transform -1 0 1304 0 -1 2610
box -4 -6 20 206
use FILL  SFILL13040x24100
timestamp 1618002947
transform -1 0 1320 0 -1 2610
box -4 -6 20 206
use FILL  SFILL13200x24100
timestamp 1618002947
transform -1 0 1336 0 -1 2610
box -4 -6 20 206
use INVX4  _1592_
timestamp 1618002947
transform -1 0 1848 0 -1 2610
box -4 -6 52 206
use NAND2X1  _1588_
timestamp 1618002947
transform 1 0 1848 0 -1 2610
box -4 -6 52 206
use INVX1  _1619_
timestamp 1618002947
transform -1 0 1928 0 -1 2610
box -4 -6 36 206
use OAI21X1  _1618_
timestamp 1618002947
transform -1 0 1992 0 -1 2610
box -4 -6 68 206
use OR2X2  _1614_
timestamp 1618002947
transform 1 0 1992 0 -1 2610
box -4 -6 68 206
use DFFSR  _1740_
timestamp 1618002947
transform -1 0 2408 0 -1 2610
box -4 -6 356 206
use NAND2X1  _1674_
timestamp 1618002947
transform -1 0 2456 0 -1 2610
box -4 -6 52 206
use DFFSR  _1062_
timestamp 1618002947
transform -1 0 2808 0 -1 2610
box -4 -6 356 206
use DFFSR  _1047_
timestamp 1618002947
transform -1 0 3224 0 -1 2610
box -4 -6 356 206
use FILL  SFILL28080x24100
timestamp 1618002947
transform -1 0 2824 0 -1 2610
box -4 -6 20 206
use FILL  SFILL28240x24100
timestamp 1618002947
transform -1 0 2840 0 -1 2610
box -4 -6 20 206
use FILL  SFILL28400x24100
timestamp 1618002947
transform -1 0 2856 0 -1 2610
box -4 -6 20 206
use FILL  SFILL28560x24100
timestamp 1618002947
transform -1 0 2872 0 -1 2610
box -4 -6 20 206
use OAI21X1  _981_
timestamp 1618002947
transform -1 0 3288 0 -1 2610
box -4 -6 68 206
use OAI21X1  _980_
timestamp 1618002947
transform -1 0 3352 0 -1 2610
box -4 -6 68 206
use INVX4  _794_
timestamp 1618002947
transform -1 0 3400 0 -1 2610
box -4 -6 52 206
use INVX1  _967_
timestamp 1618002947
transform 1 0 3400 0 -1 2610
box -4 -6 36 206
use OAI21X1  _969_
timestamp 1618002947
transform 1 0 3432 0 -1 2610
box -4 -6 68 206
use DFFSR  _1020_
timestamp 1618002947
transform 1 0 3496 0 -1 2610
box -4 -6 356 206
use INVX1  _850_
timestamp 1618002947
transform -1 0 3880 0 -1 2610
box -4 -6 36 206
use DFFSR  _1046_
timestamp 1618002947
transform -1 0 4232 0 -1 2610
box -4 -6 356 206
use INVX1  _799_
timestamp 1618002947
transform 1 0 4296 0 -1 2610
box -4 -6 36 206
use DFFSR  _1042_
timestamp 1618002947
transform -1 0 4680 0 -1 2610
box -4 -6 356 206
use FILL  SFILL42320x24100
timestamp 1618002947
transform -1 0 4248 0 -1 2610
box -4 -6 20 206
use FILL  SFILL42480x24100
timestamp 1618002947
transform -1 0 4264 0 -1 2610
box -4 -6 20 206
use FILL  SFILL42640x24100
timestamp 1618002947
transform -1 0 4280 0 -1 2610
box -4 -6 20 206
use FILL  SFILL42800x24100
timestamp 1618002947
transform -1 0 4296 0 -1 2610
box -4 -6 20 206
use AOI21X1  _803_
timestamp 1618002947
transform -1 0 4744 0 -1 2610
box -4 -6 68 206
use NOR2X1  _804_
timestamp 1618002947
transform -1 0 4792 0 -1 2610
box -4 -6 52 206
use DFFSR  _1023_
timestamp 1618002947
transform 1 0 4792 0 -1 2610
box -4 -6 356 206
use CLKBUF1  CLKBUF1_insert8
timestamp 1618002947
transform 1 0 5144 0 -1 2610
box -4 -6 148 206
use DFFPOSX1  _1018_
timestamp 1618002947
transform -1 0 5480 0 -1 2610
box -4 -6 196 206
use FILL  FILL52880x24100
timestamp 1618002947
transform -1 0 5496 0 -1 2610
box -4 -6 20 206
use FILL  FILL53040x24100
timestamp 1618002947
transform -1 0 5512 0 -1 2610
box -4 -6 20 206
use DFFSR  _1728_
timestamp 1618002947
transform -1 0 360 0 1 2610
box -4 -6 356 206
use OAI22X1  _1559_
timestamp 1618002947
transform 1 0 360 0 1 2610
box -4 -6 84 206
use NAND2X1  _1541_
timestamp 1618002947
transform -1 0 488 0 1 2610
box -4 -6 52 206
use NOR2X1  _1455_
timestamp 1618002947
transform -1 0 536 0 1 2610
box -4 -6 52 206
use AND2X2  _1456_
timestamp 1618002947
transform 1 0 536 0 1 2610
box -4 -6 68 206
use NAND2X1  _1558_
timestamp 1618002947
transform -1 0 648 0 1 2610
box -4 -6 52 206
use NAND2X1  _1556_
timestamp 1618002947
transform -1 0 696 0 1 2610
box -4 -6 52 206
use OAI21X1  _1458_
timestamp 1618002947
transform -1 0 760 0 1 2610
box -4 -6 68 206
use NOR2X1  _1457_
timestamp 1618002947
transform 1 0 760 0 1 2610
box -4 -6 52 206
use AND2X2  _1453_
timestamp 1618002947
transform 1 0 808 0 1 2610
box -4 -6 68 206
use INVX1  _1299_
timestamp 1618002947
transform 1 0 872 0 1 2610
box -4 -6 36 206
use DFFSR  _1746_
timestamp 1618002947
transform 1 0 904 0 1 2610
box -4 -6 356 206
use AOI22X1  _1658_
timestamp 1618002947
transform -1 0 1400 0 1 2610
box -4 -6 84 206
use NAND2X1  _1653_
timestamp 1618002947
transform -1 0 1448 0 1 2610
box -4 -6 52 206
use OAI21X1  _1651_
timestamp 1618002947
transform -1 0 1512 0 1 2610
box -4 -6 68 206
use FILL  SFILL12560x26100
timestamp 1618002947
transform 1 0 1256 0 1 2610
box -4 -6 20 206
use FILL  SFILL12720x26100
timestamp 1618002947
transform 1 0 1272 0 1 2610
box -4 -6 20 206
use FILL  SFILL12880x26100
timestamp 1618002947
transform 1 0 1288 0 1 2610
box -4 -6 20 206
use FILL  SFILL13040x26100
timestamp 1618002947
transform 1 0 1304 0 1 2610
box -4 -6 20 206
use AOI21X1  _1649_
timestamp 1618002947
transform -1 0 1576 0 1 2610
box -4 -6 68 206
use NOR2X1  _1258_
timestamp 1618002947
transform 1 0 1576 0 1 2610
box -4 -6 52 206
use NAND2X1  _1259_
timestamp 1618002947
transform 1 0 1624 0 1 2610
box -4 -6 52 206
use NAND2X1  _1623_
timestamp 1618002947
transform 1 0 1672 0 1 2610
box -4 -6 52 206
use NAND3X1  _1624_
timestamp 1618002947
transform 1 0 1720 0 1 2610
box -4 -6 68 206
use NAND2X1  _1622_
timestamp 1618002947
transform -1 0 1832 0 1 2610
box -4 -6 52 206
use OAI21X1  _1621_
timestamp 1618002947
transform -1 0 1896 0 1 2610
box -4 -6 68 206
use OAI21X1  _1625_
timestamp 1618002947
transform -1 0 1960 0 1 2610
box -4 -6 68 206
use NAND3X1  _1251_
timestamp 1618002947
transform 1 0 1960 0 1 2610
box -4 -6 68 206
use INVX1  _1249_
timestamp 1618002947
transform -1 0 2056 0 1 2610
box -4 -6 36 206
use NOR2X1  _1620_
timestamp 1618002947
transform 1 0 2056 0 1 2610
box -4 -6 52 206
use NOR2X1  _1250_
timestamp 1618002947
transform -1 0 2152 0 1 2610
box -4 -6 52 206
use OAI21X1  _1613_
timestamp 1618002947
transform 1 0 2152 0 1 2610
box -4 -6 68 206
use NAND2X1  _1615_
timestamp 1618002947
transform 1 0 2216 0 1 2610
box -4 -6 52 206
use INVX1  _1612_
timestamp 1618002947
transform 1 0 2264 0 1 2610
box -4 -6 36 206
use OAI21X1  _1617_
timestamp 1618002947
transform 1 0 2296 0 1 2610
box -4 -6 68 206
use AOI22X1  _1616_
timestamp 1618002947
transform -1 0 2440 0 1 2610
box -4 -6 84 206
use INVX1  _1661_
timestamp 1618002947
transform 1 0 2440 0 1 2610
box -4 -6 36 206
use OAI21X1  _1662_
timestamp 1618002947
transform 1 0 2472 0 1 2610
box -4 -6 68 206
use OAI22X1  _1589_
timestamp 1618002947
transform -1 0 2616 0 1 2610
box -4 -6 84 206
use DFFSR  _1060_
timestamp 1618002947
transform -1 0 3032 0 1 2610
box -4 -6 356 206
use FILL  SFILL26160x26100
timestamp 1618002947
transform 1 0 2616 0 1 2610
box -4 -6 20 206
use FILL  SFILL26320x26100
timestamp 1618002947
transform 1 0 2632 0 1 2610
box -4 -6 20 206
use FILL  SFILL26480x26100
timestamp 1618002947
transform 1 0 2648 0 1 2610
box -4 -6 20 206
use FILL  SFILL26640x26100
timestamp 1618002947
transform 1 0 2664 0 1 2610
box -4 -6 20 206
use DFFSR  _1052_
timestamp 1618002947
transform 1 0 3032 0 1 2610
box -4 -6 356 206
use INVX1  _979_
timestamp 1618002947
transform 1 0 3384 0 1 2610
box -4 -6 36 206
use AND2X2  _801_
timestamp 1618002947
transform 1 0 3416 0 1 2610
box -4 -6 68 206
use DFFSR  _1048_
timestamp 1618002947
transform 1 0 3480 0 1 2610
box -4 -6 356 206
use DFFSR  _1045_
timestamp 1618002947
transform 1 0 3832 0 1 2610
box -4 -6 356 206
use NOR2X1  _793_
timestamp 1618002947
transform -1 0 4232 0 1 2610
box -4 -6 52 206
use INVX1  _802_
timestamp 1618002947
transform 1 0 4296 0 1 2610
box -4 -6 36 206
use OAI21X1  _958_
timestamp 1618002947
transform 1 0 4328 0 1 2610
box -4 -6 68 206
use FILL  SFILL42320x26100
timestamp 1618002947
transform 1 0 4232 0 1 2610
box -4 -6 20 206
use FILL  SFILL42480x26100
timestamp 1618002947
transform 1 0 4248 0 1 2610
box -4 -6 20 206
use FILL  SFILL42640x26100
timestamp 1618002947
transform 1 0 4264 0 1 2610
box -4 -6 20 206
use FILL  SFILL42800x26100
timestamp 1618002947
transform 1 0 4280 0 1 2610
box -4 -6 20 206
use OAI21X1  _952_
timestamp 1618002947
transform 1 0 4392 0 1 2610
box -4 -6 68 206
use INVX1  _890_
timestamp 1618002947
transform 1 0 4456 0 1 2610
box -4 -6 36 206
use INVX1  _798_
timestamp 1618002947
transform -1 0 4520 0 1 2610
box -4 -6 36 206
use DFFSR  _1043_
timestamp 1618002947
transform -1 0 4872 0 1 2610
box -4 -6 356 206
use DFFSR  _1239_
timestamp 1618002947
transform -1 0 5224 0 1 2610
box -4 -6 356 206
use INVX1  _933_
timestamp 1618002947
transform -1 0 5256 0 1 2610
box -4 -6 36 206
use DFFPOSX1  _1015_
timestamp 1618002947
transform 1 0 5256 0 1 2610
box -4 -6 196 206
use BUFX2  _1761_
timestamp 1618002947
transform 1 0 5448 0 1 2610
box -4 -6 52 206
use FILL  FILL53040x26100
timestamp 1618002947
transform 1 0 5496 0 1 2610
box -4 -6 20 206
use NAND3X1  _1281_
timestamp 1618002947
transform -1 0 72 0 -1 3010
box -4 -6 68 206
use INVX1  _1280_
timestamp 1618002947
transform -1 0 104 0 -1 3010
box -4 -6 36 206
use NOR2X1  _1283_
timestamp 1618002947
transform 1 0 104 0 -1 3010
box -4 -6 52 206
use INVX1  _1463_
timestamp 1618002947
transform 1 0 152 0 -1 3010
box -4 -6 36 206
use INVX1  _1459_
timestamp 1618002947
transform 1 0 184 0 -1 3010
box -4 -6 36 206
use NAND3X1  _1464_
timestamp 1618002947
transform 1 0 216 0 -1 3010
box -4 -6 68 206
use NAND2X1  _1565_
timestamp 1618002947
transform -1 0 328 0 -1 3010
box -4 -6 52 206
use NOR2X1  _1540_
timestamp 1618002947
transform 1 0 328 0 -1 3010
box -4 -6 52 206
use DFFSR  _1716_
timestamp 1618002947
transform -1 0 728 0 -1 3010
box -4 -6 356 206
use DFFSR  _1725_
timestamp 1618002947
transform -1 0 1080 0 -1 3010
box -4 -6 356 206
use NAND2X1  _1659_
timestamp 1618002947
transform -1 0 1128 0 -1 3010
box -4 -6 52 206
use OAI21X1  _1657_
timestamp 1618002947
transform -1 0 1192 0 -1 3010
box -4 -6 68 206
use NOR2X1  _1256_
timestamp 1618002947
transform 1 0 1192 0 -1 3010
box -4 -6 52 206
use OAI21X1  _1665_
timestamp 1618002947
transform 1 0 1304 0 -1 3010
box -4 -6 68 206
use INVX1  _1664_
timestamp 1618002947
transform 1 0 1368 0 -1 3010
box -4 -6 36 206
use OAI21X1  _1666_
timestamp 1618002947
transform 1 0 1400 0 -1 3010
box -4 -6 68 206
use FILL  SFILL12400x28100
timestamp 1618002947
transform -1 0 1256 0 -1 3010
box -4 -6 20 206
use FILL  SFILL12560x28100
timestamp 1618002947
transform -1 0 1272 0 -1 3010
box -4 -6 20 206
use FILL  SFILL12720x28100
timestamp 1618002947
transform -1 0 1288 0 -1 3010
box -4 -6 20 206
use FILL  SFILL12880x28100
timestamp 1618002947
transform -1 0 1304 0 -1 3010
box -4 -6 20 206
use NAND3X1  _1257_
timestamp 1618002947
transform -1 0 1528 0 -1 3010
box -4 -6 68 206
use NOR2X1  _1255_
timestamp 1618002947
transform -1 0 1576 0 -1 3010
box -4 -6 52 206
use OAI21X1  _1669_
timestamp 1618002947
transform 1 0 1576 0 -1 3010
box -4 -6 68 206
use NAND2X1  _1668_
timestamp 1618002947
transform 1 0 1640 0 -1 3010
box -4 -6 52 206
use NOR2X1  _1253_
timestamp 1618002947
transform 1 0 1688 0 -1 3010
box -4 -6 52 206
use AOI22X1  _1634_
timestamp 1618002947
transform 1 0 1736 0 -1 3010
box -4 -6 84 206
use NAND2X1  _1633_
timestamp 1618002947
transform -1 0 1864 0 -1 3010
box -4 -6 52 206
use OAI21X1  _1632_
timestamp 1618002947
transform -1 0 1928 0 -1 3010
box -4 -6 68 206
use OR2X2  _1252_
timestamp 1618002947
transform -1 0 1992 0 -1 3010
box -4 -6 68 206
use AOI22X1  _1605_
timestamp 1618002947
transform -1 0 2072 0 -1 3010
box -4 -6 84 206
use OR2X2  _1608_
timestamp 1618002947
transform -1 0 2136 0 -1 3010
box -4 -6 68 206
use NAND2X1  _1609_
timestamp 1618002947
transform -1 0 2184 0 -1 3010
box -4 -6 52 206
use AOI22X1  _1610_
timestamp 1618002947
transform -1 0 2264 0 -1 3010
box -4 -6 84 206
use AOI22X1  _1601_
timestamp 1618002947
transform -1 0 2344 0 -1 3010
box -4 -6 84 206
use AOI22X1  _1596_
timestamp 1618002947
transform -1 0 2424 0 -1 3010
box -4 -6 84 206
use AND2X2  _1675_
timestamp 1618002947
transform 1 0 2424 0 -1 3010
box -4 -6 68 206
use INVX1  _1584_
timestamp 1618002947
transform 1 0 2488 0 -1 3010
box -4 -6 36 206
use AOI21X1  _1590_
timestamp 1618002947
transform 1 0 2520 0 -1 3010
box -4 -6 68 206
use INVX1  _1673_
timestamp 1618002947
transform 1 0 2584 0 -1 3010
box -4 -6 36 206
use OAI21X1  _1676_
timestamp 1618002947
transform 1 0 2616 0 -1 3010
box -4 -6 68 206
use DFFSR  _1225_
timestamp 1618002947
transform -1 0 3096 0 -1 3010
box -4 -6 356 206
use FILL  SFILL26800x28100
timestamp 1618002947
transform -1 0 2696 0 -1 3010
box -4 -6 20 206
use FILL  SFILL26960x28100
timestamp 1618002947
transform -1 0 2712 0 -1 3010
box -4 -6 20 206
use FILL  SFILL27120x28100
timestamp 1618002947
transform -1 0 2728 0 -1 3010
box -4 -6 20 206
use FILL  SFILL27280x28100
timestamp 1618002947
transform -1 0 2744 0 -1 3010
box -4 -6 20 206
use CLKBUF1  CLKBUF1_insert12
timestamp 1618002947
transform -1 0 3240 0 -1 3010
box -4 -6 148 206
use NAND3X1  _1127_
timestamp 1618002947
transform -1 0 3304 0 -1 3010
box -4 -6 68 206
use INVX1  _982_
timestamp 1618002947
transform 1 0 3304 0 -1 3010
box -4 -6 36 206
use OAI21X1  _984_
timestamp 1618002947
transform 1 0 3336 0 -1 3010
box -4 -6 68 206
use OAI21X1  _983_
timestamp 1618002947
transform -1 0 3464 0 -1 3010
box -4 -6 68 206
use NOR2X1  _1067_
timestamp 1618002947
transform -1 0 3512 0 -1 3010
box -4 -6 52 206
use NOR3X1  _1078_
timestamp 1618002947
transform 1 0 3512 0 -1 3010
box -4 -6 132 206
use AOI21X1  _1126_
timestamp 1618002947
transform -1 0 3704 0 -1 3010
box -4 -6 68 206
use INVX2  _1091_
timestamp 1618002947
transform -1 0 3736 0 -1 3010
box -4 -6 36 206
use INVX1  _1109_
timestamp 1618002947
transform -1 0 3768 0 -1 3010
box -4 -6 36 206
use OAI21X1  _1120_
timestamp 1618002947
transform -1 0 3832 0 -1 3010
box -4 -6 68 206
use NOR2X1  _1108_
timestamp 1618002947
transform 1 0 3832 0 -1 3010
box -4 -6 52 206
use NAND2X1  _1107_
timestamp 1618002947
transform -1 0 3928 0 -1 3010
box -4 -6 52 206
use OAI21X1  _1125_
timestamp 1618002947
transform 1 0 3928 0 -1 3010
box -4 -6 68 206
use NAND2X1  _1071_
timestamp 1618002947
transform 1 0 4040 0 -1 3010
box -4 -6 52 206
use NAND2X1  _1121_
timestamp 1618002947
transform -1 0 4040 0 -1 3010
box -4 -6 52 206
use AOI21X1  _1083_
timestamp 1618002947
transform -1 0 4152 0 -1 3010
box -4 -6 68 206
use NOR2X1  _1082_
timestamp 1618002947
transform 1 0 4184 0 -1 3010
box -4 -6 52 206
use INVX1  _1081_
timestamp 1618002947
transform 1 0 4152 0 -1 3010
box -4 -6 36 206
use FILL  SFILL42480x28100
timestamp 1618002947
transform -1 0 4264 0 -1 3010
box -4 -6 20 206
use FILL  SFILL42320x28100
timestamp 1618002947
transform -1 0 4248 0 -1 3010
box -4 -6 20 206
use FILL  SFILL42800x28100
timestamp 1618002947
transform -1 0 4296 0 -1 3010
box -4 -6 20 206
use FILL  SFILL42640x28100
timestamp 1618002947
transform -1 0 4280 0 -1 3010
box -4 -6 20 206
use BUFX2  BUFX2_insert21
timestamp 1618002947
transform -1 0 4344 0 -1 3010
box -4 -6 52 206
use AOI22X1  _1124_
timestamp 1618002947
transform 1 0 4344 0 -1 3010
box -4 -6 84 206
use NAND2X1  _1123_
timestamp 1618002947
transform -1 0 4472 0 -1 3010
box -4 -6 52 206
use INVX1  _1122_
timestamp 1618002947
transform 1 0 4472 0 -1 3010
box -4 -6 36 206
use DFFSR  _1236_
timestamp 1618002947
transform -1 0 4856 0 -1 3010
box -4 -6 356 206
use AOI21X1  _862_
timestamp 1618002947
transform -1 0 4920 0 -1 3010
box -4 -6 68 206
use OAI22X1  _1158_
timestamp 1618002947
transform -1 0 5000 0 -1 3010
box -4 -6 84 206
use INVX2  _1133_
timestamp 1618002947
transform -1 0 5032 0 -1 3010
box -4 -6 36 206
use NOR2X1  _1131_
timestamp 1618002947
transform 1 0 5032 0 -1 3010
box -4 -6 52 206
use NAND2X1  _1132_
timestamp 1618002947
transform -1 0 5128 0 -1 3010
box -4 -6 52 206
use DFFSR  _1237_
timestamp 1618002947
transform -1 0 5480 0 -1 3010
box -4 -6 356 206
use FILL  FILL52880x28100
timestamp 1618002947
transform -1 0 5496 0 -1 3010
box -4 -6 20 206
use FILL  FILL53040x28100
timestamp 1618002947
transform -1 0 5512 0 -1 3010
box -4 -6 20 206
use NOR2X1  _1277_
timestamp 1618002947
transform -1 0 56 0 1 3010
box -4 -6 52 206
use NAND3X1  _1461_
timestamp 1618002947
transform 1 0 56 0 1 3010
box -4 -6 68 206
use INVX1  _1460_
timestamp 1618002947
transform -1 0 152 0 1 3010
box -4 -6 36 206
use NAND3X1  _1539_
timestamp 1618002947
transform -1 0 216 0 1 3010
box -4 -6 68 206
use NAND2X1  _1525_
timestamp 1618002947
transform 1 0 216 0 1 3010
box -4 -6 52 206
use OAI21X1  _1566_
timestamp 1618002947
transform -1 0 328 0 1 3010
box -4 -6 68 206
use NOR2X1  _1462_
timestamp 1618002947
transform 1 0 328 0 1 3010
box -4 -6 52 206
use NOR2X1  _1526_
timestamp 1618002947
transform 1 0 376 0 1 3010
box -4 -6 52 206
use OAI22X1  _1568_
timestamp 1618002947
transform 1 0 424 0 1 3010
box -4 -6 84 206
use NAND2X1  _1567_
timestamp 1618002947
transform 1 0 504 0 1 3010
box -4 -6 52 206
use NAND3X1  _1527_
timestamp 1618002947
transform 1 0 552 0 1 3010
box -4 -6 68 206
use NAND2X1  _1505_
timestamp 1618002947
transform 1 0 616 0 1 3010
box -4 -6 52 206
use OAI22X1  _1557_
timestamp 1618002947
transform 1 0 664 0 1 3010
box -4 -6 84 206
use INVX1  _1452_
timestamp 1618002947
transform 1 0 744 0 1 3010
box -4 -6 36 206
use CLKBUF1  CLKBUF1_insert7
timestamp 1618002947
transform 1 0 776 0 1 3010
box -4 -6 148 206
use OAI21X1  _1553_
timestamp 1618002947
transform 1 0 920 0 1 3010
box -4 -6 68 206
use NAND2X1  _1548_
timestamp 1618002947
transform -1 0 1032 0 1 3010
box -4 -6 52 206
use INVX4  _1530_
timestamp 1618002947
transform 1 0 1032 0 1 3010
box -4 -6 52 206
use INVX1  _1660_
timestamp 1618002947
transform 1 0 1080 0 1 3010
box -4 -6 36 206
use AND2X2  _1656_
timestamp 1618002947
transform 1 0 1192 0 1 3010
box -4 -6 68 206
use NOR2X1  _1655_
timestamp 1618002947
transform 1 0 1144 0 1 3010
box -4 -6 52 206
use INVX1  _1654_
timestamp 1618002947
transform 1 0 1112 0 1 3010
box -4 -6 36 206
use FILL  SFILL13040x30100
timestamp 1618002947
transform 1 0 1304 0 1 3010
box -4 -6 20 206
use FILL  SFILL12880x30100
timestamp 1618002947
transform 1 0 1288 0 1 3010
box -4 -6 20 206
use FILL  SFILL12720x30100
timestamp 1618002947
transform 1 0 1272 0 1 3010
box -4 -6 20 206
use FILL  SFILL12560x30100
timestamp 1618002947
transform 1 0 1256 0 1 3010
box -4 -6 20 206
use OAI21X1  _1667_
timestamp 1618002947
transform 1 0 1384 0 1 3010
box -4 -6 68 206
use NAND3X1  _1663_
timestamp 1618002947
transform -1 0 1384 0 1 3010
box -4 -6 68 206
use CLKBUF1  CLKBUF1_insert11
timestamp 1618002947
transform 1 0 1448 0 1 3010
box -4 -6 148 206
use AOI21X1  _1670_
timestamp 1618002947
transform 1 0 1592 0 1 3010
box -4 -6 68 206
use OAI21X1  _1672_
timestamp 1618002947
transform -1 0 1720 0 1 3010
box -4 -6 68 206
use OAI21X1  _1635_
timestamp 1618002947
transform -1 0 1784 0 1 3010
box -4 -6 68 206
use INVX1  _1629_
timestamp 1618002947
transform 1 0 1784 0 1 3010
box -4 -6 36 206
use NAND2X1  _1631_
timestamp 1618002947
transform 1 0 1816 0 1 3010
box -4 -6 52 206
use NOR2X1  _1630_
timestamp 1618002947
transform 1 0 1864 0 1 3010
box -4 -6 52 206
use OAI21X1  _1611_
timestamp 1618002947
transform -1 0 1976 0 1 3010
box -4 -6 68 206
use INVX1  _1248_
timestamp 1618002947
transform -1 0 2008 0 1 3010
box -4 -6 36 206
use NAND2X1  _1604_
timestamp 1618002947
transform 1 0 2008 0 1 3010
box -4 -6 52 206
use OAI21X1  _1603_
timestamp 1618002947
transform -1 0 2120 0 1 3010
box -4 -6 68 206
use OAI21X1  _1607_
timestamp 1618002947
transform 1 0 2120 0 1 3010
box -4 -6 68 206
use NAND2X1  _1595_
timestamp 1618002947
transform -1 0 2232 0 1 3010
box -4 -6 52 206
use NAND2X1  _1594_
timestamp 1618002947
transform -1 0 2280 0 1 3010
box -4 -6 52 206
use NAND2X1  _1600_
timestamp 1618002947
transform -1 0 2328 0 1 3010
box -4 -6 52 206
use OAI21X1  _1599_
timestamp 1618002947
transform -1 0 2392 0 1 3010
box -4 -6 68 206
use INVX1  _1591_
timestamp 1618002947
transform 1 0 2392 0 1 3010
box -4 -6 36 206
use OAI21X1  _1597_
timestamp 1618002947
transform 1 0 2424 0 1 3010
box -4 -6 68 206
use DFFSR  _1750_
timestamp 1618002947
transform -1 0 2840 0 1 3010
box -4 -6 356 206
use FILL  SFILL28400x30100
timestamp 1618002947
transform 1 0 2840 0 1 3010
box -4 -6 20 206
use FILL  SFILL28560x30100
timestamp 1618002947
transform 1 0 2856 0 1 3010
box -4 -6 20 206
use FILL  SFILL28720x30100
timestamp 1618002947
transform 1 0 2872 0 1 3010
box -4 -6 20 206
use FILL  SFILL28880x30100
timestamp 1618002947
transform 1 0 2888 0 1 3010
box -4 -6 20 206
use DFFSR  _1053_
timestamp 1618002947
transform -1 0 3256 0 1 3010
box -4 -6 356 206
use AOI21X1  _1129_
timestamp 1618002947
transform 1 0 3256 0 1 3010
box -4 -6 68 206
use OAI21X1  _1128_
timestamp 1618002947
transform -1 0 3384 0 1 3010
box -4 -6 68 206
use INVX1  _1114_
timestamp 1618002947
transform -1 0 3416 0 1 3010
box -4 -6 36 206
use BUFX2  _1763_
timestamp 1618002947
transform -1 0 3464 0 1 3010
box -4 -6 52 206
use OAI21X1  _1116_
timestamp 1618002947
transform 1 0 3464 0 1 3010
box -4 -6 68 206
use NAND2X1  _1115_
timestamp 1618002947
transform -1 0 3576 0 1 3010
box -4 -6 52 206
use NAND3X1  _1113_
timestamp 1618002947
transform 1 0 3576 0 1 3010
box -4 -6 68 206
use INVX1  _1104_
timestamp 1618002947
transform 1 0 3640 0 1 3010
box -4 -6 36 206
use AOI22X1  _1105_
timestamp 1618002947
transform -1 0 3752 0 1 3010
box -4 -6 84 206
use NAND2X1  _1103_
timestamp 1618002947
transform -1 0 3800 0 1 3010
box -4 -6 52 206
use AOI22X1  _1112_
timestamp 1618002947
transform 1 0 3800 0 1 3010
box -4 -6 84 206
use INVX1  _1064_
timestamp 1618002947
transform -1 0 3912 0 1 3010
box -4 -6 36 206
use OAI21X1  _1111_
timestamp 1618002947
transform -1 0 3976 0 1 3010
box -4 -6 68 206
use NAND3X1  _1070_
timestamp 1618002947
transform 1 0 3976 0 1 3010
box -4 -6 68 206
use NAND3X1  _1086_
timestamp 1618002947
transform -1 0 4104 0 1 3010
box -4 -6 68 206
use INVX1  _1110_
timestamp 1618002947
transform -1 0 4136 0 1 3010
box -4 -6 36 206
use NOR2X1  _1085_
timestamp 1618002947
transform -1 0 4184 0 1 3010
box -4 -6 52 206
use NOR3X1  _1066_
timestamp 1618002947
transform 1 0 4248 0 1 3010
box -4 -6 132 206
use FILL  SFILL41840x30100
timestamp 1618002947
transform 1 0 4184 0 1 3010
box -4 -6 20 206
use FILL  SFILL42000x30100
timestamp 1618002947
transform 1 0 4200 0 1 3010
box -4 -6 20 206
use FILL  SFILL42160x30100
timestamp 1618002947
transform 1 0 4216 0 1 3010
box -4 -6 20 206
use FILL  SFILL42320x30100
timestamp 1618002947
transform 1 0 4232 0 1 3010
box -4 -6 20 206
use INVX1  _1065_
timestamp 1618002947
transform -1 0 4408 0 1 3010
box -4 -6 36 206
use DFFSR  _1222_
timestamp 1618002947
transform 1 0 4408 0 1 3010
box -4 -6 356 206
use INVX1  _1118_
timestamp 1618002947
transform 1 0 4760 0 1 3010
box -4 -6 36 206
use CLKBUF1  CLKBUF1_insert10
timestamp 1618002947
transform -1 0 4936 0 1 3010
box -4 -6 148 206
use INVX1  _1168_
timestamp 1618002947
transform 1 0 4936 0 1 3010
box -4 -6 36 206
use NOR3X1  _1076_
timestamp 1618002947
transform -1 0 5096 0 1 3010
box -4 -6 132 206
use OAI21X1  _1172_
timestamp 1618002947
transform 1 0 5096 0 1 3010
box -4 -6 68 206
use INVX1  _1136_
timestamp 1618002947
transform 1 0 5160 0 1 3010
box -4 -6 36 206
use AOI21X1  _1164_
timestamp 1618002947
transform 1 0 5192 0 1 3010
box -4 -6 68 206
use INVX1  _1159_
timestamp 1618002947
transform 1 0 5256 0 1 3010
box -4 -6 36 206
use OAI21X1  _1162_
timestamp 1618002947
transform 1 0 5288 0 1 3010
box -4 -6 68 206
use OAI21X1  _1161_
timestamp 1618002947
transform 1 0 5352 0 1 3010
box -4 -6 68 206
use NAND2X1  _894_
timestamp 1618002947
transform -1 0 5464 0 1 3010
box -4 -6 52 206
use FILL  FILL52720x30100
timestamp 1618002947
transform 1 0 5464 0 1 3010
box -4 -6 20 206
use FILL  FILL52880x30100
timestamp 1618002947
transform 1 0 5480 0 1 3010
box -4 -6 20 206
use FILL  FILL53040x30100
timestamp 1618002947
transform 1 0 5496 0 1 3010
box -4 -6 20 206
use INVX1  _1524_
timestamp 1618002947
transform 1 0 8 0 -1 3410
box -4 -6 36 206
use DFFSR  _1731_
timestamp 1618002947
transform -1 0 392 0 -1 3410
box -4 -6 356 206
use NAND2X1  _1560_
timestamp 1618002947
transform 1 0 392 0 -1 3410
box -4 -6 52 206
use OAI21X1  _1563_
timestamp 1618002947
transform -1 0 504 0 -1 3410
box -4 -6 68 206
use NAND3X1  _1550_
timestamp 1618002947
transform 1 0 504 0 -1 3410
box -4 -6 68 206
use NAND3X1  _1528_
timestamp 1618002947
transform 1 0 568 0 -1 3410
box -4 -6 68 206
use OAI21X1  _1529_
timestamp 1618002947
transform -1 0 696 0 -1 3410
box -4 -6 68 206
use NAND2X1  _1506_
timestamp 1618002947
transform -1 0 744 0 -1 3410
box -4 -6 52 206
use NAND2X1  _1562_
timestamp 1618002947
transform -1 0 792 0 -1 3410
box -4 -6 52 206
use NOR2X1  _1561_
timestamp 1618002947
transform 1 0 792 0 -1 3410
box -4 -6 52 206
use NAND3X1  _1552_
timestamp 1618002947
transform -1 0 904 0 -1 3410
box -4 -6 68 206
use INVX1  _1551_
timestamp 1618002947
transform -1 0 936 0 -1 3410
box -4 -6 36 206
use DFFSR  _1748_
timestamp 1618002947
transform -1 0 1288 0 -1 3410
box -4 -6 356 206
use DFFSR  _1749_
timestamp 1618002947
transform 1 0 1352 0 -1 3410
box -4 -6 356 206
use FILL  SFILL12880x32100
timestamp 1618002947
transform -1 0 1304 0 -1 3410
box -4 -6 20 206
use FILL  SFILL13040x32100
timestamp 1618002947
transform -1 0 1320 0 -1 3410
box -4 -6 20 206
use FILL  SFILL13200x32100
timestamp 1618002947
transform -1 0 1336 0 -1 3410
box -4 -6 20 206
use FILL  SFILL13360x32100
timestamp 1618002947
transform -1 0 1352 0 -1 3410
box -4 -6 20 206
use BUFX2  BUFX2_insert24
timestamp 1618002947
transform -1 0 1752 0 -1 3410
box -4 -6 52 206
use OAI21X1  _1606_
timestamp 1618002947
transform -1 0 1816 0 -1 3410
box -4 -6 68 206
use INVX1  _1244_
timestamp 1618002947
transform 1 0 1816 0 -1 3410
box -4 -6 36 206
use NAND3X1  _1247_
timestamp 1618002947
transform 1 0 1848 0 -1 3410
box -4 -6 68 206
use INVX1  _1245_
timestamp 1618002947
transform 1 0 1912 0 -1 3410
box -4 -6 36 206
use OAI21X1  _1602_
timestamp 1618002947
transform 1 0 1944 0 -1 3410
box -4 -6 68 206
use NAND2X1  _1598_
timestamp 1618002947
transform 1 0 2008 0 -1 3410
box -4 -6 52 206
use BUFX2  BUFX2_insert23
timestamp 1618002947
transform 1 0 2056 0 -1 3410
box -4 -6 52 206
use INVX1  _1593_
timestamp 1618002947
transform -1 0 2136 0 -1 3410
box -4 -6 36 206
use NOR2X1  _1246_
timestamp 1618002947
transform 1 0 2136 0 -1 3410
box -4 -6 52 206
use DFFSR  _1735_
timestamp 1618002947
transform -1 0 2536 0 -1 3410
box -4 -6 356 206
use CLKBUF1  CLKBUF1_insert13
timestamp 1618002947
transform 1 0 2536 0 -1 3410
box -4 -6 148 206
use DFFSR  _1228_
timestamp 1618002947
transform 1 0 2744 0 -1 3410
box -4 -6 356 206
use FILL  SFILL26800x32100
timestamp 1618002947
transform -1 0 2696 0 -1 3410
box -4 -6 20 206
use FILL  SFILL26960x32100
timestamp 1618002947
transform -1 0 2712 0 -1 3410
box -4 -6 20 206
use FILL  SFILL27120x32100
timestamp 1618002947
transform -1 0 2728 0 -1 3410
box -4 -6 20 206
use FILL  SFILL27280x32100
timestamp 1618002947
transform -1 0 2744 0 -1 3410
box -4 -6 20 206
use DFFSR  _1224_
timestamp 1618002947
transform 1 0 3096 0 -1 3410
box -4 -6 356 206
use INVX2  _1096_
timestamp 1618002947
transform 1 0 3448 0 -1 3410
box -4 -6 36 206
use NAND2X1  _1092_
timestamp 1618002947
transform 1 0 3480 0 -1 3410
box -4 -6 52 206
use AOI21X1  _1197_
timestamp 1618002947
transform 1 0 3528 0 -1 3410
box -4 -6 68 206
use OAI21X1  _1196_
timestamp 1618002947
transform -1 0 3656 0 -1 3410
box -4 -6 68 206
use OAI21X1  _1106_
timestamp 1618002947
transform -1 0 3720 0 -1 3410
box -4 -6 68 206
use INVX1  _1102_
timestamp 1618002947
transform -1 0 3752 0 -1 3410
box -4 -6 36 206
use NAND2X1  _1093_
timestamp 1618002947
transform -1 0 3800 0 -1 3410
box -4 -6 52 206
use NAND2X1  _1068_
timestamp 1618002947
transform 1 0 3800 0 -1 3410
box -4 -6 52 206
use INVX2  _1069_
timestamp 1618002947
transform 1 0 3848 0 -1 3410
box -4 -6 36 206
use OAI21X1  _1213_
timestamp 1618002947
transform -1 0 3944 0 -1 3410
box -4 -6 68 206
use NAND2X1  _1094_
timestamp 1618002947
transform -1 0 3992 0 -1 3410
box -4 -6 52 206
use NAND2X1  _1100_
timestamp 1618002947
transform -1 0 4040 0 -1 3410
box -4 -6 52 206
use OAI21X1  _1117_
timestamp 1618002947
transform -1 0 4104 0 -1 3410
box -4 -6 68 206
use NOR2X1  _1087_
timestamp 1618002947
transform -1 0 4152 0 -1 3410
box -4 -6 52 206
use INVX1  _1084_
timestamp 1618002947
transform -1 0 4184 0 -1 3410
box -4 -6 36 206
use NOR3X1  _1101_
timestamp 1618002947
transform 1 0 4248 0 -1 3410
box -4 -6 132 206
use FILL  SFILL41840x32100
timestamp 1618002947
transform -1 0 4200 0 -1 3410
box -4 -6 20 206
use FILL  SFILL42000x32100
timestamp 1618002947
transform -1 0 4216 0 -1 3410
box -4 -6 20 206
use FILL  SFILL42160x32100
timestamp 1618002947
transform -1 0 4232 0 -1 3410
box -4 -6 20 206
use FILL  SFILL42320x32100
timestamp 1618002947
transform -1 0 4248 0 -1 3410
box -4 -6 20 206
use NAND3X1  _1090_
timestamp 1618002947
transform 1 0 4376 0 -1 3410
box -4 -6 68 206
use OAI21X1  _1089_
timestamp 1618002947
transform -1 0 4504 0 -1 3410
box -4 -6 68 206
use INVX2  _1072_
timestamp 1618002947
transform -1 0 4536 0 -1 3410
box -4 -6 36 206
use NOR2X1  _1077_
timestamp 1618002947
transform -1 0 4584 0 -1 3410
box -4 -6 52 206
use DFFSR  _1227_
timestamp 1618002947
transform 1 0 4584 0 -1 3410
box -4 -6 356 206
use NAND2X1  _1170_
timestamp 1618002947
transform -1 0 4984 0 -1 3410
box -4 -6 52 206
use OAI21X1  _1169_
timestamp 1618002947
transform -1 0 5048 0 -1 3410
box -4 -6 68 206
use INVX1  _1130_
timestamp 1618002947
transform -1 0 5080 0 -1 3410
box -4 -6 36 206
use OAI21X1  _1171_
timestamp 1618002947
transform 1 0 5080 0 -1 3410
box -4 -6 68 206
use OAI21X1  _1137_
timestamp 1618002947
transform 1 0 5144 0 -1 3410
box -4 -6 68 206
use NOR2X1  _1165_
timestamp 1618002947
transform -1 0 5256 0 -1 3410
box -4 -6 52 206
use INVX1  _1163_
timestamp 1618002947
transform 1 0 5256 0 -1 3410
box -4 -6 36 206
use OAI21X1  _1167_
timestamp 1618002947
transform 1 0 5288 0 -1 3410
box -4 -6 68 206
use OAI21X1  _1166_
timestamp 1618002947
transform 1 0 5352 0 -1 3410
box -4 -6 68 206
use INVX1  _1160_
timestamp 1618002947
transform -1 0 5448 0 -1 3410
box -4 -6 36 206
use BUFX2  _1760_
timestamp 1618002947
transform -1 0 5496 0 -1 3410
box -4 -6 52 206
use FILL  FILL53040x32100
timestamp 1618002947
transform -1 0 5512 0 -1 3410
box -4 -6 20 206
use DFFSR  _1729_
timestamp 1618002947
transform -1 0 360 0 1 3410
box -4 -6 356 206
use INVX1  _1522_
timestamp 1618002947
transform -1 0 392 0 1 3410
box -4 -6 36 206
use DFFSR  _1730_
timestamp 1618002947
transform -1 0 360 0 -1 3810
box -4 -6 356 206
use DFFSR  _1727_
timestamp 1618002947
transform 1 0 360 0 -1 3810
box -4 -6 356 206
use NOR2X1  _1523_
timestamp 1618002947
transform -1 0 440 0 1 3410
box -4 -6 52 206
use NOR2X1  _1549_
timestamp 1618002947
transform -1 0 488 0 1 3410
box -4 -6 52 206
use NOR2X1  _1447_
timestamp 1618002947
transform 1 0 488 0 1 3410
box -4 -6 52 206
use NAND2X1  _1446_
timestamp 1618002947
transform 1 0 536 0 1 3410
box -4 -6 52 206
use DFFSR  _1747_
timestamp 1618002947
transform 1 0 584 0 1 3410
box -4 -6 356 206
use DFFSR  _1240_
timestamp 1618002947
transform -1 0 1064 0 -1 3810
box -4 -6 356 206
use NOR2X1  _1445_
timestamp 1618002947
transform -1 0 984 0 1 3410
box -4 -6 52 206
use DFFSR  _1743_
timestamp 1618002947
transform 1 0 984 0 1 3410
box -4 -6 356 206
use FILL  SFILL10640x36100
timestamp 1618002947
transform -1 0 1080 0 -1 3810
box -4 -6 20 206
use FILL  SFILL10800x36100
timestamp 1618002947
transform -1 0 1096 0 -1 3810
box -4 -6 20 206
use DFFSR  _1739_
timestamp 1618002947
transform 1 0 1400 0 1 3410
box -4 -6 356 206
use DFFSR  _1242_
timestamp 1618002947
transform -1 0 1480 0 -1 3810
box -4 -6 356 206
use FILL  SFILL13360x34100
timestamp 1618002947
transform 1 0 1336 0 1 3410
box -4 -6 20 206
use FILL  SFILL13520x34100
timestamp 1618002947
transform 1 0 1352 0 1 3410
box -4 -6 20 206
use FILL  SFILL13680x34100
timestamp 1618002947
transform 1 0 1368 0 1 3410
box -4 -6 20 206
use FILL  SFILL13840x34100
timestamp 1618002947
transform 1 0 1384 0 1 3410
box -4 -6 20 206
use FILL  SFILL10960x36100
timestamp 1618002947
transform -1 0 1112 0 -1 3810
box -4 -6 20 206
use FILL  SFILL11120x36100
timestamp 1618002947
transform -1 0 1128 0 -1 3810
box -4 -6 20 206
use DFFSR  _1737_
timestamp 1618002947
transform -1 0 2104 0 1 3410
box -4 -6 356 206
use DFFSR  _1738_
timestamp 1618002947
transform 1 0 1480 0 -1 3810
box -4 -6 356 206
use DFFSR  _1736_
timestamp 1618002947
transform -1 0 2456 0 1 3410
box -4 -6 356 206
use DFFSR  _1241_
timestamp 1618002947
transform 1 0 1832 0 -1 3810
box -4 -6 356 206
use NAND3X1  _1198_
timestamp 1618002947
transform -1 0 2520 0 1 3410
box -4 -6 68 206
use NAND3X1  _1193_
timestamp 1618002947
transform -1 0 2584 0 1 3410
box -4 -6 68 206
use NAND2X1  _1199_
timestamp 1618002947
transform -1 0 2232 0 -1 3810
box -4 -6 52 206
use OAI21X1  _1195_
timestamp 1618002947
transform -1 0 2296 0 -1 3810
box -4 -6 68 206
use OAI21X1  _1184_
timestamp 1618002947
transform -1 0 2360 0 -1 3810
box -4 -6 68 206
use NAND2X1  _1194_
timestamp 1618002947
transform -1 0 2408 0 -1 3810
box -4 -6 52 206
use OAI21X1  _1207_
timestamp 1618002947
transform -1 0 2472 0 -1 3810
box -4 -6 68 206
use NAND2X1  _1208_
timestamp 1618002947
transform 1 0 2472 0 -1 3810
box -4 -6 52 206
use DFFSR  _1243_
timestamp 1618002947
transform -1 0 2872 0 -1 3810
box -4 -6 356 206
use DFFSR  _1219_
timestamp 1618002947
transform 1 0 2648 0 1 3410
box -4 -6 356 206
use FILL  SFILL25840x34100
timestamp 1618002947
transform 1 0 2584 0 1 3410
box -4 -6 20 206
use FILL  SFILL26000x34100
timestamp 1618002947
transform 1 0 2600 0 1 3410
box -4 -6 20 206
use FILL  SFILL26160x34100
timestamp 1618002947
transform 1 0 2616 0 1 3410
box -4 -6 20 206
use FILL  SFILL26320x34100
timestamp 1618002947
transform 1 0 2632 0 1 3410
box -4 -6 20 206
use FILL  SFILL28720x36100
timestamp 1618002947
transform -1 0 2888 0 -1 3810
box -4 -6 20 206
use FILL  SFILL28880x36100
timestamp 1618002947
transform -1 0 2904 0 -1 3810
box -4 -6 20 206
use FILL  SFILL29200x36100
timestamp 1618002947
transform -1 0 2936 0 -1 3810
box -4 -6 20 206
use FILL  SFILL29040x36100
timestamp 1618002947
transform -1 0 2920 0 -1 3810
box -4 -6 20 206
use OAI21X1  _1216_
timestamp 1618002947
transform -1 0 3000 0 -1 3810
box -4 -6 68 206
use NAND2X1  _1217_
timestamp 1618002947
transform 1 0 3000 0 -1 3810
box -4 -6 52 206
use NAND3X1  _1215_
timestamp 1618002947
transform -1 0 3064 0 1 3410
box -4 -6 68 206
use NAND3X1  _1206_
timestamp 1618002947
transform 1 0 3080 0 -1 3810
box -4 -6 68 206
use INVX2  _1190_
timestamp 1618002947
transform -1 0 3080 0 -1 3810
box -4 -6 36 206
use NOR2X1  _1178_
timestamp 1618002947
transform -1 0 3112 0 1 3410
box -4 -6 52 206
use NOR2X1  _1189_
timestamp 1618002947
transform 1 0 3144 0 -1 3810
box -4 -6 52 206
use NAND2X1  _1187_
timestamp 1618002947
transform 1 0 3176 0 1 3410
box -4 -6 52 206
use AND2X2  _1179_
timestamp 1618002947
transform -1 0 3176 0 1 3410
box -4 -6 68 206
use OAI21X1  _1188_
timestamp 1618002947
transform 1 0 3192 0 -1 3810
box -4 -6 68 206
use NAND3X1  _1173_
timestamp 1618002947
transform -1 0 3288 0 1 3410
box -4 -6 68 206
use AND2X2  _1176_
timestamp 1618002947
transform -1 0 3480 0 -1 3810
box -4 -6 68 206
use NAND2X1  _1186_
timestamp 1618002947
transform -1 0 3416 0 -1 3810
box -4 -6 52 206
use NAND2X1  _1180_
timestamp 1618002947
transform -1 0 3368 0 -1 3810
box -4 -6 52 206
use NAND3X1  _1181_
timestamp 1618002947
transform 1 0 3256 0 -1 3810
box -4 -6 68 206
use NOR2X1  _1192_
timestamp 1618002947
transform -1 0 3464 0 1 3410
box -4 -6 52 206
use NAND3X1  _1191_
timestamp 1618002947
transform -1 0 3416 0 1 3410
box -4 -6 68 206
use AOI21X1  _1185_
timestamp 1618002947
transform -1 0 3352 0 1 3410
box -4 -6 68 206
use OAI21X1  _1183_
timestamp 1618002947
transform -1 0 3640 0 1 3410
box -4 -6 68 206
use OAI21X1  _1182_
timestamp 1618002947
transform 1 0 3512 0 1 3410
box -4 -6 68 206
use NOR2X1  _1177_
timestamp 1618002947
transform -1 0 3512 0 1 3410
box -4 -6 52 206
use DFFSR  _1218_
timestamp 1618002947
transform 1 0 3480 0 -1 3810
box -4 -6 356 206
use OAI22X1  _1095_
timestamp 1618002947
transform 1 0 3640 0 1 3410
box -4 -6 84 206
use OAI21X1  _1204_
timestamp 1618002947
transform -1 0 3784 0 1 3410
box -4 -6 68 206
use AOI21X1  _1205_
timestamp 1618002947
transform -1 0 3848 0 1 3410
box -4 -6 68 206
use INVX2  _1073_
timestamp 1618002947
transform -1 0 3880 0 1 3410
box -4 -6 36 206
use AOI21X1  _1214_
timestamp 1618002947
transform -1 0 3944 0 1 3410
box -4 -6 68 206
use AOI21X1  _1212_
timestamp 1618002947
transform 1 0 3944 0 1 3410
box -4 -6 68 206
use NOR2X1  _1175_
timestamp 1618002947
transform 1 0 3832 0 -1 3810
box -4 -6 52 206
use OAI21X1  _1174_
timestamp 1618002947
transform -1 0 3944 0 -1 3810
box -4 -6 68 206
use DFFSR  _1223_
timestamp 1618002947
transform 1 0 3944 0 -1 3810
box -4 -6 356 206
use NOR3X1  _1202_
timestamp 1618002947
transform 1 0 4072 0 1 3410
box -4 -6 132 206
use AOI21X1  _1203_
timestamp 1618002947
transform 1 0 4008 0 1 3410
box -4 -6 68 206
use NOR2X1  _1074_
timestamp 1618002947
transform -1 0 4248 0 1 3410
box -4 -6 52 206
use FILL  SFILL43280x36100
timestamp 1618002947
transform -1 0 4344 0 -1 3810
box -4 -6 20 206
use FILL  SFILL43120x36100
timestamp 1618002947
transform -1 0 4328 0 -1 3810
box -4 -6 20 206
use FILL  SFILL42960x36100
timestamp 1618002947
transform -1 0 4312 0 -1 3810
box -4 -6 20 206
use FILL  SFILL42960x34100
timestamp 1618002947
transform 1 0 4296 0 1 3410
box -4 -6 20 206
use FILL  SFILL42800x34100
timestamp 1618002947
transform 1 0 4280 0 1 3410
box -4 -6 20 206
use FILL  SFILL42640x34100
timestamp 1618002947
transform 1 0 4264 0 1 3410
box -4 -6 20 206
use FILL  SFILL42480x34100
timestamp 1618002947
transform 1 0 4248 0 1 3410
box -4 -6 20 206
use NAND2X1  _1075_
timestamp 1618002947
transform 1 0 4312 0 1 3410
box -4 -6 52 206
use NAND2X1  _1088_
timestamp 1618002947
transform 1 0 4360 0 1 3410
box -4 -6 52 206
use NAND3X1  _1080_
timestamp 1618002947
transform 1 0 4408 0 1 3410
box -4 -6 68 206
use OAI21X1  _1079_
timestamp 1618002947
transform 1 0 4472 0 1 3410
box -4 -6 68 206
use OAI22X1  _1099_
timestamp 1618002947
transform 1 0 4536 0 1 3410
box -4 -6 84 206
use OAI21X1  _1098_
timestamp 1618002947
transform -1 0 4680 0 1 3410
box -4 -6 68 206
use INVX1  _866_
timestamp 1618002947
transform -1 0 4712 0 1 3410
box -4 -6 36 206
use DFFSR  _1220_
timestamp 1618002947
transform -1 0 4712 0 -1 3810
box -4 -6 356 206
use FILL  SFILL43440x36100
timestamp 1618002947
transform -1 0 4360 0 -1 3810
box -4 -6 20 206
use OAI21X1  _1201_
timestamp 1618002947
transform 1 0 4712 0 1 3410
box -4 -6 68 206
use OAI21X1  _1211_
timestamp 1618002947
transform 1 0 4776 0 1 3410
box -4 -6 68 206
use INVX1  _1097_
timestamp 1618002947
transform 1 0 4840 0 1 3410
box -4 -6 36 206
use INVX1  _1209_
timestamp 1618002947
transform 1 0 4872 0 1 3410
box -4 -6 36 206
use NAND3X1  _1210_
timestamp 1618002947
transform 1 0 4904 0 1 3410
box -4 -6 68 206
use NAND3X1  _1200_
timestamp 1618002947
transform 1 0 4968 0 1 3410
box -4 -6 68 206
use NOR2X1  _868_
timestamp 1618002947
transform -1 0 5080 0 1 3410
box -4 -6 52 206
use DFFSR  _1221_
timestamp 1618002947
transform 1 0 4712 0 -1 3810
box -4 -6 356 206
use AOI21X1  _1119_
timestamp 1618002947
transform -1 0 5144 0 1 3410
box -4 -6 68 206
use DFFSR  _1238_
timestamp 1618002947
transform -1 0 5496 0 1 3410
box -4 -6 356 206
use NAND2X1  _869_
timestamp 1618002947
transform 1 0 5064 0 -1 3810
box -4 -6 52 206
use DFFSR  _1226_
timestamp 1618002947
transform -1 0 5464 0 -1 3810
box -4 -6 356 206
use INVX1  _887_
timestamp 1618002947
transform -1 0 5496 0 -1 3810
box -4 -6 36 206
use FILL  FILL53040x34100
timestamp 1618002947
transform 1 0 5496 0 1 3410
box -4 -6 20 206
use FILL  FILL53040x36100
timestamp 1618002947
transform -1 0 5512 0 -1 3810
box -4 -6 20 206
<< labels >>
flabel metal4 s 2720 -10 2784 0 7 FreeSans 24 270 0 0 gnd
port 0 nsew
flabel metal4 s 1216 -10 1280 0 7 FreeSans 24 270 0 0 vdd
port 1 nsew
flabel metal2 s 2061 3857 2067 3863 3 FreeSans 24 90 0 0 arst_i
port 2 nsew
flabel metal2 s 3293 -23 3299 -17 7 FreeSans 24 270 0 0 scl_pad_i
port 3 nsew
flabel metal2 s 1741 -23 1747 -17 7 FreeSans 24 270 0 0 scl_pad_o
port 4 nsew
flabel metal3 s -35 1497 -29 1503 7 FreeSans 24 0 0 0 scl_padoen_o
port 5 nsew
flabel metal2 s 765 -23 771 -17 7 FreeSans 24 270 0 0 sda_pad_i
port 6 nsew
flabel metal2 s 1789 -23 1795 -17 7 FreeSans 24 270 0 0 sda_pad_o
port 7 nsew
flabel metal2 s 733 -23 739 -17 7 FreeSans 24 270 0 0 sda_padoen_o
port 8 nsew
flabel metal3 s 5549 2397 5555 2403 3 FreeSans 24 0 0 0 wb_ack_o
port 9 nsew
flabel metal3 s 5549 1757 5555 1763 3 FreeSans 24 0 0 0 wb_adr_i[2]
port 10 nsew
flabel metal3 s 5549 1797 5555 1803 3 FreeSans 24 0 0 0 wb_adr_i[1]
port 11 nsew
flabel metal3 s 5549 1697 5555 1703 3 FreeSans 24 0 0 0 wb_adr_i[0]
port 12 nsew
flabel metal2 s 5165 -23 5171 -17 7 FreeSans 24 270 0 0 wb_clk_i
port 13 nsew
flabel metal3 s 5549 3117 5555 3123 3 FreeSans 24 0 0 0 wb_cyc_i
port 14 nsew
flabel metal3 s 5549 2357 5555 2363 3 FreeSans 24 0 0 0 wb_dat_i[7]
port 15 nsew
flabel metal2 s 3437 3857 3443 3863 3 FreeSans 24 90 0 0 wb_dat_i[6]
port 16 nsew
flabel metal3 s 5549 2277 5555 2283 3 FreeSans 24 0 0 0 wb_dat_i[5]
port 17 nsew
flabel metal2 s 3261 -23 3267 -17 7 FreeSans 24 270 0 0 wb_dat_i[4]
port 18 nsew
flabel metal2 s 4701 -23 4707 -17 7 FreeSans 24 270 0 0 wb_dat_i[3]
port 19 nsew
flabel metal2 s 3165 -23 3171 -17 7 FreeSans 24 270 0 0 wb_dat_i[2]
port 20 nsew
flabel metal2 s 3517 -23 3523 -17 7 FreeSans 24 270 0 0 wb_dat_i[1]
port 21 nsew
flabel metal2 s 3213 -23 3219 -17 7 FreeSans 24 270 0 0 wb_dat_i[0]
port 22 nsew
flabel metal2 s 3405 3857 3411 3863 3 FreeSans 24 90 0 0 wb_dat_o[7]
port 23 nsew
flabel metal3 s 5549 97 5555 103 3 FreeSans 24 0 0 0 wb_dat_o[6]
port 24 nsew
flabel metal3 s 5549 2697 5555 2703 3 FreeSans 24 0 0 0 wb_dat_o[5]
port 25 nsew
flabel metal3 s 5549 3297 5555 3303 3 FreeSans 24 0 0 0 wb_dat_o[4]
port 26 nsew
flabel metal2 s 4589 -23 4595 -17 7 FreeSans 24 270 0 0 wb_dat_o[3]
port 27 nsew
flabel metal3 s 5549 1497 5555 1503 3 FreeSans 24 0 0 0 wb_dat_o[2]
port 28 nsew
flabel metal2 s 4637 -23 4643 -17 7 FreeSans 24 270 0 0 wb_dat_o[1]
port 29 nsew
flabel metal2 s 3741 -23 3747 -17 7 FreeSans 24 270 0 0 wb_dat_o[0]
port 30 nsew
flabel metal2 s 5421 -23 5427 -17 7 FreeSans 24 270 0 0 wb_inta_o
port 31 nsew
flabel metal2 s 2813 -23 2819 -17 7 FreeSans 24 270 0 0 wb_rst_i
port 32 nsew
flabel metal3 s 5549 3077 5555 3083 3 FreeSans 24 0 0 0 wb_stb_i
port 33 nsew
flabel metal3 s 5549 2317 5555 2323 3 FreeSans 24 0 0 0 wb_we_i
port 34 nsew
<< end >>
