* NGSPICE file created from map9v3.ext - technology: scmos

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR Q CLK R S D gnd vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

.subckt map9v3 gnd vdd N[8] N[7] N[6] N[5] N[4] N[3] N[2] N[1] N[0] clock counter[7]
+ counter[6] counter[5] counter[4] counter[3] counter[2] counter[1] counter[0] done
+ dp[8] dp[7] dp[6] dp[5] dp[4] dp[3] dp[2] dp[1] dp[0] reset sr[7] sr[6] sr[5] sr[4]
+ sr[3] sr[2] sr[1] sr[0] start
X_294_ _320_/A _291_/CLK _297_/R vdd _294_/D gnd vdd DFFSR
XSFILL18640x10100 gnd vdd FILL
XSFILL17840x6100 gnd vdd FILL
X_200_ N[5] _200_/B N[6] gnd _203_/C vdd OAI21X1
X_277_ _303_/A _275_/CLK _275_/R vdd _181_/Y gnd vdd DFFSR
XSFILL6320x6100 gnd vdd FILL
X_293_ _233_/A _291_/CLK _297_/R vdd _264_/Y gnd vdd DFFSR
X_276_ _302_/A _275_/CLK _275_/R vdd _172_/Y gnd vdd DFFSR
XSFILL18640x2100 gnd vdd FILL
X_259_ _257_/Y _198_/B _259_/C gnd _259_/Y vdd OAI21X1
X_292_ _258_/A _292_/CLK _275_/R vdd _259_/Y gnd vdd DFFSR
X_275_ _275_/Q _275_/CLK _275_/R vdd _163_/Y gnd vdd DFFSR
X_258_ _258_/A _160_/B gnd _259_/C vdd NAND2X1
XFILL23760x12100 gnd vdd FILL
X_189_ _200_/B gnd _190_/B vdd INVX1
XSFILL5200x100 gnd vdd FILL
XSFILL18640x8100 gnd vdd FILL
XSFILL8080x4100 gnd vdd FILL
XSFILL8400x4100 gnd vdd FILL
X_291_ _318_/A _291_/CLK _297_/R vdd _291_/D gnd vdd DFFSR
X_274_ _274_/Q _282_/CLK _269_/R vdd _154_/A gnd vdd DFFSR
X_326_ _326_/A gnd sr[7] vdd BUFX2
X_309_ _258_/A gnd done vdd BUFX2
X_188_ _188_/A _167_/Y _187_/Y gnd _200_/B vdd OAI21X1
XSFILL18320x12100 gnd vdd FILL
X_257_ _257_/A _257_/B gnd _257_/Y vdd NAND2X1
XSFILL5840x6100 gnd vdd FILL
X_290_ _252_/A _275_/CLK _275_/R vdd _253_/Y gnd vdd DFFSR
X_187_ N[3] N[4] gnd _187_/Y vdd NOR2X1
X_325_ _325_/A gnd sr[6] vdd BUFX2
X_256_ _256_/A _244_/B _255_/Y gnd _291_/D vdd AOI21X1
X_273_ _154_/A _296_/CLK _273_/R vdd start gnd vdd DFFSR
X_239_ _295_/Q gnd _136_/C vdd INVX1
X_308_ _218_/A gnd counter[7] vdd BUFX2
XSFILL18800x14100 gnd vdd FILL
X_272_ _257_/A _282_/CLK _269_/R vdd _229_/A gnd vdd DFFSR
X_255_ _318_/A _244_/B gnd _255_/Y vdd NOR2X1
X_186_ N[3] _175_/Y N[4] gnd _191_/C vdd OAI21X1
X_324_ _260_/B gnd sr[5] vdd BUFX2
XBUFX2_insert5 _141_/Y gnd _269_/R vdd BUFX2
XSFILL7920x4100 gnd vdd FILL
X_169_ N[1] N[2] gnd _169_/Y vdd NAND2X1
XFILL23920x10100 gnd vdd FILL
XSFILL6640x8100 gnd vdd FILL
X_238_ _236_/Y _238_/B _238_/C gnd _285_/D vdd AOI21X1
XSFILL6160x2100 gnd vdd FILL
X_307_ _147_/A gnd counter[6] vdd BUFX2
XSFILL6800x12100 gnd vdd FILL
X_254_ _326_/A gnd _256_/A vdd INVX1
X_185_ _185_/A gnd _191_/B vdd INVX1
X_323_ _245_/A gnd sr[4] vdd BUFX2
XSFILL18960x4100 gnd vdd FILL
X_271_ _164_/A _292_/CLK _299_/R vdd _271_/D gnd vdd DFFSR
X_306_ _213_/A gnd counter[5] vdd BUFX2
X_168_ _188_/A _167_/Y gnd _170_/A vdd NAND2X1
XSFILL5360x100 gnd vdd FILL
X_237_ _312_/A _238_/B gnd _238_/C vdd NOR2X1
XBUFX2_insert6 _141_/Y gnd _297_/R vdd BUFX2
XSFILL6000x2100 gnd vdd FILL
X_270_ _229_/A _292_/CLK _299_/R vdd _270_/D gnd vdd DFFSR
X_253_ _251_/Y _253_/B _252_/Y gnd _253_/Y vdd AOI21X1
X_184_ _304_/A _183_/Y gnd _192_/C vdd NAND2X1
XBUFX2_insert7 _141_/Y gnd _275_/R vdd BUFX2
X_322_ _261_/B gnd sr[3] vdd BUFX2
X_305_ _305_/A gnd counter[4] vdd BUFX2
X_167_ N[2] gnd _167_/Y vdd INVX1
X_236_ _320_/A gnd _236_/Y vdd INVX1
X_219_ N[7] _209_/Y N[8] gnd _219_/Y vdd OAI21X1
XSFILL18800x4100 gnd vdd FILL
XSFILL18480x10100 gnd vdd FILL
X_252_ _252_/A _253_/B gnd _252_/Y vdd NOR2X1
X_235_ _235_/A _253_/B _235_/C gnd _284_/D vdd AOI21X1
X_166_ N[1] gnd _188_/A vdd INVX1
X_183_ _173_/A _179_/Y _198_/B gnd _183_/Y vdd OAI21X1
XSFILL5680x2100 gnd vdd FILL
X_304_ _304_/A gnd counter[3] vdd BUFX2
X_321_ _295_/Q gnd sr[2] vdd BUFX2
XBUFX2_insert8 _141_/Y gnd _273_/R vdd BUFX2
X_149_ _147_/Y _148_/Y gnd _150_/B vdd NAND2X1
X_218_ _218_/A gnd _227_/A vdd INVX1
XCLKBUF1_insert0 clock gnd _282_/CLK vdd CLKBUF1
X_251_ _325_/A gnd _251_/Y vdd INVX1
X_182_ _162_/B gnd _198_/B vdd INVX4
X_320_ _320_/A gnd sr[1] vdd BUFX2
XBUFX2_insert9 _141_/Y gnd _299_/R vdd BUFX2
X_303_ _303_/A gnd counter[2] vdd BUFX2
X_165_ _302_/A _164_/Y gnd _172_/C vdd NAND2X1
X_234_ _311_/A _253_/B gnd _235_/C vdd NOR2X1
X_148_ _213_/A _305_/A gnd _148_/Y vdd NOR2X1
XCLKBUF1_insert1 clock gnd _292_/CLK vdd CLKBUF1
X_217_ _217_/A _212_/Y _217_/C gnd _281_/D vdd NAND3X1
XSFILL8400x14100 gnd vdd FILL
XSFILL19120x100 gnd vdd FILL
X_302_ _302_/A gnd counter[1] vdd BUFX2
X_233_ _233_/A gnd _235_/A vdd INVX1
X_164_ _164_/A _173_/A _160_/Y gnd _164_/Y vdd OAI21X1
X_181_ _162_/B _180_/Y _181_/C gnd _181_/Y vdd OAI21X1
X_250_ _248_/Y _231_/B _249_/Y gnd _289_/D vdd AOI21X1
XFILL23920x2100 gnd vdd FILL
X_147_ _147_/A _218_/A gnd _147_/Y vdd NOR2X1
X_216_ _225_/B _215_/Y _265_/A gnd _217_/C vdd OAI21X1
XCLKBUF1_insert2 clock gnd _275_/CLK vdd CLKBUF1
XSFILL6960x10100 gnd vdd FILL
X_180_ _160_/B _179_/Y _180_/C gnd _180_/Y vdd AOI21X1
X_301_ _275_/Q gnd counter[0] vdd BUFX2
X_163_ _162_/B _161_/Y _163_/C gnd _163_/Y vdd OAI21X1
XFILL23920x8100 gnd vdd FILL
X_232_ _228_/Y _231_/B _232_/C gnd _232_/Y vdd OAI21X1
X_146_ _144_/Y _145_/Y gnd _185_/A vdd NAND2X1
X_215_ _215_/A gnd _215_/Y vdd INVX1
XCLKBUF1_insert3 clock gnd _296_/CLK vdd CLKBUF1
XSFILL5520x100 gnd vdd FILL
X_162_ _275_/Q _162_/B gnd _163_/C vdd NAND2X1
X_300_ _326_/A _291_/CLK _297_/R vdd _140_/Y gnd vdd DFFSR
X_231_ N[0] _231_/B gnd _232_/C vdd NAND2X1
X_145_ _304_/A _303_/A gnd _145_/Y vdd NOR2X1
X_214_ _213_/A _206_/B _147_/A gnd _215_/A vdd OAI21X1
XCLKBUF1_insert4 clock gnd _291_/CLK vdd CLKBUF1
X_161_ _160_/B N[1] _160_/Y gnd _161_/Y vdd OAI21X1
X_230_ _257_/B _198_/B gnd _230_/Y vdd NOR2X1
X_144_ _302_/A _275_/Q gnd _144_/Y vdd NOR2X1
XFILL23760x10100 gnd vdd FILL
X_213_ _213_/A _147_/A _206_/B gnd _225_/B vdd NOR3X1
XSFILL6160x16100 gnd vdd FILL
XSFILL6640x12100 gnd vdd FILL
XSFILL19280x100 gnd vdd FILL
X_160_ _275_/Q _160_/B gnd _160_/Y vdd NAND2X1
XBUFX2_insert10 _230_/Y gnd _253_/B vdd BUFX2
X_143_ _173_/A gnd _160_/B vdd INVX4
X_289_ _316_/A _296_/CLK _273_/R vdd _289_/D gnd vdd DFFSR
X_212_ _147_/A _162_/B gnd _212_/Y vdd NAND2X1
XSFILL18320x10100 gnd vdd FILL
XSFILL18160x6100 gnd vdd FILL
X_288_ _246_/A _275_/CLK _297_/R vdd _247_/Y gnd vdd DFFSR
XBUFX2_insert11 _230_/Y gnd _244_/B vdd BUFX2
X_142_ _164_/A gnd _196_/B vdd INVX1
X_211_ _173_/A _211_/B gnd _217_/A vdd NAND2X1
XSFILL18800x12100 gnd vdd FILL
XSFILL5680x100 gnd vdd FILL
X_287_ _243_/A _291_/CLK _297_/R vdd _287_/D gnd vdd DFFSR
X_210_ _209_/Y N[7] gnd _211_/B vdd XOR2X1
XSFILL18000x6100 gnd vdd FILL
XBUFX2_insert12 _230_/Y gnd _238_/B vdd BUFX2
X_141_ reset gnd _141_/Y vdd INVX8
XSFILL19280x16100 gnd vdd FILL
X_286_ _240_/A _296_/CLK _273_/R vdd _286_/D gnd vdd DFFSR
XBUFX2_insert13 _230_/Y gnd _231_/B vdd BUFX2
X_140_ _256_/A _198_/B _251_/Y _140_/D gnd _140_/Y vdd OAI22X1
X_269_ _153_/A _282_/CLK _269_/R vdd _269_/D gnd vdd DFFSR
XSFILL6800x10100 gnd vdd FILL
XSFILL8240x14100 gnd vdd FILL
XFILL23920x14100 gnd vdd FILL
X_285_ _312_/A _296_/CLK _273_/R vdd _285_/D gnd vdd DFFSR
XSFILL6160x6100 gnd vdd FILL
X_199_ _199_/A _173_/A _199_/C gnd _199_/Y vdd AOI21X1
X_268_ _173_/A _282_/CLK vdd _269_/R _157_/Y gnd vdd DFFSR
XSFILL18480x2100 gnd vdd FILL
XSFILL18800x2100 gnd vdd FILL
X_284_ _311_/A _292_/CLK _299_/R vdd _284_/D gnd vdd DFFSR
XSFILL5840x16100 gnd vdd FILL
X_198_ _305_/A _198_/B _197_/Y _195_/Y gnd _199_/C vdd OAI22X1
X_267_ _136_/C _198_/B _236_/Y _140_/D gnd _295_/D vdd OAI22X1
XSFILL6000x6100 gnd vdd FILL
X_319_ _233_/A gnd sr[0] vdd BUFX2
XSFILL18320x2100 gnd vdd FILL
XSFILL19440x100 gnd vdd FILL
XSFILL18800x8100 gnd vdd FILL
XSFILL18480x8100 gnd vdd FILL
X_283_ _283_/Q _282_/CLK _269_/R vdd _232_/Y gnd vdd DFFSR
XSFILL8240x4100 gnd vdd FILL
XSFILL6000x16100 gnd vdd FILL
X_318_ _318_/A gnd dp[8] vdd BUFX2
X_266_ _236_/Y _198_/B _235_/A _140_/D gnd _294_/D vdd OAI22X1
X_197_ _305_/A _185_/A _265_/A gnd _197_/Y vdd OAI21X1
X_249_ _316_/A _231_/B gnd _249_/Y vdd NOR2X1
XSFILL18320x8100 gnd vdd FILL
X_196_ _173_/A _196_/B gnd _265_/A vdd NOR2X1
X_282_ _218_/A _282_/CLK _269_/R vdd _282_/D gnd vdd DFFSR
X_265_ _265_/A gnd _140_/D vdd INVX4
X_317_ _252_/A gnd dp[7] vdd BUFX2
X_179_ _144_/Y _179_/B gnd _179_/Y vdd AND2X2
X_248_ _260_/B gnd _248_/Y vdd INVX1
XSFILL18960x16100 gnd vdd FILL
XSFILL6480x12100 gnd vdd FILL
X_281_ _147_/A _282_/CLK _269_/R vdd _281_/D gnd vdd DFFSR
X_247_ _247_/A _244_/B _247_/C gnd _247_/Y vdd AOI21X1
X_264_ _235_/A _198_/B _262_/Y _263_/Y gnd _264_/Y vdd OAI22X1
X_195_ _195_/A _191_/B gnd _195_/Y vdd NOR2X1
X_316_ _316_/A gnd dp[6] vdd BUFX2
XSFILL19120x4100 gnd vdd FILL
X_178_ _303_/A gnd _179_/B vdd INVX1
XSFILL7920x14100 gnd vdd FILL
X_263_ _260_/Y _262_/A _265_/A gnd _263_/Y vdd OAI21X1
X_194_ _305_/A gnd _195_/A vdd INVX1
X_280_ _213_/A _292_/CLK _299_/R vdd _280_/D gnd vdd DFFSR
XSFILL6800x8100 gnd vdd FILL
XSFILL6480x8100 gnd vdd FILL
XSFILL19120x16100 gnd vdd FILL
X_315_ _246_/A gnd dp[5] vdd BUFX2
X_246_ _246_/A _253_/B gnd _247_/C vdd NOR2X1
X_177_ N[3] _175_/Y _176_/Y gnd _180_/C vdd AOI21X1
X_229_ _229_/A gnd _257_/B vdd INVX1
XSFILL18640x12100 gnd vdd FILL
X_193_ _200_/B N[5] gnd _199_/A vdd XNOR2X1
X_262_ _262_/A _260_/Y gnd _262_/Y vdd AND2X2
X_159_ _164_/A _173_/A gnd _162_/B vdd NOR2X1
X_314_ _243_/A gnd dp[4] vdd BUFX2
X_176_ N[3] _175_/Y _173_/A gnd _176_/Y vdd OAI21X1
XSFILL6320x8100 gnd vdd FILL
X_245_ _245_/A gnd _247_/A vdd INVX1
X_228_ _283_/Q gnd _228_/Y vdd INVX1
X_192_ _162_/B _192_/B _192_/C gnd _278_/D vdd OAI21X1
X_261_ _245_/A _261_/B gnd _262_/A vdd XOR2X1
XSFILL18640x4100 gnd vdd FILL
X_175_ _169_/Y gnd _175_/Y vdd INVX1
XSFILL6640x10100 gnd vdd FILL
X_244_ _244_/A _244_/B _244_/C gnd _287_/D vdd AOI21X1
X_313_ _240_/A gnd dp[3] vdd BUFX2
XSFILL8080x14100 gnd vdd FILL
X_227_ _227_/A _162_/B _227_/C _226_/Y gnd _282_/D vdd AOI22X1
X_158_ _150_/Y _164_/A gnd _270_/D vdd AND2X2
XSFILL19600x100 gnd vdd FILL
XSFILL5840x2100 gnd vdd FILL
X_191_ _160_/B _191_/B _191_/C _191_/D gnd _192_/B vdd AOI22X1
X_260_ _326_/A _260_/B gnd _260_/Y vdd XNOR2X1
X_174_ _162_/B _174_/B _303_/A gnd _181_/C vdd OAI21X1
X_243_ _243_/A _244_/B gnd _244_/C vdd NOR2X1
X_226_ _160_/B _150_/Y _225_/Y gnd _226_/Y vdd AOI21X1
X_312_ _312_/A gnd dp[2] vdd BUFX2
X_157_ _157_/A _153_/A gnd _157_/Y vdd AND2X2
X_209_ _169_/Y _187_/Y _209_/C gnd _209_/Y vdd NAND3X1
XSFILL5680x16100 gnd vdd FILL
X_311_ _311_/A gnd dp[1] vdd BUFX2
X_173_ _173_/A _144_/Y gnd _174_/B vdd NOR2X1
XSFILL18800x10100 gnd vdd FILL
X_190_ _160_/B _190_/B gnd _191_/D vdd NOR2X1
X_242_ _261_/B gnd _244_/A vdd INVX1
X_225_ _225_/A _225_/B _198_/B gnd _225_/Y vdd OAI21X1
X_156_ _156_/A _157_/A _152_/Y gnd _269_/D vdd OAI21X1
X_208_ _208_/A _173_/A _207_/Y gnd _280_/D vdd AOI21X1
X_139_ _251_/Y _198_/B _248_/Y _140_/D gnd _139_/Y vdd OAI22X1
XFILL23760x2100 gnd vdd FILL
XSFILL19280x14100 gnd vdd FILL
X_172_ _162_/B _171_/Y _172_/C gnd _172_/Y vdd OAI21X1
X_224_ _218_/A _160_/B gnd _225_/A vdd NAND2X1
X_241_ _136_/C _238_/B _240_/Y gnd _286_/D vdd AOI21X1
X_310_ _283_/Q gnd dp[0] vdd BUFX2
X_155_ _274_/Q _154_/Y gnd _157_/A vdd NOR2X1
XSFILL18800x16100 gnd vdd FILL
XSFILL6320x12100 gnd vdd FILL
X_207_ _213_/A _198_/B _205_/Y _206_/Y gnd _207_/Y vdd OAI22X1
X_138_ _248_/Y _198_/B _247_/A _140_/D gnd _138_/Y vdd OAI22X1
X_171_ _160_/B _144_/Y _171_/C gnd _171_/Y vdd AOI21X1
X_240_ _240_/A _238_/B gnd _240_/Y vdd NOR2X1
XFILL23920x12100 gnd vdd FILL
X_223_ _173_/A _219_/Y _222_/Y gnd _227_/C vdd NAND3X1
X_154_ _154_/A gnd _154_/Y vdd INVX1
X_206_ _213_/A _206_/B _265_/A gnd _206_/Y vdd OAI21X1
X_137_ _247_/A _198_/B _244_/A _140_/D gnd _297_/D vdd OAI22X1
X_170_ _170_/A _169_/Y _160_/B gnd _171_/C vdd AOI21X1
X_299_ _325_/A _292_/CLK _299_/R vdd _139_/Y gnd vdd DFFSR
X_205_ _206_/B _213_/A gnd _205_/Y vdd AND2X2
X_153_ _153_/A gnd _156_/A vdd INVX1
X_222_ _220_/Y _222_/B gnd _222_/Y vdd NAND2X1
X_136_ _244_/A _198_/B _136_/C _140_/D gnd _296_/D vdd OAI22X1
X_298_ _260_/B _292_/CLK _299_/R vdd _138_/Y gnd vdd DFFSR
X_221_ N[7] _209_/Y gnd _222_/B vdd NOR2X1
X_152_ _257_/A gnd _152_/Y vdd INVX1
X_204_ _195_/A _144_/Y _145_/Y gnd _206_/B vdd NAND3X1
XSFILL18480x12100 gnd vdd FILL
X_297_ _245_/A _291_/CLK _297_/R vdd _297_/D gnd vdd DFFSR
X_203_ _200_/B _203_/B _203_/C gnd _208_/A vdd OAI21X1
X_151_ _196_/B _150_/Y _160_/B gnd _271_/D vdd OAI21X1
XSFILL18320x6100 gnd vdd FILL
X_220_ N[8] gnd _220_/Y vdd INVX1
X_279_ _305_/A _275_/CLK _275_/R vdd _199_/Y gnd vdd DFFSR
XSFILL6480x10100 gnd vdd FILL
X_150_ _185_/A _150_/B gnd _150_/Y vdd NOR2X1
X_296_ _261_/B _296_/CLK _273_/R vdd _296_/D gnd vdd DFFSR
X_202_ _209_/C gnd _203_/B vdd INVX1
XSFILL18960x14100 gnd vdd FILL
X_295_ _295_/Q _296_/CLK _273_/R vdd _295_/D gnd vdd DFFSR
X_201_ N[5] N[6] gnd _209_/C vdd NOR2X1
X_278_ _304_/A _275_/CLK _275_/R vdd _278_/D gnd vdd DFFSR
XSFILL19120x14100 gnd vdd FILL
.ends

