VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO map9v3
  CLASS BLOCK ;
  FOREIGN map9v3 ;
  ORIGIN 3.500 2.300 ;
  SIZE 261.400 BY 188.600 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.400 180.400 254.000 181.600 ;
        RECT 2.800 175.800 3.600 180.400 ;
        RECT 6.000 177.800 6.800 180.400 ;
        RECT 12.400 175.800 13.200 180.400 ;
        RECT 23.600 177.800 24.400 180.400 ;
        RECT 26.800 177.800 27.600 180.400 ;
        RECT 36.400 175.800 37.200 180.400 ;
        RECT 41.200 177.800 42.000 180.400 ;
        RECT 44.400 177.800 45.200 180.400 ;
        RECT 46.000 177.800 46.800 180.400 ;
        RECT 50.200 175.800 51.000 180.400 ;
        RECT 54.000 175.800 54.800 180.400 ;
        RECT 66.800 175.800 67.600 180.400 ;
        RECT 76.400 177.800 77.200 180.400 ;
        RECT 79.600 177.800 80.400 180.400 ;
        RECT 90.800 175.800 91.600 180.400 ;
        RECT 97.200 177.800 98.000 180.400 ;
        RECT 100.400 175.800 101.200 180.400 ;
        RECT 105.200 175.800 106.000 180.400 ;
        RECT 108.400 177.800 109.200 180.400 ;
        RECT 114.800 175.800 115.600 180.400 ;
        RECT 126.000 177.800 126.800 180.400 ;
        RECT 129.200 177.800 130.000 180.400 ;
        RECT 138.800 175.800 139.600 180.400 ;
        RECT 145.200 175.800 146.000 180.400 ;
        RECT 150.000 175.800 150.800 180.400 ;
        RECT 156.400 175.800 157.200 180.400 ;
        RECT 166.000 177.800 166.800 180.400 ;
        RECT 169.200 177.800 170.000 180.400 ;
        RECT 180.400 175.800 181.200 180.400 ;
        RECT 186.800 177.800 187.600 180.400 ;
        RECT 196.400 175.800 197.200 180.400 ;
        RECT 202.800 175.800 203.600 180.400 ;
        RECT 212.400 177.800 213.200 180.400 ;
        RECT 215.600 177.800 216.400 180.400 ;
        RECT 226.800 175.800 227.600 180.400 ;
        RECT 233.200 177.800 234.000 180.400 ;
        RECT 236.400 175.800 237.200 180.400 ;
        RECT 239.600 177.800 240.400 180.400 ;
        RECT 242.800 177.800 243.600 180.400 ;
        RECT 247.600 175.800 248.400 180.400 ;
        RECT 250.800 175.800 251.600 180.400 ;
        RECT 2.800 141.600 3.600 146.200 ;
        RECT 6.000 141.600 6.800 144.200 ;
        RECT 12.400 141.600 13.200 146.200 ;
        RECT 23.600 141.600 24.400 144.200 ;
        RECT 26.800 141.600 27.600 144.200 ;
        RECT 36.400 141.600 37.200 146.200 ;
        RECT 41.200 141.600 42.000 144.200 ;
        RECT 47.600 141.600 48.400 146.200 ;
        RECT 57.200 141.600 58.000 144.200 ;
        RECT 60.400 141.600 61.200 144.200 ;
        RECT 71.600 141.600 72.400 146.200 ;
        RECT 78.000 141.600 78.800 144.200 ;
        RECT 86.600 141.600 87.400 146.200 ;
        RECT 90.800 141.600 91.600 144.200 ;
        RECT 92.400 141.600 93.200 144.200 ;
        RECT 95.600 141.600 96.400 144.200 ;
        RECT 97.800 141.600 98.600 146.200 ;
        RECT 102.000 141.600 102.800 144.200 ;
        RECT 105.200 141.600 106.000 146.200 ;
        RECT 108.400 141.600 109.200 144.200 ;
        RECT 111.600 141.600 112.400 144.200 ;
        RECT 114.800 141.600 115.600 146.200 ;
        RECT 118.000 141.600 118.800 144.200 ;
        RECT 121.200 141.600 122.000 144.200 ;
        RECT 122.800 141.600 123.600 144.200 ;
        RECT 127.000 141.600 127.800 146.200 ;
        RECT 130.800 141.600 131.600 144.200 ;
        RECT 134.000 141.600 134.800 146.200 ;
        RECT 137.200 141.600 138.000 146.200 ;
        RECT 145.200 141.600 146.000 146.200 ;
        RECT 154.800 141.600 155.600 144.200 ;
        RECT 158.000 141.600 158.800 144.200 ;
        RECT 169.200 141.600 170.000 146.200 ;
        RECT 175.600 141.600 176.400 144.200 ;
        RECT 178.800 141.600 179.600 146.200 ;
        RECT 183.600 141.600 184.400 145.400 ;
        RECT 198.000 141.600 198.800 146.200 ;
        RECT 199.600 141.600 200.400 144.200 ;
        RECT 202.800 141.600 203.600 144.200 ;
        RECT 207.600 141.600 208.400 146.200 ;
        RECT 210.800 141.600 211.600 145.400 ;
        RECT 218.800 141.600 219.600 146.200 ;
        RECT 222.000 142.200 223.000 145.600 ;
        RECT 222.200 141.600 223.000 142.200 ;
        RECT 228.200 141.600 229.200 145.600 ;
        RECT 233.200 141.600 234.000 145.400 ;
        RECT 239.600 141.600 240.400 145.400 ;
        RECT 246.000 141.600 246.800 144.200 ;
        RECT 247.600 141.600 248.400 144.200 ;
        RECT 250.800 141.600 251.600 144.200 ;
        RECT 0.400 140.400 254.000 141.600 ;
        RECT 2.800 135.800 3.600 140.400 ;
        RECT 6.000 137.800 6.800 140.400 ;
        RECT 12.400 135.800 13.200 140.400 ;
        RECT 23.600 137.800 24.400 140.400 ;
        RECT 26.800 137.800 27.600 140.400 ;
        RECT 36.400 135.800 37.200 140.400 ;
        RECT 41.200 137.800 42.000 140.400 ;
        RECT 46.000 136.600 46.800 140.400 ;
        RECT 54.000 136.600 54.800 140.400 ;
        RECT 62.000 137.800 62.800 140.400 ;
        RECT 71.600 136.600 72.400 140.400 ;
        RECT 79.600 135.800 80.400 140.400 ;
        RECT 86.000 135.800 86.800 140.400 ;
        RECT 95.600 137.800 96.400 140.400 ;
        RECT 98.800 137.800 99.600 140.400 ;
        RECT 110.000 135.800 110.800 140.400 ;
        RECT 116.400 137.800 117.200 140.400 ;
        RECT 118.000 137.800 118.800 140.400 ;
        RECT 124.400 135.800 125.200 140.400 ;
        RECT 135.600 137.800 136.400 140.400 ;
        RECT 138.800 137.800 139.600 140.400 ;
        RECT 148.400 135.800 149.200 140.400 ;
        RECT 153.200 135.800 154.000 140.400 ;
        RECT 156.400 135.800 157.200 140.400 ;
        RECT 158.600 135.800 159.400 140.400 ;
        RECT 162.800 137.800 163.600 140.400 ;
        RECT 169.200 136.600 170.000 140.400 ;
        RECT 172.400 135.800 173.200 140.400 ;
        RECT 175.600 135.800 176.400 140.400 ;
        RECT 178.800 136.600 179.600 140.400 ;
        RECT 190.600 135.800 191.400 140.400 ;
        RECT 194.800 137.800 195.600 140.400 ;
        RECT 196.400 137.800 197.200 140.400 ;
        RECT 199.600 137.800 200.400 140.400 ;
        RECT 202.800 136.600 203.600 140.400 ;
        RECT 210.800 136.600 211.600 140.400 ;
        RECT 215.600 137.800 216.400 140.400 ;
        RECT 217.200 137.800 218.000 140.400 ;
        RECT 221.400 135.800 222.200 140.400 ;
        RECT 223.600 137.800 224.400 140.400 ;
        RECT 226.800 135.800 227.600 140.400 ;
        RECT 233.200 136.600 234.000 140.400 ;
        RECT 238.000 137.800 238.800 140.400 ;
        RECT 241.200 137.800 242.000 140.400 ;
        RECT 244.400 133.800 245.200 140.400 ;
        RECT 2.800 101.600 3.600 106.200 ;
        RECT 6.000 101.600 6.800 104.200 ;
        RECT 12.400 101.600 13.200 106.200 ;
        RECT 23.600 101.600 24.400 104.200 ;
        RECT 26.800 101.600 27.600 104.200 ;
        RECT 36.400 101.600 37.200 106.200 ;
        RECT 41.800 101.600 42.600 106.200 ;
        RECT 46.000 101.600 46.800 104.200 ;
        RECT 47.600 101.600 48.400 104.200 ;
        RECT 50.800 101.600 51.600 104.200 ;
        RECT 54.000 101.600 54.800 105.400 ;
        RECT 61.400 101.600 62.200 106.000 ;
        RECT 73.200 101.600 74.000 106.200 ;
        RECT 78.000 101.600 79.000 105.600 ;
        RECT 84.200 102.200 85.200 105.600 ;
        RECT 84.200 101.600 85.000 102.200 ;
        RECT 92.400 101.600 93.200 105.400 ;
        RECT 98.800 101.600 99.600 106.200 ;
        RECT 108.400 101.600 109.200 104.200 ;
        RECT 111.600 101.600 112.400 104.200 ;
        RECT 122.800 101.600 123.600 106.200 ;
        RECT 129.200 101.600 130.000 104.200 ;
        RECT 133.000 101.600 133.800 106.000 ;
        RECT 140.400 101.600 141.200 105.400 ;
        RECT 145.200 101.600 146.000 105.400 ;
        RECT 154.800 101.600 155.600 105.400 ;
        RECT 158.000 101.600 158.800 104.200 ;
        RECT 162.200 101.600 163.000 106.200 ;
        RECT 167.600 101.600 168.400 105.400 ;
        RECT 170.800 101.600 171.600 104.200 ;
        RECT 174.000 101.600 174.800 104.200 ;
        RECT 175.600 101.600 176.400 104.200 ;
        RECT 178.800 101.600 179.600 104.200 ;
        RECT 182.000 101.600 182.800 104.200 ;
        RECT 190.400 101.600 191.200 106.200 ;
        RECT 196.400 101.600 197.200 106.200 ;
        RECT 198.000 101.600 198.800 104.200 ;
        RECT 201.200 101.600 202.000 104.200 ;
        RECT 206.000 101.600 206.800 105.400 ;
        RECT 212.400 101.600 213.200 106.200 ;
        RECT 222.000 101.600 222.800 104.200 ;
        RECT 225.200 101.600 226.000 104.200 ;
        RECT 236.400 101.600 237.200 106.200 ;
        RECT 242.800 101.600 243.600 104.200 ;
        RECT 246.000 101.600 246.800 105.400 ;
        RECT 0.400 100.400 254.000 101.600 ;
        RECT 2.800 95.800 3.600 100.400 ;
        RECT 6.000 97.800 6.800 100.400 ;
        RECT 12.400 95.800 13.200 100.400 ;
        RECT 23.600 97.800 24.400 100.400 ;
        RECT 26.800 97.800 27.600 100.400 ;
        RECT 36.400 95.800 37.200 100.400 ;
        RECT 46.000 96.600 46.800 100.400 ;
        RECT 50.800 96.400 51.800 100.400 ;
        RECT 57.000 99.800 57.800 100.400 ;
        RECT 57.000 96.400 58.000 99.800 ;
        RECT 60.400 97.800 61.200 100.400 ;
        RECT 74.800 96.600 75.600 100.400 ;
        RECT 79.600 97.800 80.400 100.400 ;
        RECT 81.200 97.800 82.000 100.400 ;
        RECT 87.600 95.800 88.400 100.400 ;
        RECT 98.800 97.800 99.600 100.400 ;
        RECT 102.000 97.800 102.800 100.400 ;
        RECT 111.600 95.800 112.400 100.400 ;
        RECT 119.600 95.800 120.400 100.400 ;
        RECT 129.200 97.800 130.000 100.400 ;
        RECT 132.400 97.800 133.200 100.400 ;
        RECT 143.600 95.800 144.400 100.400 ;
        RECT 150.000 97.800 150.800 100.400 ;
        RECT 154.800 96.600 155.600 100.400 ;
        RECT 158.000 97.800 158.800 100.400 ;
        RECT 161.200 97.800 162.000 100.400 ;
        RECT 164.400 97.800 165.200 100.400 ;
        RECT 166.000 97.800 166.800 100.400 ;
        RECT 169.200 97.800 170.000 100.400 ;
        RECT 170.800 97.800 171.600 100.400 ;
        RECT 174.000 97.800 174.800 100.400 ;
        RECT 178.800 95.800 179.600 100.400 ;
        RECT 180.400 97.800 181.200 100.400 ;
        RECT 190.000 93.800 190.800 100.400 ;
        RECT 199.600 95.800 200.400 100.400 ;
        RECT 202.800 96.600 203.600 100.400 ;
        RECT 210.800 96.600 211.600 100.400 ;
        RECT 217.200 95.800 218.000 100.400 ;
        RECT 218.800 97.800 219.600 100.400 ;
        RECT 222.000 97.800 222.800 100.400 ;
        RECT 224.200 95.800 225.000 100.400 ;
        RECT 228.400 97.800 229.200 100.400 ;
        RECT 232.200 96.000 233.000 100.400 ;
        RECT 238.000 97.800 238.800 100.400 ;
        RECT 242.800 96.600 243.600 100.400 ;
        RECT 246.000 97.800 246.800 100.400 ;
        RECT 250.200 95.800 251.000 100.400 ;
        RECT 2.800 61.600 3.600 66.200 ;
        RECT 6.000 61.600 6.800 66.200 ;
        RECT 9.200 61.600 10.000 66.200 ;
        RECT 12.400 61.600 13.200 66.200 ;
        RECT 15.600 61.600 16.400 66.200 ;
        RECT 18.800 61.600 19.600 66.200 ;
        RECT 20.400 61.600 21.200 66.200 ;
        RECT 23.600 61.600 24.400 66.200 ;
        RECT 26.800 61.600 27.600 66.200 ;
        RECT 30.000 61.600 30.800 66.200 ;
        RECT 33.200 61.600 34.000 66.200 ;
        RECT 34.800 61.600 35.600 64.200 ;
        RECT 39.600 61.600 40.400 65.400 ;
        RECT 50.800 61.600 51.600 65.400 ;
        RECT 54.000 61.600 54.800 66.200 ;
        RECT 57.200 61.600 58.000 66.200 ;
        RECT 65.200 61.600 66.000 66.200 ;
        RECT 68.400 61.600 69.200 66.200 ;
        RECT 71.600 61.600 72.400 66.200 ;
        RECT 74.800 61.600 75.600 66.200 ;
        RECT 78.000 61.600 78.800 66.200 ;
        RECT 81.200 61.600 82.000 66.200 ;
        RECT 87.600 61.600 88.400 66.200 ;
        RECT 97.200 61.600 98.000 64.200 ;
        RECT 100.400 61.600 101.200 64.200 ;
        RECT 111.600 61.600 112.400 66.200 ;
        RECT 118.000 61.600 118.800 64.200 ;
        RECT 121.800 61.600 122.600 66.000 ;
        RECT 127.600 61.600 128.400 66.200 ;
        RECT 137.200 61.600 138.000 63.800 ;
        RECT 140.400 61.600 141.200 64.200 ;
        RECT 145.200 61.600 146.000 65.400 ;
        RECT 151.600 61.600 152.400 65.400 ;
        RECT 158.000 61.600 158.800 65.400 ;
        RECT 166.000 61.600 166.800 66.200 ;
        RECT 167.600 61.600 168.400 64.200 ;
        RECT 171.800 61.600 172.600 66.200 ;
        RECT 174.000 61.600 174.800 64.200 ;
        RECT 177.200 61.600 178.000 64.200 ;
        RECT 188.400 61.600 189.200 66.200 ;
        RECT 198.000 61.600 198.800 64.200 ;
        RECT 201.200 61.600 202.000 64.200 ;
        RECT 212.400 61.600 213.200 66.200 ;
        RECT 218.800 61.600 219.600 64.200 ;
        RECT 220.800 61.600 221.600 66.200 ;
        RECT 226.800 61.600 227.600 66.200 ;
        RECT 230.000 61.600 230.800 64.200 ;
        RECT 233.200 62.200 234.200 65.600 ;
        RECT 233.400 61.600 234.200 62.200 ;
        RECT 239.400 61.600 240.400 65.600 ;
        RECT 242.800 61.600 243.600 68.200 ;
        RECT 249.200 61.600 250.000 64.200 ;
        RECT 252.400 61.600 253.200 64.200 ;
        RECT 0.400 60.400 254.000 61.600 ;
        RECT 2.800 55.800 3.600 60.400 ;
        RECT 6.000 57.800 6.800 60.400 ;
        RECT 9.200 57.800 10.000 60.400 ;
        RECT 15.600 55.800 16.400 60.400 ;
        RECT 26.800 57.800 27.600 60.400 ;
        RECT 30.000 57.800 30.800 60.400 ;
        RECT 39.600 55.800 40.400 60.400 ;
        RECT 44.400 57.800 45.200 60.400 ;
        RECT 50.800 55.800 51.600 60.400 ;
        RECT 62.000 57.800 62.800 60.400 ;
        RECT 65.200 57.800 66.000 60.400 ;
        RECT 74.800 55.800 75.600 60.400 ;
        RECT 87.600 55.800 88.400 60.400 ;
        RECT 92.400 55.800 93.200 60.400 ;
        RECT 97.200 55.800 98.000 60.400 ;
        RECT 100.400 57.800 101.200 60.400 ;
        RECT 103.600 57.800 104.400 60.400 ;
        RECT 108.400 55.800 109.200 60.400 ;
        RECT 118.000 57.800 118.800 60.400 ;
        RECT 121.200 57.800 122.000 60.400 ;
        RECT 132.400 55.800 133.200 60.400 ;
        RECT 138.800 57.800 139.600 60.400 ;
        RECT 142.000 57.800 142.800 60.400 ;
        RECT 146.800 55.800 147.600 60.400 ;
        RECT 148.400 57.800 149.200 60.400 ;
        RECT 151.600 57.800 152.400 60.400 ;
        RECT 158.000 55.800 158.800 60.400 ;
        RECT 169.200 57.800 170.000 60.400 ;
        RECT 172.400 57.800 173.200 60.400 ;
        RECT 182.000 55.800 182.800 60.400 ;
        RECT 193.200 55.800 194.000 60.400 ;
        RECT 202.800 53.800 203.600 60.400 ;
        RECT 204.400 55.800 205.200 60.400 ;
        RECT 212.400 55.800 213.200 60.400 ;
        RECT 222.000 57.800 222.800 60.400 ;
        RECT 225.200 57.800 226.000 60.400 ;
        RECT 236.400 55.800 237.200 60.400 ;
        RECT 242.800 57.800 243.600 60.400 ;
        RECT 246.000 55.800 246.800 60.400 ;
        RECT 252.400 55.800 253.200 60.400 ;
        RECT 2.800 21.600 3.600 26.200 ;
        RECT 6.000 21.600 6.800 24.200 ;
        RECT 12.400 21.600 13.200 26.200 ;
        RECT 23.600 21.600 24.400 24.200 ;
        RECT 26.800 21.600 27.600 24.200 ;
        RECT 36.400 21.600 37.200 26.200 ;
        RECT 41.200 21.600 42.000 24.200 ;
        RECT 45.400 21.600 46.200 26.200 ;
        RECT 47.600 21.600 48.400 24.200 ;
        RECT 50.800 21.600 51.600 24.200 ;
        RECT 54.000 21.600 54.800 26.200 ;
        RECT 66.800 21.600 67.600 26.200 ;
        RECT 76.400 21.600 77.200 24.200 ;
        RECT 79.600 21.600 80.400 24.200 ;
        RECT 90.800 21.600 91.600 26.200 ;
        RECT 97.200 21.600 98.000 24.200 ;
        RECT 98.800 21.600 99.600 24.200 ;
        RECT 102.000 21.600 102.800 24.200 ;
        RECT 103.600 21.600 104.400 24.200 ;
        RECT 107.800 21.600 108.600 26.200 ;
        RECT 110.000 21.600 110.800 26.200 ;
        RECT 113.200 21.600 114.000 26.200 ;
        RECT 116.400 21.600 117.200 26.200 ;
        RECT 119.600 21.600 120.400 26.200 ;
        RECT 122.800 21.600 123.600 26.200 ;
        RECT 127.600 21.600 128.400 26.200 ;
        RECT 129.200 21.600 130.000 26.200 ;
        RECT 132.400 21.600 133.200 26.200 ;
        RECT 135.600 21.600 136.400 26.200 ;
        RECT 138.800 21.600 139.600 26.200 ;
        RECT 142.000 21.600 142.800 26.200 ;
        RECT 145.200 21.600 146.000 26.200 ;
        RECT 151.600 21.600 152.400 26.200 ;
        RECT 161.200 21.600 162.000 24.200 ;
        RECT 164.400 21.600 165.200 24.200 ;
        RECT 175.600 21.600 176.400 26.200 ;
        RECT 182.000 21.600 182.800 24.200 ;
        RECT 191.600 21.600 192.400 26.200 ;
        RECT 194.800 21.600 195.600 24.200 ;
        RECT 201.200 21.600 202.000 25.400 ;
        RECT 206.000 21.600 206.800 24.200 ;
        RECT 210.800 21.600 211.600 26.200 ;
        RECT 220.400 21.600 221.200 24.200 ;
        RECT 223.600 21.600 224.400 24.200 ;
        RECT 234.800 21.600 235.600 26.200 ;
        RECT 241.200 21.600 242.000 24.200 ;
        RECT 244.400 21.600 245.200 24.200 ;
        RECT 247.600 21.600 248.400 26.200 ;
        RECT 0.400 20.400 254.000 21.600 ;
        RECT 2.800 15.800 3.600 20.400 ;
        RECT 6.000 17.800 6.800 20.400 ;
        RECT 12.400 15.800 13.200 20.400 ;
        RECT 23.600 17.800 24.400 20.400 ;
        RECT 26.800 17.800 27.600 20.400 ;
        RECT 36.400 15.800 37.200 20.400 ;
        RECT 41.200 17.800 42.000 20.400 ;
        RECT 44.400 17.800 45.200 20.400 ;
        RECT 46.000 17.800 46.800 20.400 ;
        RECT 50.200 15.800 51.000 20.400 ;
        RECT 62.000 15.800 62.800 20.400 ;
        RECT 71.600 17.800 72.400 20.400 ;
        RECT 74.800 17.800 75.600 20.400 ;
        RECT 86.000 15.800 86.800 20.400 ;
        RECT 92.400 17.800 93.200 20.400 ;
        RECT 95.600 15.800 96.400 20.400 ;
        RECT 98.800 15.800 99.600 20.400 ;
        RECT 102.000 15.800 102.800 20.400 ;
        RECT 105.200 15.800 106.000 20.400 ;
        RECT 108.400 15.800 109.200 20.400 ;
        RECT 111.600 17.800 112.400 20.400 ;
        RECT 116.400 16.600 117.200 20.400 ;
        RECT 121.200 17.800 122.000 20.400 ;
        RECT 127.600 15.800 128.400 20.400 ;
        RECT 138.800 17.800 139.600 20.400 ;
        RECT 142.000 17.800 142.800 20.400 ;
        RECT 151.600 15.800 152.400 20.400 ;
        RECT 159.600 15.800 160.400 20.400 ;
        RECT 169.200 17.800 170.000 20.400 ;
        RECT 172.400 17.800 173.200 20.400 ;
        RECT 183.600 15.800 184.400 20.400 ;
        RECT 190.000 17.800 190.800 20.400 ;
        RECT 198.000 17.800 198.800 20.400 ;
        RECT 201.200 17.800 202.000 20.400 ;
        RECT 204.400 17.800 205.200 20.400 ;
        RECT 208.600 16.000 209.400 20.400 ;
        RECT 215.600 15.800 216.400 20.400 ;
        RECT 225.200 17.800 226.000 20.400 ;
        RECT 228.400 17.800 229.200 20.400 ;
        RECT 239.600 15.800 240.400 20.400 ;
        RECT 246.000 17.800 246.800 20.400 ;
        RECT 249.200 16.600 250.000 20.400 ;
      LAYER via1 ;
        RECT 184.300 180.600 185.100 181.400 ;
        RECT 185.300 180.600 186.100 181.400 ;
        RECT 186.300 180.600 187.100 181.400 ;
        RECT 187.300 180.600 188.100 181.400 ;
        RECT 188.300 180.600 189.100 181.400 ;
        RECT 189.300 180.600 190.100 181.400 ;
        RECT 184.300 140.600 185.100 141.400 ;
        RECT 185.300 140.600 186.100 141.400 ;
        RECT 186.300 140.600 187.100 141.400 ;
        RECT 187.300 140.600 188.100 141.400 ;
        RECT 188.300 140.600 189.100 141.400 ;
        RECT 189.300 140.600 190.100 141.400 ;
        RECT 184.300 100.600 185.100 101.400 ;
        RECT 185.300 100.600 186.100 101.400 ;
        RECT 186.300 100.600 187.100 101.400 ;
        RECT 187.300 100.600 188.100 101.400 ;
        RECT 188.300 100.600 189.100 101.400 ;
        RECT 189.300 100.600 190.100 101.400 ;
        RECT 184.300 60.600 185.100 61.400 ;
        RECT 185.300 60.600 186.100 61.400 ;
        RECT 186.300 60.600 187.100 61.400 ;
        RECT 187.300 60.600 188.100 61.400 ;
        RECT 188.300 60.600 189.100 61.400 ;
        RECT 189.300 60.600 190.100 61.400 ;
        RECT 184.300 20.600 185.100 21.400 ;
        RECT 185.300 20.600 186.100 21.400 ;
        RECT 186.300 20.600 187.100 21.400 ;
        RECT 187.300 20.600 188.100 21.400 ;
        RECT 188.300 20.600 189.100 21.400 ;
        RECT 189.300 20.600 190.100 21.400 ;
      LAYER metal2 ;
        RECT 186.600 181.400 187.800 181.600 ;
        RECT 184.300 180.600 190.100 181.400 ;
        RECT 186.600 180.400 187.800 180.600 ;
        RECT 186.600 141.400 187.800 141.600 ;
        RECT 184.300 140.600 190.100 141.400 ;
        RECT 186.600 140.400 187.800 140.600 ;
        RECT 186.600 101.400 187.800 101.600 ;
        RECT 184.300 100.600 190.100 101.400 ;
        RECT 186.600 100.400 187.800 100.600 ;
        RECT 186.600 61.400 187.800 61.600 ;
        RECT 184.300 60.600 190.100 61.400 ;
        RECT 186.600 60.400 187.800 60.600 ;
        RECT 186.600 21.400 187.800 21.600 ;
        RECT 184.300 20.600 190.100 21.400 ;
        RECT 186.600 20.400 187.800 20.600 ;
      LAYER via2 ;
        RECT 185.300 180.600 186.100 181.400 ;
        RECT 186.300 180.600 187.100 181.400 ;
        RECT 187.300 180.600 188.100 181.400 ;
        RECT 188.300 180.600 189.100 181.400 ;
        RECT 189.300 180.600 190.100 181.400 ;
        RECT 185.300 140.600 186.100 141.400 ;
        RECT 186.300 140.600 187.100 141.400 ;
        RECT 187.300 140.600 188.100 141.400 ;
        RECT 188.300 140.600 189.100 141.400 ;
        RECT 189.300 140.600 190.100 141.400 ;
        RECT 185.300 100.600 186.100 101.400 ;
        RECT 186.300 100.600 187.100 101.400 ;
        RECT 187.300 100.600 188.100 101.400 ;
        RECT 188.300 100.600 189.100 101.400 ;
        RECT 189.300 100.600 190.100 101.400 ;
        RECT 185.300 60.600 186.100 61.400 ;
        RECT 186.300 60.600 187.100 61.400 ;
        RECT 187.300 60.600 188.100 61.400 ;
        RECT 188.300 60.600 189.100 61.400 ;
        RECT 189.300 60.600 190.100 61.400 ;
        RECT 185.300 20.600 186.100 21.400 ;
        RECT 186.300 20.600 187.100 21.400 ;
        RECT 187.300 20.600 188.100 21.400 ;
        RECT 188.300 20.600 189.100 21.400 ;
        RECT 189.300 20.600 190.100 21.400 ;
      LAYER metal3 ;
        RECT 184.200 180.400 190.200 181.600 ;
        RECT 184.200 140.400 190.200 141.600 ;
        RECT 184.200 100.400 190.200 101.600 ;
        RECT 184.200 60.400 190.200 61.600 ;
        RECT 184.200 20.400 190.200 21.600 ;
      LAYER via3 ;
        RECT 184.400 180.600 185.200 181.400 ;
        RECT 185.600 180.600 186.400 181.400 ;
        RECT 186.800 180.600 187.600 181.400 ;
        RECT 188.000 180.600 188.800 181.400 ;
        RECT 189.200 180.600 190.000 181.400 ;
        RECT 184.400 140.600 185.200 141.400 ;
        RECT 185.600 140.600 186.400 141.400 ;
        RECT 186.800 140.600 187.600 141.400 ;
        RECT 188.000 140.600 188.800 141.400 ;
        RECT 189.200 140.600 190.000 141.400 ;
        RECT 184.400 100.600 185.200 101.400 ;
        RECT 185.600 100.600 186.400 101.400 ;
        RECT 186.800 100.600 187.600 101.400 ;
        RECT 188.000 100.600 188.800 101.400 ;
        RECT 189.200 100.600 190.000 101.400 ;
        RECT 184.400 60.600 185.200 61.400 ;
        RECT 185.600 60.600 186.400 61.400 ;
        RECT 186.800 60.600 187.600 61.400 ;
        RECT 188.000 60.600 188.800 61.400 ;
        RECT 189.200 60.600 190.000 61.400 ;
        RECT 184.400 20.600 185.200 21.400 ;
        RECT 185.600 20.600 186.400 21.400 ;
        RECT 186.800 20.600 187.600 21.400 ;
        RECT 188.000 20.600 188.800 21.400 ;
        RECT 189.200 20.600 190.000 21.400 ;
      LAYER metal4 ;
        RECT 184.000 -1.000 190.400 181.600 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 10.200 170.800 11.000 171.000 ;
        RECT 93.000 170.800 93.800 171.000 ;
        RECT 10.200 170.200 37.200 170.800 ;
        RECT 66.800 170.200 93.800 170.800 ;
        RECT 112.600 170.800 113.400 171.000 ;
        RECT 182.600 170.800 183.400 171.000 ;
        RECT 229.000 170.800 229.800 171.000 ;
        RECT 112.600 170.200 139.600 170.800 ;
        RECT 33.000 170.000 33.800 170.200 ;
        RECT 36.400 169.600 37.200 170.200 ;
        RECT 2.800 161.600 3.600 169.000 ;
        RECT 6.000 161.600 6.800 166.200 ;
        RECT 9.200 161.600 10.000 166.200 ;
        RECT 12.400 161.600 13.200 166.200 ;
        RECT 15.600 161.600 16.400 166.200 ;
        RECT 23.600 161.600 24.400 166.200 ;
        RECT 26.800 161.600 27.600 166.200 ;
        RECT 33.200 161.600 34.000 166.200 ;
        RECT 36.400 161.600 37.200 166.200 ;
        RECT 39.600 161.600 40.400 166.200 ;
        RECT 41.200 161.600 42.000 170.200 ;
        RECT 66.800 169.600 67.600 170.200 ;
        RECT 70.000 170.000 71.000 170.200 ;
        RECT 135.400 170.000 136.400 170.200 ;
        RECT 138.800 169.600 139.600 170.200 ;
        RECT 156.400 170.200 183.400 170.800 ;
        RECT 202.800 170.200 229.800 170.800 ;
        RECT 156.400 169.600 157.200 170.200 ;
        RECT 159.600 170.000 160.600 170.200 ;
        RECT 202.800 169.600 203.600 170.200 ;
        RECT 206.200 170.000 207.000 170.200 ;
        RECT 49.200 161.600 50.000 169.000 ;
        RECT 54.000 161.600 54.800 169.000 ;
        RECT 63.600 161.600 64.400 166.200 ;
        RECT 66.800 161.600 67.600 166.200 ;
        RECT 70.000 161.600 70.800 166.200 ;
        RECT 76.400 161.600 77.200 166.200 ;
        RECT 79.600 161.600 80.400 166.200 ;
        RECT 87.600 161.600 88.400 166.200 ;
        RECT 90.800 161.600 91.600 166.200 ;
        RECT 94.000 161.600 94.800 166.200 ;
        RECT 97.200 161.600 98.000 166.200 ;
        RECT 100.400 161.600 101.200 169.000 ;
        RECT 105.200 161.600 106.000 169.000 ;
        RECT 108.400 161.600 109.200 166.200 ;
        RECT 111.600 161.600 112.400 166.200 ;
        RECT 114.800 161.600 115.600 166.200 ;
        RECT 118.000 161.600 118.800 166.200 ;
        RECT 126.000 161.600 126.800 166.200 ;
        RECT 129.200 161.600 130.000 166.200 ;
        RECT 135.600 161.600 136.400 166.200 ;
        RECT 138.800 161.600 139.600 166.200 ;
        RECT 142.000 161.600 142.800 166.200 ;
        RECT 145.200 161.600 146.000 169.000 ;
        RECT 150.000 161.600 150.800 169.000 ;
        RECT 153.200 161.600 154.000 166.200 ;
        RECT 156.400 161.600 157.200 166.200 ;
        RECT 159.600 161.600 160.400 166.200 ;
        RECT 166.000 161.600 166.800 166.200 ;
        RECT 169.200 161.600 170.000 166.200 ;
        RECT 177.200 161.600 178.000 166.200 ;
        RECT 180.400 161.600 181.200 166.200 ;
        RECT 183.600 161.600 184.400 166.200 ;
        RECT 186.800 161.600 187.600 166.200 ;
        RECT 196.400 161.600 197.200 169.000 ;
        RECT 199.600 161.600 200.400 166.200 ;
        RECT 202.800 161.600 203.600 166.200 ;
        RECT 206.000 161.600 206.800 166.200 ;
        RECT 212.400 161.600 213.200 166.200 ;
        RECT 215.600 161.600 216.400 166.200 ;
        RECT 223.600 161.600 224.400 166.200 ;
        RECT 226.800 161.600 227.600 166.200 ;
        RECT 230.000 161.600 230.800 166.200 ;
        RECT 233.200 161.600 234.000 166.200 ;
        RECT 236.400 161.600 237.200 169.000 ;
        RECT 239.600 161.600 240.400 170.200 ;
        RECT 244.400 161.600 245.200 166.200 ;
        RECT 247.600 161.600 248.400 166.200 ;
        RECT 250.800 161.600 251.600 169.000 ;
        RECT 0.400 160.400 254.000 161.600 ;
        RECT 2.800 153.000 3.600 160.400 ;
        RECT 6.000 155.800 6.800 160.400 ;
        RECT 9.200 155.800 10.000 160.400 ;
        RECT 12.400 155.800 13.200 160.400 ;
        RECT 15.600 155.800 16.400 160.400 ;
        RECT 23.600 155.800 24.400 160.400 ;
        RECT 26.800 155.800 27.600 160.400 ;
        RECT 33.200 155.800 34.000 160.400 ;
        RECT 36.400 155.800 37.200 160.400 ;
        RECT 39.600 155.800 40.400 160.400 ;
        RECT 41.200 155.800 42.000 160.400 ;
        RECT 44.400 155.800 45.200 160.400 ;
        RECT 47.600 155.800 48.400 160.400 ;
        RECT 50.800 155.800 51.600 160.400 ;
        RECT 57.200 155.800 58.000 160.400 ;
        RECT 60.400 155.800 61.200 160.400 ;
        RECT 68.400 155.800 69.200 160.400 ;
        RECT 71.600 155.800 72.400 160.400 ;
        RECT 74.800 155.800 75.600 160.400 ;
        RECT 78.000 155.800 78.800 160.400 ;
        RECT 87.600 153.000 88.400 160.400 ;
        RECT 33.000 151.800 33.800 152.000 ;
        RECT 36.400 151.800 37.200 152.400 ;
        RECT 10.200 151.200 37.200 151.800 ;
        RECT 47.600 151.800 48.400 152.400 ;
        RECT 51.000 151.800 51.800 152.000 ;
        RECT 92.400 151.800 93.200 160.400 ;
        RECT 98.800 153.000 99.600 160.400 ;
        RECT 105.200 153.000 106.000 160.400 ;
        RECT 111.600 151.800 112.400 160.400 ;
        RECT 114.800 153.000 115.600 160.400 ;
        RECT 118.000 151.800 118.800 160.400 ;
        RECT 126.000 153.000 126.800 160.400 ;
        RECT 130.800 155.800 131.600 160.400 ;
        RECT 134.000 153.000 134.800 160.400 ;
        RECT 137.200 155.800 138.000 160.400 ;
        RECT 140.400 155.800 141.200 160.400 ;
        RECT 142.000 155.800 142.800 160.400 ;
        RECT 145.200 155.800 146.000 160.400 ;
        RECT 148.400 155.800 149.200 160.400 ;
        RECT 154.800 155.800 155.600 160.400 ;
        RECT 158.000 155.800 158.800 160.400 ;
        RECT 166.000 155.800 166.800 160.400 ;
        RECT 169.200 155.800 170.000 160.400 ;
        RECT 172.400 155.800 173.200 160.400 ;
        RECT 175.600 155.800 176.400 160.400 ;
        RECT 178.800 153.000 179.600 160.400 ;
        RECT 145.200 151.800 146.000 152.400 ;
        RECT 148.400 151.800 149.400 152.000 ;
        RECT 182.000 151.800 182.800 160.400 ;
        RECT 186.200 155.800 187.000 160.400 ;
        RECT 194.800 155.800 195.600 160.400 ;
        RECT 198.000 155.800 198.800 160.400 ;
        RECT 199.600 151.800 200.400 160.400 ;
        RECT 204.400 155.800 205.200 160.400 ;
        RECT 207.600 155.800 208.400 160.400 ;
        RECT 209.200 151.800 210.000 160.400 ;
        RECT 213.400 155.800 214.200 160.400 ;
        RECT 215.600 155.800 216.400 160.400 ;
        RECT 218.800 155.800 219.600 160.400 ;
        RECT 222.200 159.800 223.000 160.400 ;
        RECT 222.000 153.200 223.000 159.800 ;
        RECT 228.200 153.200 229.200 160.400 ;
        RECT 231.600 151.800 232.400 160.400 ;
        RECT 235.800 155.800 236.600 160.400 ;
        RECT 238.000 151.800 238.800 160.400 ;
        RECT 242.200 155.800 243.000 160.400 ;
        RECT 246.000 155.800 246.800 160.400 ;
        RECT 247.600 151.800 248.400 160.400 ;
        RECT 47.600 151.200 74.600 151.800 ;
        RECT 145.200 151.200 172.200 151.800 ;
        RECT 10.200 151.000 11.000 151.200 ;
        RECT 73.800 151.000 74.600 151.200 ;
        RECT 171.400 151.000 172.200 151.200 ;
        RECT 10.200 130.800 11.000 131.000 ;
        RECT 112.200 130.800 113.000 131.000 ;
        RECT 10.200 130.200 37.200 130.800 ;
        RECT 86.000 130.200 113.000 130.800 ;
        RECT 122.200 130.800 123.000 131.000 ;
        RECT 122.200 130.200 149.200 130.800 ;
        RECT 33.000 130.000 33.800 130.200 ;
        RECT 36.400 129.600 37.200 130.200 ;
        RECT 2.800 121.600 3.600 129.000 ;
        RECT 6.000 121.600 6.800 126.200 ;
        RECT 9.200 121.600 10.000 126.200 ;
        RECT 12.400 121.600 13.200 126.200 ;
        RECT 15.600 121.600 16.400 126.200 ;
        RECT 23.600 121.600 24.400 126.200 ;
        RECT 26.800 121.600 27.600 126.200 ;
        RECT 33.200 121.600 34.000 126.200 ;
        RECT 36.400 121.600 37.200 126.200 ;
        RECT 39.600 121.600 40.400 126.200 ;
        RECT 41.200 121.600 42.000 126.200 ;
        RECT 44.400 121.600 45.200 130.200 ;
        RECT 50.800 121.600 51.600 130.200 ;
        RECT 52.400 121.600 53.200 130.200 ;
        RECT 58.800 121.600 59.600 130.200 ;
        RECT 62.000 121.600 62.800 126.200 ;
        RECT 70.000 121.600 70.800 130.200 ;
        RECT 76.400 121.600 77.200 130.200 ;
        RECT 86.000 129.600 86.800 130.200 ;
        RECT 89.200 130.000 90.200 130.200 ;
        RECT 145.000 130.000 146.000 130.200 ;
        RECT 148.400 129.600 149.200 130.200 ;
        RECT 79.600 121.600 80.400 129.000 ;
        RECT 82.800 121.600 83.600 126.200 ;
        RECT 86.000 121.600 86.800 126.200 ;
        RECT 89.200 121.600 90.000 126.200 ;
        RECT 95.600 121.600 96.400 126.200 ;
        RECT 98.800 121.600 99.600 126.200 ;
        RECT 106.800 121.600 107.600 126.200 ;
        RECT 110.000 121.600 110.800 126.200 ;
        RECT 113.200 121.600 114.000 126.200 ;
        RECT 116.400 121.600 117.200 126.200 ;
        RECT 118.000 121.600 118.800 126.200 ;
        RECT 121.200 121.600 122.000 126.200 ;
        RECT 124.400 121.600 125.200 126.200 ;
        RECT 127.600 121.600 128.400 126.200 ;
        RECT 135.600 121.600 136.400 126.200 ;
        RECT 138.800 121.600 139.600 126.200 ;
        RECT 145.200 121.600 146.000 126.200 ;
        RECT 148.400 121.600 149.200 126.200 ;
        RECT 151.600 121.600 152.400 126.200 ;
        RECT 153.200 121.600 154.000 130.200 ;
        RECT 156.400 121.600 157.200 130.200 ;
        RECT 159.600 121.600 160.400 129.000 ;
        RECT 164.400 121.600 165.200 130.200 ;
        RECT 170.800 121.600 171.600 130.200 ;
        RECT 172.400 121.600 173.200 130.200 ;
        RECT 175.600 121.600 176.400 130.200 ;
        RECT 177.200 121.600 178.000 130.200 ;
        RECT 181.400 121.600 182.200 126.200 ;
        RECT 191.600 121.600 192.400 129.000 ;
        RECT 196.400 121.600 197.200 130.200 ;
        RECT 201.200 121.600 202.000 130.200 ;
        RECT 205.400 121.600 206.200 126.200 ;
        RECT 208.200 121.600 209.000 126.200 ;
        RECT 212.400 121.600 213.200 130.200 ;
        RECT 215.600 121.600 216.400 126.200 ;
        RECT 220.400 121.600 221.200 129.000 ;
        RECT 223.600 121.600 224.400 126.200 ;
        RECT 226.800 121.600 227.600 126.200 ;
        RECT 230.000 121.600 230.800 126.200 ;
        RECT 231.600 121.600 232.400 130.200 ;
        RECT 235.800 121.600 236.600 126.200 ;
        RECT 238.000 121.600 238.800 126.200 ;
        RECT 241.200 121.600 242.000 126.200 ;
        RECT 244.400 121.600 245.200 126.200 ;
        RECT 247.600 121.600 248.400 125.800 ;
        RECT 0.400 120.400 254.000 121.600 ;
        RECT 2.800 113.000 3.600 120.400 ;
        RECT 6.000 115.800 6.800 120.400 ;
        RECT 9.200 115.800 10.000 120.400 ;
        RECT 12.400 115.800 13.200 120.400 ;
        RECT 15.600 115.800 16.400 120.400 ;
        RECT 23.600 115.800 24.400 120.400 ;
        RECT 26.800 115.800 27.600 120.400 ;
        RECT 33.200 115.800 34.000 120.400 ;
        RECT 36.400 115.800 37.200 120.400 ;
        RECT 39.600 115.800 40.400 120.400 ;
        RECT 42.800 113.000 43.600 120.400 ;
        RECT 33.000 111.800 33.800 112.000 ;
        RECT 36.400 111.800 37.200 112.400 ;
        RECT 47.600 111.800 48.400 120.400 ;
        RECT 52.400 111.800 53.200 120.400 ;
        RECT 56.600 115.800 57.400 120.400 ;
        RECT 58.800 115.800 59.600 120.400 ;
        RECT 62.000 112.200 62.800 120.400 ;
        RECT 73.200 113.000 74.000 120.400 ;
        RECT 78.000 113.200 79.000 120.400 ;
        RECT 84.200 119.800 85.000 120.400 ;
        RECT 84.200 113.200 85.200 119.800 ;
        RECT 87.600 111.800 88.400 120.400 ;
        RECT 94.000 111.800 94.800 120.400 ;
        RECT 95.600 115.800 96.400 120.400 ;
        RECT 98.800 115.800 99.600 120.400 ;
        RECT 102.000 115.800 102.800 120.400 ;
        RECT 108.400 115.800 109.200 120.400 ;
        RECT 111.600 115.800 112.400 120.400 ;
        RECT 119.600 115.800 120.400 120.400 ;
        RECT 122.800 115.800 123.600 120.400 ;
        RECT 126.000 115.800 126.800 120.400 ;
        RECT 129.200 115.800 130.000 120.400 ;
        RECT 98.800 111.800 99.600 112.400 ;
        RECT 132.400 112.200 133.200 120.400 ;
        RECT 135.600 115.800 136.400 120.400 ;
        RECT 137.800 115.800 138.600 120.400 ;
        RECT 102.200 111.800 103.000 112.000 ;
        RECT 142.000 111.800 142.800 120.400 ;
        RECT 143.600 111.800 144.400 120.400 ;
        RECT 147.800 115.800 148.600 120.400 ;
        RECT 150.000 111.800 150.800 120.400 ;
        RECT 156.400 111.800 157.200 120.400 ;
        RECT 161.200 113.000 162.000 120.400 ;
        RECT 165.000 115.800 165.800 120.400 ;
        RECT 169.200 111.800 170.000 120.400 ;
        RECT 170.800 111.800 171.600 120.400 ;
        RECT 175.600 115.800 176.400 120.400 ;
        RECT 182.000 111.800 182.800 120.400 ;
        RECT 191.600 113.000 192.400 120.400 ;
        RECT 198.000 111.800 198.800 120.400 ;
        RECT 203.400 115.800 204.200 120.400 ;
        RECT 207.600 111.800 208.400 120.400 ;
        RECT 209.200 115.800 210.000 120.400 ;
        RECT 212.400 115.800 213.200 120.400 ;
        RECT 215.600 115.800 216.400 120.400 ;
        RECT 222.000 115.800 222.800 120.400 ;
        RECT 225.200 115.800 226.000 120.400 ;
        RECT 233.200 115.800 234.000 120.400 ;
        RECT 236.400 115.800 237.200 120.400 ;
        RECT 239.600 115.800 240.400 120.400 ;
        RECT 242.800 115.800 243.600 120.400 ;
        RECT 212.400 111.800 213.200 112.400 ;
        RECT 215.600 111.800 216.600 112.000 ;
        RECT 244.400 111.800 245.200 120.400 ;
        RECT 248.600 115.800 249.400 120.400 ;
        RECT 10.200 111.200 37.200 111.800 ;
        RECT 98.800 111.200 125.800 111.800 ;
        RECT 212.400 111.200 239.400 111.800 ;
        RECT 10.200 111.000 11.000 111.200 ;
        RECT 125.000 111.000 125.800 111.200 ;
        RECT 238.600 111.000 239.400 111.200 ;
        RECT 10.200 90.800 11.000 91.000 ;
        RECT 85.400 90.800 86.200 91.000 ;
        RECT 145.800 90.800 146.600 91.000 ;
        RECT 10.200 90.200 37.200 90.800 ;
        RECT 85.400 90.200 112.400 90.800 ;
        RECT 33.000 90.000 33.800 90.200 ;
        RECT 36.400 89.600 37.200 90.200 ;
        RECT 2.800 81.600 3.600 89.000 ;
        RECT 6.000 81.600 6.800 86.200 ;
        RECT 9.200 81.600 10.000 86.200 ;
        RECT 12.400 81.600 13.200 86.200 ;
        RECT 15.600 81.600 16.400 86.200 ;
        RECT 23.600 81.600 24.400 86.200 ;
        RECT 26.800 81.600 27.600 86.200 ;
        RECT 33.200 81.600 34.000 86.200 ;
        RECT 36.400 81.600 37.200 86.200 ;
        RECT 39.600 81.600 40.400 86.200 ;
        RECT 41.200 81.600 42.000 90.200 ;
        RECT 47.600 81.600 48.400 90.200 ;
        RECT 50.800 81.600 51.800 88.800 ;
        RECT 57.000 82.200 58.000 88.800 ;
        RECT 57.000 81.600 57.800 82.200 ;
        RECT 60.400 81.600 61.200 86.200 ;
        RECT 70.000 81.600 70.800 90.200 ;
        RECT 76.400 81.600 77.200 90.200 ;
        RECT 108.200 90.000 109.000 90.200 ;
        RECT 111.600 89.600 112.400 90.200 ;
        RECT 119.600 90.200 146.600 90.800 ;
        RECT 119.600 89.600 120.400 90.200 ;
        RECT 122.800 90.000 123.800 90.200 ;
        RECT 79.600 81.600 80.400 86.200 ;
        RECT 81.200 81.600 82.000 86.200 ;
        RECT 84.400 81.600 85.200 86.200 ;
        RECT 87.600 81.600 88.400 86.200 ;
        RECT 90.800 81.600 91.600 86.200 ;
        RECT 98.800 81.600 99.600 86.200 ;
        RECT 102.000 81.600 102.800 86.200 ;
        RECT 108.400 81.600 109.200 86.200 ;
        RECT 111.600 81.600 112.400 86.200 ;
        RECT 114.800 81.600 115.600 86.200 ;
        RECT 116.400 81.600 117.200 86.200 ;
        RECT 119.600 81.600 120.400 86.200 ;
        RECT 122.800 81.600 123.600 86.200 ;
        RECT 129.200 81.600 130.000 86.200 ;
        RECT 132.400 81.600 133.200 86.200 ;
        RECT 140.400 81.600 141.200 86.200 ;
        RECT 143.600 81.600 144.400 86.200 ;
        RECT 146.800 81.600 147.600 86.200 ;
        RECT 150.000 81.600 150.800 86.200 ;
        RECT 152.200 81.600 153.000 86.200 ;
        RECT 156.400 81.600 157.200 90.200 ;
        RECT 158.000 81.600 158.800 86.200 ;
        RECT 164.400 81.600 165.200 90.200 ;
        RECT 166.000 81.600 166.800 90.200 ;
        RECT 170.800 81.600 171.600 90.200 ;
        RECT 175.600 81.600 176.400 86.200 ;
        RECT 178.800 81.600 179.600 86.200 ;
        RECT 180.400 81.600 181.200 86.200 ;
        RECT 190.000 81.600 190.800 86.200 ;
        RECT 193.200 81.600 194.000 85.800 ;
        RECT 196.400 81.600 197.200 86.200 ;
        RECT 199.600 81.600 200.400 86.200 ;
        RECT 201.200 81.600 202.000 90.200 ;
        RECT 205.400 81.600 206.200 86.200 ;
        RECT 208.200 81.600 209.000 86.200 ;
        RECT 212.400 81.600 213.200 90.200 ;
        RECT 214.000 81.600 214.800 86.200 ;
        RECT 217.200 81.600 218.000 86.200 ;
        RECT 222.000 81.600 222.800 90.200 ;
        RECT 225.200 81.600 226.000 89.000 ;
        RECT 231.600 81.600 232.400 89.800 ;
        RECT 234.800 81.600 235.600 86.200 ;
        RECT 238.000 81.600 238.800 86.200 ;
        RECT 240.200 81.600 241.000 86.200 ;
        RECT 244.400 81.600 245.200 90.200 ;
        RECT 249.200 81.600 250.000 89.000 ;
        RECT 0.400 80.400 254.000 81.600 ;
        RECT 2.800 73.000 3.600 80.400 ;
        RECT 6.000 71.800 6.800 80.400 ;
        RECT 9.200 71.800 10.000 80.400 ;
        RECT 12.400 71.800 13.200 80.400 ;
        RECT 15.600 71.800 16.400 80.400 ;
        RECT 18.800 71.800 19.600 80.400 ;
        RECT 20.400 71.800 21.200 80.400 ;
        RECT 23.600 71.800 24.400 80.400 ;
        RECT 26.800 71.800 27.600 80.400 ;
        RECT 30.000 71.800 30.800 80.400 ;
        RECT 33.200 71.800 34.000 80.400 ;
        RECT 34.800 75.800 35.600 80.400 ;
        RECT 38.000 71.800 38.800 80.400 ;
        RECT 44.400 71.800 45.200 80.400 ;
        RECT 46.000 71.800 46.800 80.400 ;
        RECT 52.400 71.800 53.200 80.400 ;
        RECT 54.000 71.800 54.800 80.400 ;
        RECT 57.200 71.800 58.000 80.400 ;
        RECT 65.200 71.800 66.000 80.400 ;
        RECT 68.400 71.800 69.200 80.400 ;
        RECT 71.600 71.800 72.400 80.400 ;
        RECT 74.800 71.800 75.600 80.400 ;
        RECT 78.000 71.800 78.800 80.400 ;
        RECT 81.200 73.000 82.000 80.400 ;
        RECT 84.400 75.800 85.200 80.400 ;
        RECT 87.600 75.800 88.400 80.400 ;
        RECT 90.800 75.800 91.600 80.400 ;
        RECT 97.200 75.800 98.000 80.400 ;
        RECT 100.400 75.800 101.200 80.400 ;
        RECT 108.400 75.800 109.200 80.400 ;
        RECT 111.600 75.800 112.400 80.400 ;
        RECT 114.800 75.800 115.600 80.400 ;
        RECT 118.000 75.800 118.800 80.400 ;
        RECT 87.600 71.800 88.400 72.400 ;
        RECT 121.200 72.200 122.000 80.400 ;
        RECT 124.400 75.800 125.200 80.400 ;
        RECT 127.600 73.000 128.400 80.400 ;
        RECT 140.400 73.800 141.200 80.400 ;
        RECT 91.000 71.800 91.800 72.000 ;
        RECT 143.600 71.800 144.400 80.400 ;
        RECT 147.800 75.800 148.600 80.400 ;
        RECT 150.000 71.800 150.800 80.400 ;
        RECT 154.200 75.800 155.000 80.400 ;
        RECT 156.400 71.800 157.200 80.400 ;
        RECT 160.600 75.800 161.400 80.400 ;
        RECT 162.800 75.800 163.600 80.400 ;
        RECT 166.000 75.800 166.800 80.400 ;
        RECT 170.800 73.000 171.600 80.400 ;
        RECT 174.000 71.800 174.800 80.400 ;
        RECT 185.200 75.800 186.000 80.400 ;
        RECT 188.400 75.800 189.200 80.400 ;
        RECT 191.600 75.800 192.400 80.400 ;
        RECT 198.000 75.800 198.800 80.400 ;
        RECT 201.200 75.800 202.000 80.400 ;
        RECT 209.200 75.800 210.000 80.400 ;
        RECT 212.400 75.800 213.200 80.400 ;
        RECT 215.600 75.800 216.400 80.400 ;
        RECT 218.800 75.800 219.600 80.400 ;
        RECT 222.000 73.000 222.800 80.400 ;
        RECT 230.000 75.800 230.800 80.400 ;
        RECT 233.400 79.800 234.200 80.400 ;
        RECT 233.200 73.200 234.200 79.800 ;
        RECT 239.400 73.200 240.400 80.400 ;
        RECT 242.800 75.800 243.600 80.400 ;
        RECT 246.000 76.200 246.800 80.400 ;
        RECT 188.400 71.800 189.200 72.400 ;
        RECT 191.600 71.800 192.600 72.000 ;
        RECT 252.400 71.800 253.200 80.400 ;
        RECT 87.600 71.200 114.600 71.800 ;
        RECT 188.400 71.200 215.400 71.800 ;
        RECT 113.800 71.000 114.600 71.200 ;
        RECT 214.600 71.000 215.400 71.200 ;
        RECT 13.400 50.800 14.200 51.000 ;
        RECT 48.600 50.800 49.400 51.000 ;
        RECT 134.600 50.800 135.400 51.000 ;
        RECT 13.400 50.200 40.400 50.800 ;
        RECT 48.600 50.200 75.600 50.800 ;
        RECT 108.400 50.200 135.400 50.800 ;
        RECT 155.800 50.800 156.600 51.000 ;
        RECT 238.600 50.800 239.400 51.000 ;
        RECT 155.800 50.200 182.800 50.800 ;
        RECT 36.200 50.000 37.000 50.200 ;
        RECT 39.600 49.600 40.400 50.200 ;
        RECT 71.400 50.000 72.200 50.200 ;
        RECT 74.800 49.600 75.600 50.200 ;
        RECT 2.800 41.600 3.600 49.000 ;
        RECT 6.000 41.600 6.800 46.200 ;
        RECT 9.200 41.600 10.000 46.200 ;
        RECT 12.400 41.600 13.200 46.200 ;
        RECT 15.600 41.600 16.400 46.200 ;
        RECT 18.800 41.600 19.600 46.200 ;
        RECT 26.800 41.600 27.600 46.200 ;
        RECT 30.000 41.600 30.800 46.200 ;
        RECT 36.400 41.600 37.200 46.200 ;
        RECT 39.600 41.600 40.400 46.200 ;
        RECT 42.800 41.600 43.600 46.200 ;
        RECT 44.400 41.600 45.200 46.200 ;
        RECT 47.600 41.600 48.400 46.200 ;
        RECT 50.800 41.600 51.600 46.200 ;
        RECT 54.000 41.600 54.800 46.200 ;
        RECT 62.000 41.600 62.800 46.200 ;
        RECT 65.200 41.600 66.000 46.200 ;
        RECT 71.600 41.600 72.400 46.200 ;
        RECT 74.800 41.600 75.600 46.200 ;
        RECT 78.000 41.600 78.800 46.200 ;
        RECT 87.600 41.600 88.400 49.000 ;
        RECT 92.400 41.600 93.200 49.000 ;
        RECT 97.200 41.600 98.000 49.000 ;
        RECT 103.600 41.600 104.400 50.200 ;
        RECT 108.400 49.600 109.200 50.200 ;
        RECT 111.600 50.000 112.600 50.200 ;
        RECT 178.600 50.000 179.600 50.200 ;
        RECT 182.000 49.600 182.800 50.200 ;
        RECT 212.400 50.200 239.400 50.800 ;
        RECT 212.400 49.600 213.200 50.200 ;
        RECT 215.600 50.000 216.600 50.200 ;
        RECT 105.200 41.600 106.000 46.200 ;
        RECT 108.400 41.600 109.200 46.200 ;
        RECT 111.600 41.600 112.400 46.200 ;
        RECT 118.000 41.600 118.800 46.200 ;
        RECT 121.200 41.600 122.000 46.200 ;
        RECT 129.200 41.600 130.000 46.200 ;
        RECT 132.400 41.600 133.200 46.200 ;
        RECT 135.600 41.600 136.400 46.200 ;
        RECT 138.800 41.600 139.600 46.200 ;
        RECT 142.000 41.600 142.800 46.200 ;
        RECT 143.600 41.600 144.400 46.200 ;
        RECT 146.800 41.600 147.600 46.200 ;
        RECT 148.400 41.600 149.200 46.200 ;
        RECT 151.600 41.600 152.400 46.200 ;
        RECT 154.800 41.600 155.600 46.200 ;
        RECT 158.000 41.600 158.800 46.200 ;
        RECT 161.200 41.600 162.000 46.200 ;
        RECT 169.200 41.600 170.000 46.200 ;
        RECT 172.400 41.600 173.200 46.200 ;
        RECT 178.800 41.600 179.600 46.200 ;
        RECT 182.000 41.600 182.800 46.200 ;
        RECT 185.200 41.600 186.000 46.200 ;
        RECT 193.200 41.600 194.000 46.200 ;
        RECT 196.400 41.600 197.200 46.200 ;
        RECT 199.600 41.600 200.400 45.800 ;
        RECT 202.800 41.600 203.600 46.200 ;
        RECT 204.400 41.600 205.200 46.200 ;
        RECT 207.600 41.600 208.400 46.200 ;
        RECT 209.200 41.600 210.000 46.200 ;
        RECT 212.400 41.600 213.200 46.200 ;
        RECT 215.600 41.600 216.400 46.200 ;
        RECT 222.000 41.600 222.800 46.200 ;
        RECT 225.200 41.600 226.000 46.200 ;
        RECT 233.200 41.600 234.000 46.200 ;
        RECT 236.400 41.600 237.200 46.200 ;
        RECT 239.600 41.600 240.400 46.200 ;
        RECT 242.800 41.600 243.600 46.200 ;
        RECT 246.000 41.600 246.800 49.000 ;
        RECT 249.200 41.600 250.000 46.200 ;
        RECT 252.400 41.600 253.200 46.200 ;
        RECT 0.400 40.400 254.000 41.600 ;
        RECT 2.800 33.000 3.600 40.400 ;
        RECT 6.000 35.800 6.800 40.400 ;
        RECT 9.200 35.800 10.000 40.400 ;
        RECT 12.400 35.800 13.200 40.400 ;
        RECT 15.600 35.800 16.400 40.400 ;
        RECT 23.600 35.800 24.400 40.400 ;
        RECT 26.800 35.800 27.600 40.400 ;
        RECT 33.200 35.800 34.000 40.400 ;
        RECT 36.400 35.800 37.200 40.400 ;
        RECT 39.600 35.800 40.400 40.400 ;
        RECT 44.400 33.000 45.200 40.400 ;
        RECT 33.000 31.800 33.800 32.000 ;
        RECT 36.400 31.800 37.200 32.400 ;
        RECT 47.600 31.800 48.400 40.400 ;
        RECT 54.000 33.000 54.800 40.400 ;
        RECT 63.600 35.800 64.400 40.400 ;
        RECT 66.800 35.800 67.600 40.400 ;
        RECT 70.000 35.800 70.800 40.400 ;
        RECT 76.400 35.800 77.200 40.400 ;
        RECT 79.600 35.800 80.400 40.400 ;
        RECT 87.600 35.800 88.400 40.400 ;
        RECT 90.800 35.800 91.600 40.400 ;
        RECT 94.000 35.800 94.800 40.400 ;
        RECT 97.200 35.800 98.000 40.400 ;
        RECT 66.800 31.800 67.600 32.400 ;
        RECT 70.000 31.800 71.000 32.000 ;
        RECT 98.800 31.800 99.600 40.400 ;
        RECT 106.800 33.000 107.600 40.400 ;
        RECT 110.000 31.800 110.800 40.400 ;
        RECT 113.200 31.800 114.000 40.400 ;
        RECT 116.400 31.800 117.200 40.400 ;
        RECT 119.600 31.800 120.400 40.400 ;
        RECT 122.800 31.800 123.600 40.400 ;
        RECT 124.400 35.800 125.200 40.400 ;
        RECT 127.600 35.800 128.400 40.400 ;
        RECT 129.200 31.800 130.000 40.400 ;
        RECT 132.400 31.800 133.200 40.400 ;
        RECT 135.600 31.800 136.400 40.400 ;
        RECT 138.800 31.800 139.600 40.400 ;
        RECT 142.000 31.800 142.800 40.400 ;
        RECT 145.200 33.000 146.000 40.400 ;
        RECT 148.400 35.800 149.200 40.400 ;
        RECT 151.600 35.800 152.400 40.400 ;
        RECT 154.800 35.800 155.600 40.400 ;
        RECT 161.200 35.800 162.000 40.400 ;
        RECT 164.400 35.800 165.200 40.400 ;
        RECT 172.400 35.800 173.200 40.400 ;
        RECT 175.600 35.800 176.400 40.400 ;
        RECT 178.800 35.800 179.600 40.400 ;
        RECT 182.000 35.800 182.800 40.400 ;
        RECT 191.600 33.000 192.400 40.400 ;
        RECT 194.800 35.800 195.600 40.400 ;
        RECT 198.600 35.800 199.400 40.400 ;
        RECT 151.600 31.800 152.400 32.400 ;
        RECT 155.000 31.800 155.800 32.000 ;
        RECT 202.800 31.800 203.600 40.400 ;
        RECT 206.000 35.800 206.800 40.400 ;
        RECT 207.600 35.800 208.400 40.400 ;
        RECT 210.800 35.800 211.600 40.400 ;
        RECT 214.000 35.800 214.800 40.400 ;
        RECT 220.400 35.600 221.200 40.400 ;
        RECT 223.600 35.800 224.400 40.400 ;
        RECT 231.600 35.800 232.400 40.400 ;
        RECT 234.800 35.800 235.600 40.400 ;
        RECT 238.000 35.800 238.800 40.400 ;
        RECT 241.200 35.800 242.000 40.400 ;
        RECT 244.400 35.800 245.200 40.400 ;
        RECT 247.600 33.000 248.400 40.400 ;
        RECT 10.200 31.200 37.200 31.800 ;
        RECT 66.800 31.200 93.800 31.800 ;
        RECT 151.600 31.200 178.600 31.800 ;
        RECT 10.200 31.000 11.000 31.200 ;
        RECT 93.000 31.000 93.800 31.200 ;
        RECT 177.800 31.000 178.600 31.200 ;
        RECT 209.000 30.000 232.400 30.600 ;
        RECT 209.000 29.800 209.800 30.000 ;
        RECT 214.000 29.600 214.800 30.000 ;
        RECT 220.400 29.600 221.200 30.000 ;
        RECT 231.600 29.400 232.400 30.000 ;
        RECT 10.200 10.800 11.000 11.000 ;
        RECT 88.200 10.800 89.000 11.000 ;
        RECT 10.200 10.200 37.200 10.800 ;
        RECT 62.000 10.200 89.000 10.800 ;
        RECT 125.400 10.800 126.200 11.000 ;
        RECT 185.800 10.800 186.600 11.000 ;
        RECT 241.800 10.800 242.600 11.000 ;
        RECT 125.400 10.200 152.400 10.800 ;
        RECT 33.000 10.000 34.000 10.200 ;
        RECT 36.400 9.600 37.200 10.200 ;
        RECT 2.800 1.600 3.600 9.000 ;
        RECT 6.000 1.600 6.800 6.200 ;
        RECT 9.200 1.600 10.000 6.200 ;
        RECT 12.400 1.600 13.200 6.200 ;
        RECT 15.600 1.600 16.400 6.200 ;
        RECT 23.600 1.600 24.400 6.200 ;
        RECT 26.800 1.600 27.600 6.200 ;
        RECT 33.200 1.600 34.000 6.200 ;
        RECT 36.400 1.600 37.200 6.200 ;
        RECT 39.600 1.600 40.400 6.200 ;
        RECT 41.200 1.600 42.000 10.200 ;
        RECT 62.000 9.600 62.800 10.200 ;
        RECT 65.200 10.000 66.200 10.200 ;
        RECT 49.200 1.600 50.000 9.000 ;
        RECT 58.800 1.600 59.600 6.200 ;
        RECT 62.000 1.600 62.800 6.200 ;
        RECT 65.200 1.600 66.000 6.200 ;
        RECT 71.600 1.600 72.400 6.200 ;
        RECT 74.800 1.600 75.600 6.200 ;
        RECT 82.800 1.600 83.600 6.200 ;
        RECT 86.000 1.600 86.800 6.200 ;
        RECT 89.200 1.600 90.000 6.200 ;
        RECT 92.400 1.600 93.200 6.200 ;
        RECT 95.600 1.600 96.400 9.000 ;
        RECT 98.800 1.600 99.600 10.200 ;
        RECT 102.000 1.600 102.800 10.200 ;
        RECT 105.200 1.600 106.000 10.200 ;
        RECT 108.400 1.600 109.200 9.000 ;
        RECT 111.600 1.600 112.400 6.200 ;
        RECT 114.800 1.600 115.600 10.200 ;
        RECT 148.200 10.000 149.200 10.200 ;
        RECT 151.600 9.600 152.400 10.200 ;
        RECT 159.600 10.200 186.600 10.800 ;
        RECT 215.600 10.200 242.600 10.800 ;
        RECT 159.600 9.600 160.400 10.200 ;
        RECT 162.800 10.000 163.800 10.200 ;
        RECT 119.000 1.600 119.800 6.200 ;
        RECT 121.200 1.600 122.000 6.200 ;
        RECT 124.400 1.600 125.200 6.200 ;
        RECT 127.600 1.600 128.400 6.200 ;
        RECT 130.800 1.600 131.600 6.200 ;
        RECT 138.800 1.600 139.600 6.200 ;
        RECT 142.000 1.600 142.800 6.200 ;
        RECT 148.400 1.600 149.200 6.200 ;
        RECT 151.600 1.600 152.400 6.200 ;
        RECT 154.800 1.600 155.600 6.200 ;
        RECT 156.400 1.600 157.200 6.200 ;
        RECT 159.600 1.600 160.400 6.200 ;
        RECT 162.800 1.600 163.600 6.200 ;
        RECT 169.200 1.600 170.000 6.200 ;
        RECT 172.400 1.600 173.200 6.200 ;
        RECT 180.400 1.600 181.200 6.200 ;
        RECT 183.600 1.600 184.400 6.200 ;
        RECT 186.800 1.600 187.600 6.200 ;
        RECT 190.000 1.600 190.800 6.200 ;
        RECT 198.000 1.600 198.800 6.200 ;
        RECT 201.200 1.600 202.000 10.200 ;
        RECT 206.000 1.600 206.800 6.200 ;
        RECT 209.200 1.600 210.000 9.800 ;
        RECT 215.600 9.600 216.400 10.200 ;
        RECT 218.800 10.000 219.800 10.200 ;
        RECT 212.400 1.600 213.200 6.200 ;
        RECT 215.600 1.600 216.400 6.200 ;
        RECT 218.800 1.600 219.600 6.200 ;
        RECT 225.200 1.600 226.000 6.200 ;
        RECT 228.400 1.600 229.200 6.200 ;
        RECT 236.400 1.600 237.200 6.200 ;
        RECT 239.600 1.600 240.400 6.200 ;
        RECT 242.800 1.600 243.600 6.200 ;
        RECT 246.000 1.600 246.800 6.200 ;
        RECT 247.600 1.600 248.400 10.200 ;
        RECT 251.800 1.600 252.600 6.200 ;
        RECT 0.400 0.400 254.000 1.600 ;
      LAYER via1 ;
        RECT 36.400 163.600 37.200 164.400 ;
        RECT 135.600 170.000 136.400 170.800 ;
        RECT 70.000 165.400 70.800 166.200 ;
        RECT 135.600 163.600 136.400 164.400 ;
        RECT 159.600 165.400 160.400 166.200 ;
        RECT 202.800 163.600 203.600 164.400 ;
        RECT 64.300 160.600 65.100 161.400 ;
        RECT 65.300 160.600 66.100 161.400 ;
        RECT 66.300 160.600 67.100 161.400 ;
        RECT 67.300 160.600 68.100 161.400 ;
        RECT 68.300 160.600 69.100 161.400 ;
        RECT 69.300 160.600 70.100 161.400 ;
        RECT 36.400 157.600 37.200 158.400 ;
        RECT 47.600 157.600 48.400 158.400 ;
        RECT 36.400 151.600 37.200 152.400 ;
        RECT 47.600 151.600 48.400 152.400 ;
        RECT 148.400 151.200 149.200 152.000 ;
        RECT 36.400 123.600 37.200 124.400 ;
        RECT 145.200 130.000 146.000 130.800 ;
        RECT 89.200 125.400 90.000 126.200 ;
        RECT 145.200 125.400 146.000 126.200 ;
        RECT 64.300 120.600 65.100 121.400 ;
        RECT 65.300 120.600 66.100 121.400 ;
        RECT 66.300 120.600 67.100 121.400 ;
        RECT 67.300 120.600 68.100 121.400 ;
        RECT 68.300 120.600 69.100 121.400 ;
        RECT 69.300 120.600 70.100 121.400 ;
        RECT 36.400 117.600 37.200 118.400 ;
        RECT 36.400 111.600 37.200 112.400 ;
        RECT 98.800 117.600 99.600 118.400 ;
        RECT 98.800 111.600 99.600 112.400 ;
        RECT 215.600 111.200 216.400 112.000 ;
        RECT 36.400 83.600 37.200 84.400 ;
        RECT 111.600 83.600 112.400 84.400 ;
        RECT 122.800 83.600 123.600 84.400 ;
        RECT 64.300 80.600 65.100 81.400 ;
        RECT 65.300 80.600 66.100 81.400 ;
        RECT 66.300 80.600 67.100 81.400 ;
        RECT 67.300 80.600 68.100 81.400 ;
        RECT 68.300 80.600 69.100 81.400 ;
        RECT 69.300 80.600 70.100 81.400 ;
        RECT 87.600 77.600 88.400 78.400 ;
        RECT 87.600 71.600 88.400 72.400 ;
        RECT 191.600 71.200 192.400 72.000 ;
        RECT 39.600 43.600 40.400 44.400 ;
        RECT 74.800 43.600 75.600 44.400 ;
        RECT 178.800 50.000 179.600 50.800 ;
        RECT 111.600 45.400 112.400 46.200 ;
        RECT 178.800 45.400 179.600 46.200 ;
        RECT 215.600 45.400 216.400 46.200 ;
        RECT 64.300 40.600 65.100 41.400 ;
        RECT 65.300 40.600 66.100 41.400 ;
        RECT 66.300 40.600 67.100 41.400 ;
        RECT 67.300 40.600 68.100 41.400 ;
        RECT 68.300 40.600 69.100 41.400 ;
        RECT 69.300 40.600 70.100 41.400 ;
        RECT 36.400 37.600 37.200 38.400 ;
        RECT 36.400 31.600 37.200 32.400 ;
        RECT 70.000 31.200 70.800 32.000 ;
        RECT 151.600 37.600 152.400 38.400 ;
        RECT 151.600 31.600 152.400 32.400 ;
        RECT 33.200 10.000 34.000 10.800 ;
        RECT 33.200 3.600 34.000 4.400 ;
        RECT 65.200 5.400 66.000 6.200 ;
        RECT 148.400 10.000 149.200 10.800 ;
        RECT 148.400 3.600 149.200 4.400 ;
        RECT 162.800 3.600 163.600 4.400 ;
        RECT 218.800 3.600 219.600 4.400 ;
        RECT 64.300 0.600 65.100 1.400 ;
        RECT 65.300 0.600 66.100 1.400 ;
        RECT 66.300 0.600 67.100 1.400 ;
        RECT 67.300 0.600 68.100 1.400 ;
        RECT 68.300 0.600 69.100 1.400 ;
        RECT 69.300 0.600 70.100 1.400 ;
      LAYER metal2 ;
        RECT 36.400 169.600 37.200 170.400 ;
        RECT 70.000 170.000 70.800 170.800 ;
        RECT 135.600 170.000 136.400 170.800 ;
        RECT 159.600 170.000 160.400 170.800 ;
        RECT 36.500 164.400 37.100 169.600 ;
        RECT 70.100 166.200 70.700 170.000 ;
        RECT 70.000 165.400 70.800 166.200 ;
        RECT 135.700 164.400 136.300 170.000 ;
        RECT 159.700 166.200 160.300 170.000 ;
        RECT 202.800 169.600 203.600 170.400 ;
        RECT 159.600 165.400 160.400 166.200 ;
        RECT 202.900 164.400 203.500 169.600 ;
        RECT 36.400 163.600 37.200 164.400 ;
        RECT 135.600 163.600 136.400 164.400 ;
        RECT 202.800 163.600 203.600 164.400 ;
        RECT 66.600 161.400 67.800 161.600 ;
        RECT 64.300 160.600 70.100 161.400 ;
        RECT 66.600 160.400 67.800 160.600 ;
        RECT 36.400 157.600 37.200 158.400 ;
        RECT 47.600 157.600 48.400 158.400 ;
        RECT 36.500 152.400 37.100 157.600 ;
        RECT 47.700 152.400 48.300 157.600 ;
        RECT 148.400 155.800 149.200 156.600 ;
        RECT 36.400 151.600 37.200 152.400 ;
        RECT 47.600 151.600 48.400 152.400 ;
        RECT 148.500 152.000 149.100 155.800 ;
        RECT 148.400 151.200 149.200 152.000 ;
        RECT 36.400 129.600 37.200 130.400 ;
        RECT 89.200 130.000 90.000 130.800 ;
        RECT 145.200 130.000 146.000 130.800 ;
        RECT 36.500 124.400 37.100 129.600 ;
        RECT 89.300 126.200 89.900 130.000 ;
        RECT 145.300 126.200 145.900 130.000 ;
        RECT 89.200 125.400 90.000 126.200 ;
        RECT 145.200 125.400 146.000 126.200 ;
        RECT 36.400 123.600 37.200 124.400 ;
        RECT 66.600 121.400 67.800 121.600 ;
        RECT 64.300 120.600 70.100 121.400 ;
        RECT 66.600 120.400 67.800 120.600 ;
        RECT 36.400 117.600 37.200 118.400 ;
        RECT 98.800 117.600 99.600 118.400 ;
        RECT 36.500 112.400 37.100 117.600 ;
        RECT 98.900 112.400 99.500 117.600 ;
        RECT 215.600 115.800 216.400 116.600 ;
        RECT 36.400 111.600 37.200 112.400 ;
        RECT 98.800 111.600 99.600 112.400 ;
        RECT 215.700 112.000 216.300 115.800 ;
        RECT 215.600 111.200 216.400 112.000 ;
        RECT 36.400 89.600 37.200 90.400 ;
        RECT 111.600 89.600 112.400 90.400 ;
        RECT 122.800 90.000 123.600 90.800 ;
        RECT 36.500 84.400 37.100 89.600 ;
        RECT 111.700 84.400 112.300 89.600 ;
        RECT 122.900 84.400 123.500 90.000 ;
        RECT 36.400 83.600 37.200 84.400 ;
        RECT 111.600 83.600 112.400 84.400 ;
        RECT 122.800 83.600 123.600 84.400 ;
        RECT 66.600 81.400 67.800 81.600 ;
        RECT 64.300 80.600 70.100 81.400 ;
        RECT 66.600 80.400 67.800 80.600 ;
        RECT 87.600 77.600 88.400 78.400 ;
        RECT 87.700 72.400 88.300 77.600 ;
        RECT 191.600 75.800 192.400 76.600 ;
        RECT 87.600 71.600 88.400 72.400 ;
        RECT 191.700 72.000 192.300 75.800 ;
        RECT 191.600 71.200 192.400 72.000 ;
        RECT 39.600 49.600 40.400 50.400 ;
        RECT 74.800 49.600 75.600 50.400 ;
        RECT 111.600 50.000 112.400 50.800 ;
        RECT 178.800 50.000 179.600 50.800 ;
        RECT 215.600 50.000 216.400 50.800 ;
        RECT 39.700 44.400 40.300 49.600 ;
        RECT 74.900 44.400 75.500 49.600 ;
        RECT 111.700 46.200 112.300 50.000 ;
        RECT 178.900 46.200 179.500 50.000 ;
        RECT 215.700 46.200 216.300 50.000 ;
        RECT 111.600 45.400 112.400 46.200 ;
        RECT 178.800 45.400 179.600 46.200 ;
        RECT 215.600 45.400 216.400 46.200 ;
        RECT 39.600 43.600 40.400 44.400 ;
        RECT 74.800 43.600 75.600 44.400 ;
        RECT 66.600 41.400 67.800 41.600 ;
        RECT 64.300 40.600 70.100 41.400 ;
        RECT 66.600 40.400 67.800 40.600 ;
        RECT 36.400 37.600 37.200 38.400 ;
        RECT 151.600 37.600 152.400 38.400 ;
        RECT 36.500 32.400 37.100 37.600 ;
        RECT 70.000 35.800 70.800 36.600 ;
        RECT 36.400 31.600 37.200 32.400 ;
        RECT 70.100 32.000 70.700 35.800 ;
        RECT 151.700 32.400 152.300 37.600 ;
        RECT 220.400 35.600 221.200 36.400 ;
        RECT 70.000 31.200 70.800 32.000 ;
        RECT 151.600 31.600 152.400 32.400 ;
        RECT 220.500 30.400 221.100 35.600 ;
        RECT 220.400 29.600 221.200 30.400 ;
        RECT 33.200 10.000 34.000 10.800 ;
        RECT 65.200 10.000 66.000 10.800 ;
        RECT 148.400 10.000 149.200 10.800 ;
        RECT 162.800 10.000 163.600 10.800 ;
        RECT 218.800 10.000 219.600 10.800 ;
        RECT 33.300 4.400 33.900 10.000 ;
        RECT 65.300 6.200 65.900 10.000 ;
        RECT 65.200 5.400 66.000 6.200 ;
        RECT 148.500 4.400 149.100 10.000 ;
        RECT 162.900 4.400 163.500 10.000 ;
        RECT 218.900 4.400 219.500 10.000 ;
        RECT 33.200 3.600 34.000 4.400 ;
        RECT 148.400 3.600 149.200 4.400 ;
        RECT 162.800 3.600 163.600 4.400 ;
        RECT 218.800 3.600 219.600 4.400 ;
        RECT 66.600 1.400 67.800 1.600 ;
        RECT 64.300 0.600 70.100 1.400 ;
        RECT 66.600 0.400 67.800 0.600 ;
      LAYER via2 ;
        RECT 65.300 160.600 66.100 161.400 ;
        RECT 66.300 160.600 67.100 161.400 ;
        RECT 67.300 160.600 68.100 161.400 ;
        RECT 68.300 160.600 69.100 161.400 ;
        RECT 69.300 160.600 70.100 161.400 ;
        RECT 65.300 120.600 66.100 121.400 ;
        RECT 66.300 120.600 67.100 121.400 ;
        RECT 67.300 120.600 68.100 121.400 ;
        RECT 68.300 120.600 69.100 121.400 ;
        RECT 69.300 120.600 70.100 121.400 ;
        RECT 65.300 80.600 66.100 81.400 ;
        RECT 66.300 80.600 67.100 81.400 ;
        RECT 67.300 80.600 68.100 81.400 ;
        RECT 68.300 80.600 69.100 81.400 ;
        RECT 69.300 80.600 70.100 81.400 ;
        RECT 65.300 40.600 66.100 41.400 ;
        RECT 66.300 40.600 67.100 41.400 ;
        RECT 67.300 40.600 68.100 41.400 ;
        RECT 68.300 40.600 69.100 41.400 ;
        RECT 69.300 40.600 70.100 41.400 ;
        RECT 65.300 0.600 66.100 1.400 ;
        RECT 66.300 0.600 67.100 1.400 ;
        RECT 67.300 0.600 68.100 1.400 ;
        RECT 68.300 0.600 69.100 1.400 ;
        RECT 69.300 0.600 70.100 1.400 ;
      LAYER metal3 ;
        RECT 64.200 160.400 70.200 161.600 ;
        RECT 64.200 120.400 70.200 121.600 ;
        RECT 64.200 80.400 70.200 81.600 ;
        RECT 64.200 40.400 70.200 41.600 ;
        RECT 64.200 0.400 70.200 1.600 ;
      LAYER via3 ;
        RECT 64.400 160.600 65.200 161.400 ;
        RECT 65.600 160.600 66.400 161.400 ;
        RECT 66.800 160.600 67.600 161.400 ;
        RECT 68.000 160.600 68.800 161.400 ;
        RECT 69.200 160.600 70.000 161.400 ;
        RECT 64.400 120.600 65.200 121.400 ;
        RECT 65.600 120.600 66.400 121.400 ;
        RECT 66.800 120.600 67.600 121.400 ;
        RECT 68.000 120.600 68.800 121.400 ;
        RECT 69.200 120.600 70.000 121.400 ;
        RECT 64.400 80.600 65.200 81.400 ;
        RECT 65.600 80.600 66.400 81.400 ;
        RECT 66.800 80.600 67.600 81.400 ;
        RECT 68.000 80.600 68.800 81.400 ;
        RECT 69.200 80.600 70.000 81.400 ;
        RECT 64.400 40.600 65.200 41.400 ;
        RECT 65.600 40.600 66.400 41.400 ;
        RECT 66.800 40.600 67.600 41.400 ;
        RECT 68.000 40.600 68.800 41.400 ;
        RECT 69.200 40.600 70.000 41.400 ;
        RECT 64.400 0.600 65.200 1.400 ;
        RECT 65.600 0.600 66.400 1.400 ;
        RECT 66.800 0.600 67.600 1.400 ;
        RECT 68.000 0.600 68.800 1.400 ;
        RECT 69.200 0.600 70.000 1.400 ;
      LAYER metal4 ;
        RECT 64.000 -1.000 70.400 181.600 ;
    END
  END vdd
  PIN N[8]
    PORT
      LAYER metal1 ;
        RECT 244.400 24.800 245.200 26.400 ;
        RECT 252.400 10.300 253.200 10.400 ;
        RECT 254.000 10.300 254.800 10.400 ;
        RECT 252.400 10.200 254.800 10.300 ;
        RECT 251.800 9.700 254.800 10.200 ;
        RECT 251.800 9.600 253.200 9.700 ;
        RECT 254.000 9.600 254.800 9.700 ;
        RECT 251.800 8.400 252.400 9.600 ;
        RECT 251.600 7.600 252.400 8.400 ;
      LAYER via1 ;
        RECT 244.400 25.600 245.200 26.400 ;
      LAYER metal2 ;
        RECT 244.400 25.600 245.200 26.400 ;
        RECT 254.000 25.600 254.800 26.400 ;
        RECT 254.100 10.400 254.700 25.600 ;
        RECT 254.000 9.600 254.800 10.400 ;
      LAYER metal3 ;
        RECT 244.400 26.300 245.200 26.400 ;
        RECT 254.000 26.300 254.800 26.400 ;
        RECT 244.400 25.700 254.800 26.300 ;
        RECT 244.400 25.600 245.200 25.700 ;
        RECT 254.000 25.600 254.800 25.700 ;
        RECT 254.000 10.300 254.800 10.400 ;
        RECT 254.000 9.700 257.900 10.300 ;
        RECT 254.000 9.600 254.800 9.700 ;
    END
  END N[8]
  PIN N[7]
    PORT
      LAYER metal1 ;
        RECT 240.400 67.600 242.000 68.400 ;
        RECT 252.400 64.800 253.200 66.400 ;
        RECT 248.400 14.400 249.200 14.800 ;
        RECT 247.600 13.800 249.200 14.400 ;
        RECT 247.600 13.600 248.400 13.800 ;
      LAYER via1 ;
        RECT 241.200 67.600 242.000 68.400 ;
        RECT 252.400 65.600 253.200 66.400 ;
      LAYER metal2 ;
        RECT 241.200 67.600 242.000 68.400 ;
        RECT 241.300 66.400 241.900 67.600 ;
        RECT 241.200 65.600 242.000 66.400 ;
        RECT 252.400 65.600 253.200 66.400 ;
        RECT 247.600 13.600 248.400 14.400 ;
      LAYER metal3 ;
        RECT 241.200 66.300 242.000 66.400 ;
        RECT 247.600 66.300 248.400 66.400 ;
        RECT 252.400 66.300 253.200 66.400 ;
        RECT 241.200 65.700 257.900 66.300 ;
        RECT 241.200 65.600 242.000 65.700 ;
        RECT 247.600 65.600 248.400 65.700 ;
        RECT 252.400 65.600 253.200 65.700 ;
        RECT 247.600 13.600 248.400 14.400 ;
      LAYER metal4 ;
        RECT 247.400 13.400 248.600 66.600 ;
    END
  END N[7]
  PIN N[6]
    PORT
      LAYER metal1 ;
        RECT 242.000 153.600 242.800 154.400 ;
        RECT 242.200 152.400 242.800 153.600 ;
        RECT 242.200 151.800 243.600 152.400 ;
        RECT 242.800 151.600 243.600 151.800 ;
        RECT 250.800 149.600 251.600 151.200 ;
      LAYER metal2 ;
        RECT 250.800 159.600 251.600 160.400 ;
        RECT 242.800 151.600 243.600 152.400 ;
        RECT 242.900 150.400 243.500 151.600 ;
        RECT 250.900 150.400 251.500 159.600 ;
        RECT 242.800 149.600 243.600 150.400 ;
        RECT 250.800 149.600 251.600 150.400 ;
      LAYER metal3 ;
        RECT 250.800 160.300 251.600 160.400 ;
        RECT 250.800 159.700 257.900 160.300 ;
        RECT 250.800 159.600 251.600 159.700 ;
        RECT 242.800 150.300 243.600 150.400 ;
        RECT 250.800 150.300 251.600 150.400 ;
        RECT 242.800 149.700 251.600 150.300 ;
        RECT 242.800 149.600 243.600 149.700 ;
        RECT 250.800 149.600 251.600 149.700 ;
    END
  END N[6]
  PIN N[5]
    PORT
      LAYER metal1 ;
        RECT 229.200 147.600 230.800 148.400 ;
        RECT 238.000 148.200 238.800 148.400 ;
        RECT 238.000 147.600 239.600 148.200 ;
        RECT 238.800 147.200 239.600 147.600 ;
        RECT 247.600 144.800 248.400 146.400 ;
      LAYER via1 ;
        RECT 230.000 147.600 230.800 148.400 ;
        RECT 247.600 145.600 248.400 146.400 ;
      LAYER metal2 ;
        RECT 230.000 147.600 230.800 148.400 ;
        RECT 238.000 147.600 238.800 148.400 ;
        RECT 230.100 146.400 230.700 147.600 ;
        RECT 238.100 146.400 238.700 147.600 ;
        RECT 230.000 145.600 230.800 146.400 ;
        RECT 238.000 145.600 238.800 146.400 ;
        RECT 247.600 145.600 248.400 146.400 ;
      LAYER metal3 ;
        RECT 247.700 147.700 257.900 148.300 ;
        RECT 247.700 146.400 248.300 147.700 ;
        RECT 230.000 146.300 230.800 146.400 ;
        RECT 238.000 146.300 238.800 146.400 ;
        RECT 247.600 146.300 248.400 146.400 ;
        RECT 230.000 145.700 248.400 146.300 ;
        RECT 230.000 145.600 230.800 145.700 ;
        RECT 238.000 145.600 238.800 145.700 ;
        RECT 247.600 145.600 248.400 145.700 ;
    END
  END N[5]
  PIN N[4]
    PORT
      LAYER metal1 ;
        RECT 242.800 172.300 243.600 172.400 ;
        RECT 244.400 172.300 245.200 172.400 ;
        RECT 242.800 171.700 245.200 172.300 ;
        RECT 242.800 170.800 243.600 171.700 ;
        RECT 244.400 171.600 245.200 171.700 ;
        RECT 248.400 114.300 249.200 114.400 ;
        RECT 254.000 114.300 254.800 114.400 ;
        RECT 248.400 113.700 254.800 114.300 ;
        RECT 248.400 113.600 249.200 113.700 ;
        RECT 254.000 113.600 254.800 113.700 ;
        RECT 248.600 112.400 249.200 113.600 ;
        RECT 248.600 111.800 250.000 112.400 ;
        RECT 249.200 111.600 250.000 111.800 ;
      LAYER metal2 ;
        RECT 244.400 172.300 245.200 172.400 ;
        RECT 244.400 171.700 246.700 172.300 ;
        RECT 244.400 171.600 245.200 171.700 ;
        RECT 246.100 152.400 246.700 171.700 ;
        RECT 246.000 151.600 246.800 152.400 ;
        RECT 254.000 151.600 254.800 152.400 ;
        RECT 254.100 114.400 254.700 151.600 ;
        RECT 254.000 113.600 254.800 114.400 ;
      LAYER metal3 ;
        RECT 246.000 152.300 246.800 152.400 ;
        RECT 254.000 152.300 254.800 152.400 ;
        RECT 246.000 151.700 257.900 152.300 ;
        RECT 246.000 151.600 246.800 151.700 ;
        RECT 254.000 151.600 254.800 151.700 ;
    END
  END N[4]
  PIN N[3]
    PORT
      LAYER metal1 ;
        RECT 239.600 175.600 240.400 177.200 ;
        RECT 244.400 108.200 245.200 108.400 ;
        RECT 244.400 107.600 246.000 108.200 ;
        RECT 245.200 107.200 246.000 107.600 ;
        RECT 243.600 94.400 244.400 94.800 ;
        RECT 243.600 93.800 245.200 94.400 ;
        RECT 244.400 93.600 245.200 93.800 ;
        RECT 250.800 92.200 251.600 92.400 ;
        RECT 250.000 91.600 251.600 92.200 ;
        RECT 250.000 91.200 250.800 91.600 ;
      LAYER via1 ;
        RECT 250.800 91.600 251.600 92.400 ;
      LAYER metal2 ;
        RECT 239.600 175.600 240.400 176.400 ;
        RECT 244.400 127.600 245.200 128.400 ;
        RECT 244.500 108.400 245.100 127.600 ;
        RECT 244.400 107.600 245.200 108.400 ;
        RECT 244.500 94.400 245.100 107.600 ;
        RECT 244.400 93.600 245.200 94.400 ;
        RECT 244.500 92.400 245.100 93.600 ;
        RECT 244.400 91.600 245.200 92.400 ;
        RECT 250.800 91.600 251.600 92.400 ;
      LAYER metal3 ;
        RECT 239.600 176.300 240.400 176.400 ;
        RECT 244.400 176.300 245.200 176.400 ;
        RECT 239.600 175.700 245.200 176.300 ;
        RECT 239.600 175.600 240.400 175.700 ;
        RECT 244.400 175.600 245.200 175.700 ;
        RECT 244.400 127.600 245.200 128.400 ;
        RECT 244.400 92.300 245.200 92.400 ;
        RECT 250.800 92.300 251.600 92.400 ;
        RECT 244.400 91.700 257.900 92.300 ;
        RECT 244.400 91.600 245.200 91.700 ;
        RECT 250.800 91.600 251.600 91.700 ;
      LAYER metal4 ;
        RECT 244.200 127.400 245.400 176.600 ;
    END
  END N[3]
  PIN N[2]
    PORT
      LAYER metal1 ;
        RECT 244.400 168.800 245.200 170.400 ;
        RECT 238.000 135.600 238.800 137.200 ;
      LAYER via1 ;
        RECT 244.400 169.600 245.200 170.400 ;
      LAYER metal2 ;
        RECT 244.400 169.600 245.200 170.400 ;
        RECT 244.500 156.400 245.100 169.600 ;
        RECT 244.400 155.600 245.200 156.400 ;
        RECT 238.000 143.600 238.800 144.400 ;
        RECT 238.100 136.400 238.700 143.600 ;
        RECT 238.000 135.600 238.800 136.400 ;
      LAYER metal3 ;
        RECT 244.400 156.300 245.200 156.400 ;
        RECT 247.600 156.300 248.400 156.400 ;
        RECT 244.400 155.700 257.900 156.300 ;
        RECT 244.400 155.600 245.200 155.700 ;
        RECT 247.600 155.600 248.400 155.700 ;
        RECT 238.000 144.300 238.800 144.400 ;
        RECT 247.600 144.300 248.400 144.400 ;
        RECT 238.000 143.700 248.400 144.300 ;
        RECT 238.000 143.600 238.800 143.700 ;
        RECT 247.600 143.600 248.400 143.700 ;
      LAYER metal4 ;
        RECT 247.400 143.400 248.600 156.600 ;
    END
  END N[2]
  PIN N[1]
    PORT
      LAYER metal1 ;
        RECT 247.600 173.600 248.400 175.200 ;
        RECT 223.600 135.600 224.400 137.200 ;
        RECT 210.800 131.600 211.600 133.200 ;
      LAYER metal2 ;
        RECT 247.600 173.600 248.400 174.400 ;
        RECT 210.800 137.600 211.600 138.400 ;
        RECT 223.600 137.600 224.400 138.400 ;
        RECT 210.900 132.400 211.500 137.600 ;
        RECT 223.700 136.400 224.300 137.600 ;
        RECT 223.600 135.600 224.400 136.400 ;
        RECT 210.800 131.600 211.600 132.400 ;
      LAYER metal3 ;
        RECT 228.400 174.300 229.200 174.400 ;
        RECT 247.600 174.300 248.400 174.400 ;
        RECT 228.400 173.700 257.900 174.300 ;
        RECT 228.400 173.600 229.200 173.700 ;
        RECT 247.600 173.600 248.400 173.700 ;
        RECT 210.800 138.300 211.600 138.400 ;
        RECT 223.600 138.300 224.400 138.400 ;
        RECT 228.400 138.300 229.200 138.400 ;
        RECT 210.800 137.700 229.200 138.300 ;
        RECT 210.800 137.600 211.600 137.700 ;
        RECT 223.600 137.600 224.400 137.700 ;
        RECT 228.400 137.600 229.200 137.700 ;
      LAYER metal4 ;
        RECT 228.200 137.400 229.400 174.600 ;
    END
  END N[1]
  PIN N[0]
    PORT
      LAYER metal1 ;
        RECT 127.600 26.800 128.400 28.400 ;
      LAYER via1 ;
        RECT 127.600 27.600 128.400 28.400 ;
      LAYER metal2 ;
        RECT 127.600 27.600 128.400 28.400 ;
        RECT 127.700 -1.700 128.300 27.600 ;
        RECT 126.100 -2.300 128.300 -1.700 ;
    END
  END N[0]
  PIN clock
    PORT
      LAYER metal1 ;
        RECT 6.000 68.200 7.800 69.000 ;
        RECT 20.400 68.200 22.200 69.000 ;
        RECT 65.200 68.200 67.000 69.000 ;
        RECT 6.000 67.600 6.800 68.200 ;
        RECT 20.400 67.600 21.200 68.200 ;
        RECT 65.200 67.600 66.000 68.200 ;
        RECT 110.000 28.200 111.800 29.000 ;
        RECT 129.200 28.200 131.000 29.000 ;
        RECT 110.000 27.600 110.800 28.200 ;
        RECT 129.200 27.600 130.000 28.200 ;
      LAYER metal2 ;
        RECT 6.000 67.600 6.800 68.400 ;
        RECT 20.400 67.600 21.200 68.400 ;
        RECT 65.200 67.600 66.000 68.400 ;
        RECT 65.300 66.400 65.900 67.600 ;
        RECT 65.200 65.600 66.000 66.400 ;
        RECT 65.300 56.400 65.900 65.600 ;
        RECT 65.200 55.600 66.000 56.400 ;
        RECT 110.000 55.600 110.800 56.400 ;
        RECT 110.100 28.400 110.700 55.600 ;
        RECT 110.000 27.600 110.800 28.400 ;
        RECT 129.200 27.600 130.000 28.400 ;
      LAYER metal3 ;
        RECT 6.000 68.300 6.800 68.400 ;
        RECT 20.400 68.300 21.200 68.400 ;
        RECT -3.500 67.700 21.200 68.300 ;
        RECT 6.000 67.600 6.800 67.700 ;
        RECT 20.400 67.600 21.200 67.700 ;
        RECT 20.500 66.300 21.100 67.600 ;
        RECT 65.200 66.300 66.000 66.400 ;
        RECT 20.500 65.700 66.000 66.300 ;
        RECT 65.200 65.600 66.000 65.700 ;
        RECT 65.200 56.300 66.000 56.400 ;
        RECT 110.000 56.300 110.800 56.400 ;
        RECT 65.200 55.700 110.800 56.300 ;
        RECT 65.200 55.600 66.000 55.700 ;
        RECT 110.000 55.600 110.800 55.700 ;
        RECT 110.000 28.300 110.800 28.400 ;
        RECT 129.200 28.300 130.000 28.400 ;
        RECT 110.000 27.700 130.000 28.300 ;
        RECT 110.000 27.600 110.800 27.700 ;
        RECT 129.200 27.600 130.000 27.700 ;
    END
  END clock
  PIN counter[7]
    PORT
      LAYER metal1 ;
        RECT 247.600 52.400 248.400 59.800 ;
        RECT 247.800 50.200 248.400 52.400 ;
        RECT 247.600 42.200 248.400 50.200 ;
      LAYER via1 ;
        RECT 247.600 47.600 248.400 48.400 ;
      LAYER metal2 ;
        RECT 247.600 49.600 248.400 50.400 ;
        RECT 247.700 48.400 248.300 49.600 ;
        RECT 247.600 47.600 248.400 48.400 ;
      LAYER metal3 ;
        RECT 247.600 50.300 248.400 50.400 ;
        RECT 247.600 49.700 257.900 50.300 ;
        RECT 247.600 49.600 248.400 49.700 ;
    END
  END counter[7]
  PIN counter[6]
    PORT
      LAYER metal1 ;
        RECT 190.000 31.800 190.800 39.800 ;
        RECT 190.000 29.600 190.600 31.800 ;
        RECT 190.000 22.200 190.800 29.600 ;
      LAYER via1 ;
        RECT 190.000 23.600 190.800 24.400 ;
      LAYER metal2 ;
        RECT 190.000 23.600 190.800 24.400 ;
        RECT 193.200 23.600 194.000 24.400 ;
        RECT 193.300 -2.300 193.900 23.600 ;
      LAYER metal3 ;
        RECT 190.000 24.300 190.800 24.400 ;
        RECT 193.200 24.300 194.000 24.400 ;
        RECT 190.000 23.700 194.000 24.300 ;
        RECT 190.000 23.600 190.800 23.700 ;
        RECT 193.200 23.600 194.000 23.700 ;
    END
  END counter[6]
  PIN counter[5]
    PORT
      LAYER metal1 ;
        RECT 151.600 172.400 152.400 179.800 ;
        RECT 151.800 170.200 152.400 172.400 ;
        RECT 151.600 162.200 152.400 170.200 ;
      LAYER via1 ;
        RECT 151.600 177.600 152.400 178.400 ;
      LAYER metal2 ;
        RECT 150.100 185.700 152.300 186.300 ;
        RECT 151.700 178.400 152.300 185.700 ;
        RECT 151.600 177.600 152.400 178.400 ;
    END
  END counter[5]
  PIN counter[4]
    PORT
      LAYER metal1 ;
        RECT 177.200 151.800 178.000 159.800 ;
        RECT 177.200 149.600 177.800 151.800 ;
        RECT 177.200 142.200 178.000 149.600 ;
      LAYER via1 ;
        RECT 177.200 157.600 178.000 158.400 ;
      LAYER metal2 ;
        RECT 177.300 185.700 179.500 186.300 ;
        RECT 177.300 158.400 177.900 185.700 ;
        RECT 177.200 157.600 178.000 158.400 ;
    END
  END counter[4]
  PIN counter[3]
    PORT
      LAYER metal1 ;
        RECT 249.200 31.800 250.000 39.800 ;
        RECT 249.400 29.600 250.000 31.800 ;
        RECT 249.200 28.300 250.000 29.600 ;
        RECT 254.000 28.300 254.800 28.400 ;
        RECT 249.200 27.700 254.800 28.300 ;
        RECT 249.200 22.200 250.000 27.700 ;
        RECT 254.000 27.600 254.800 27.700 ;
      LAYER metal2 ;
        RECT 254.000 29.600 254.800 30.400 ;
        RECT 254.100 28.400 254.700 29.600 ;
        RECT 254.000 27.600 254.800 28.400 ;
      LAYER metal3 ;
        RECT 254.000 30.300 254.800 30.400 ;
        RECT 254.000 29.700 257.900 30.300 ;
        RECT 254.000 29.600 254.800 29.700 ;
    END
  END counter[3]
  PIN counter[2]
    PORT
      LAYER metal1 ;
        RECT 252.400 172.400 253.200 179.800 ;
        RECT 252.600 170.200 253.200 172.400 ;
        RECT 252.400 168.300 253.200 170.200 ;
        RECT 254.000 168.300 254.800 168.400 ;
        RECT 252.400 167.700 254.800 168.300 ;
        RECT 252.400 162.200 253.200 167.700 ;
        RECT 254.000 167.600 254.800 167.700 ;
      LAYER metal2 ;
        RECT 254.000 169.600 254.800 170.400 ;
        RECT 254.100 168.400 254.700 169.600 ;
        RECT 254.000 167.600 254.800 168.400 ;
      LAYER metal3 ;
        RECT 254.000 170.300 254.800 170.400 ;
        RECT 254.000 169.700 257.900 170.300 ;
        RECT 254.000 169.600 254.800 169.700 ;
    END
  END counter[2]
  PIN counter[1]
    PORT
      LAYER metal1 ;
        RECT 198.000 172.400 198.800 179.800 ;
        RECT 198.200 170.200 198.800 172.400 ;
        RECT 198.000 162.200 198.800 170.200 ;
      LAYER via1 ;
        RECT 198.000 177.600 198.800 178.400 ;
      LAYER metal2 ;
        RECT 196.500 185.700 198.700 186.300 ;
        RECT 198.100 178.400 198.700 185.700 ;
        RECT 198.000 177.600 198.800 178.400 ;
    END
  END counter[1]
  PIN counter[0]
    PORT
      LAYER metal1 ;
        RECT 238.000 172.400 238.800 179.800 ;
        RECT 238.200 170.200 238.800 172.400 ;
        RECT 238.000 162.200 238.800 170.200 ;
      LAYER via1 ;
        RECT 238.000 177.600 238.800 178.400 ;
      LAYER metal2 ;
        RECT 236.500 185.700 238.700 186.300 ;
        RECT 238.100 178.400 238.700 185.700 ;
        RECT 238.000 177.600 238.800 178.400 ;
    END
  END counter[0]
  PIN done
    PORT
      LAYER metal1 ;
        RECT 135.600 151.800 136.400 159.800 ;
        RECT 135.800 149.600 136.400 151.800 ;
        RECT 135.600 142.200 136.400 149.600 ;
      LAYER via1 ;
        RECT 135.600 157.600 136.400 158.400 ;
      LAYER metal2 ;
        RECT 134.100 182.400 134.700 186.300 ;
        RECT 134.000 181.600 134.800 182.400 ;
        RECT 135.600 161.600 136.400 162.400 ;
        RECT 135.700 158.400 136.300 161.600 ;
        RECT 135.600 157.600 136.400 158.400 ;
      LAYER metal3 ;
        RECT 134.000 182.300 134.800 182.400 ;
        RECT 135.600 182.300 136.400 182.400 ;
        RECT 134.000 181.700 136.400 182.300 ;
        RECT 134.000 181.600 134.800 181.700 ;
        RECT 135.600 181.600 136.400 181.700 ;
        RECT 135.600 161.600 136.400 162.400 ;
      LAYER metal4 ;
        RECT 135.400 161.400 136.600 182.600 ;
    END
  END done
  PIN dp[8]
    PORT
      LAYER metal1 ;
        RECT 1.200 172.400 2.000 179.800 ;
        RECT 1.200 170.200 1.800 172.400 ;
        RECT 1.200 162.200 2.000 170.200 ;
      LAYER via1 ;
        RECT 1.200 167.600 2.000 168.400 ;
      LAYER metal2 ;
        RECT 1.200 169.600 2.000 170.400 ;
        RECT 1.300 168.400 1.900 169.600 ;
        RECT 1.200 167.600 2.000 168.400 ;
      LAYER metal3 ;
        RECT 1.200 170.300 2.000 170.400 ;
        RECT -3.500 169.700 2.000 170.300 ;
        RECT 1.200 169.600 2.000 169.700 ;
    END
  END dp[8]
  PIN dp[7]
    PORT
      LAYER metal1 ;
        RECT 103.600 172.400 104.400 179.800 ;
        RECT 103.600 170.200 104.200 172.400 ;
        RECT 103.600 162.200 104.400 170.200 ;
      LAYER via1 ;
        RECT 103.600 177.600 104.400 178.400 ;
      LAYER metal2 ;
        RECT 103.700 185.700 105.900 186.300 ;
        RECT 103.700 178.400 104.300 185.700 ;
        RECT 103.600 177.600 104.400 178.400 ;
    END
  END dp[7]
  PIN dp[6]
    PORT
      LAYER metal1 ;
        RECT 97.200 12.400 98.000 19.800 ;
        RECT 97.400 10.200 98.000 12.400 ;
        RECT 97.200 2.200 98.000 10.200 ;
      LAYER via1 ;
        RECT 97.200 3.600 98.000 4.400 ;
      LAYER metal2 ;
        RECT 97.200 3.600 98.000 4.400 ;
        RECT 97.300 -1.700 97.900 3.600 ;
        RECT 95.700 -2.300 97.900 -1.700 ;
    END
  END dp[6]
  PIN dp[5]
    PORT
      LAYER metal1 ;
        RECT 102.000 172.400 102.800 179.800 ;
        RECT 102.200 170.200 102.800 172.400 ;
        RECT 102.000 162.200 102.800 170.200 ;
      LAYER via1 ;
        RECT 102.000 177.600 102.800 178.400 ;
      LAYER metal2 ;
        RECT 100.500 185.700 102.700 186.300 ;
        RECT 102.100 178.400 102.700 185.700 ;
        RECT 102.000 177.600 102.800 178.400 ;
    END
  END dp[5]
  PIN dp[4]
    PORT
      LAYER metal1 ;
        RECT 1.200 111.800 2.000 119.800 ;
        RECT 1.200 109.600 1.800 111.800 ;
        RECT 1.200 102.200 2.000 109.600 ;
      LAYER via1 ;
        RECT 1.200 107.600 2.000 108.400 ;
      LAYER metal2 ;
        RECT 1.200 109.600 2.000 110.400 ;
        RECT 1.300 108.400 1.900 109.600 ;
        RECT 1.200 107.600 2.000 108.400 ;
      LAYER metal3 ;
        RECT 1.200 110.300 2.000 110.400 ;
        RECT -3.500 109.700 2.000 110.300 ;
        RECT 1.200 109.600 2.000 109.700 ;
    END
  END dp[4]
  PIN dp[3]
    PORT
      LAYER metal1 ;
        RECT 1.200 31.800 2.000 39.800 ;
        RECT 1.200 29.600 1.800 31.800 ;
        RECT 1.200 22.200 2.000 29.600 ;
      LAYER via1 ;
        RECT 1.200 27.600 2.000 28.400 ;
      LAYER metal2 ;
        RECT 1.200 29.600 2.000 30.400 ;
        RECT 1.300 28.400 1.900 29.600 ;
        RECT 1.200 27.600 2.000 28.400 ;
      LAYER metal3 ;
        RECT 1.200 30.300 2.000 30.400 ;
        RECT -3.500 29.700 2.000 30.300 ;
        RECT 1.200 29.600 2.000 29.700 ;
    END
  END dp[3]
  PIN dp[2]
    PORT
      LAYER metal1 ;
        RECT 1.200 12.400 2.000 19.800 ;
        RECT 1.200 10.200 1.800 12.400 ;
        RECT 1.200 2.200 2.000 10.200 ;
      LAYER via1 ;
        RECT 1.200 7.600 2.000 8.400 ;
      LAYER metal2 ;
        RECT 1.200 9.600 2.000 10.400 ;
        RECT 1.300 8.400 1.900 9.600 ;
        RECT 1.200 7.600 2.000 8.400 ;
      LAYER metal3 ;
        RECT 1.200 10.300 2.000 10.400 ;
        RECT -3.500 9.700 2.000 10.300 ;
        RECT 1.200 9.600 2.000 9.700 ;
    END
  END dp[2]
  PIN dp[1]
    PORT
      LAYER metal1 ;
        RECT 116.400 151.800 117.200 159.800 ;
        RECT 116.600 149.600 117.200 151.800 ;
        RECT 116.400 142.200 117.200 149.600 ;
      LAYER via1 ;
        RECT 116.400 157.600 117.200 158.400 ;
      LAYER metal2 ;
        RECT 114.900 185.700 117.100 186.300 ;
        RECT 116.500 158.400 117.100 185.700 ;
        RECT 116.400 157.600 117.200 158.400 ;
    END
  END dp[1]
  PIN dp[0]
    PORT
      LAYER metal1 ;
        RECT 106.800 12.400 107.600 19.800 ;
        RECT 106.800 10.200 107.400 12.400 ;
        RECT 106.800 2.200 107.600 10.200 ;
      LAYER via1 ;
        RECT 106.800 3.600 107.600 4.400 ;
      LAYER metal2 ;
        RECT 106.800 3.600 107.600 4.400 ;
        RECT 106.900 -2.300 107.500 3.600 ;
    END
  END dp[0]
  PIN reset
    PORT
      LAYER metal1 ;
        RECT 105.200 13.600 106.000 15.200 ;
      LAYER metal2 ;
        RECT 105.200 13.600 106.000 14.400 ;
        RECT 105.300 2.400 105.900 13.600 ;
        RECT 105.200 1.600 106.000 2.400 ;
        RECT 110.000 1.600 110.800 2.400 ;
        RECT 110.100 -2.300 110.700 1.600 ;
      LAYER metal3 ;
        RECT 105.200 2.300 106.000 2.400 ;
        RECT 110.000 2.300 110.800 2.400 ;
        RECT 105.200 1.700 110.800 2.300 ;
        RECT 105.200 1.600 106.000 1.700 ;
        RECT 110.000 1.600 110.800 1.700 ;
    END
  END reset
  PIN sr[7]
    PORT
      LAYER metal1 ;
        RECT 52.400 172.400 53.200 179.800 ;
        RECT 52.400 170.200 53.000 172.400 ;
        RECT 52.400 162.200 53.200 170.200 ;
      LAYER via1 ;
        RECT 52.400 177.600 53.200 178.400 ;
      LAYER metal2 ;
        RECT 52.500 185.700 54.700 186.300 ;
        RECT 52.500 178.400 53.100 185.700 ;
        RECT 52.400 177.600 53.200 178.400 ;
    END
  END sr[7]
  PIN sr[6]
    PORT
      LAYER metal1 ;
        RECT 146.800 172.400 147.600 179.800 ;
        RECT 147.000 170.200 147.600 172.400 ;
        RECT 146.800 162.200 147.600 170.200 ;
      LAYER via1 ;
        RECT 146.800 177.600 147.600 178.400 ;
      LAYER metal2 ;
        RECT 145.300 185.700 147.500 186.300 ;
        RECT 146.900 178.400 147.500 185.700 ;
        RECT 146.800 177.600 147.600 178.400 ;
    END
  END sr[6]
  PIN sr[5]
    PORT
      LAYER metal1 ;
        RECT 65.200 114.300 66.000 114.400 ;
        RECT 71.600 114.300 72.400 119.800 ;
        RECT 65.200 113.700 72.400 114.300 ;
        RECT 65.200 113.600 66.000 113.700 ;
        RECT 71.600 111.800 72.400 113.700 ;
        RECT 71.600 109.600 72.200 111.800 ;
        RECT 71.600 102.200 72.400 109.600 ;
      LAYER metal2 ;
        RECT 65.200 113.600 66.000 114.400 ;
      LAYER metal3 ;
        RECT 65.200 114.300 66.000 114.400 ;
        RECT -3.500 113.700 66.000 114.300 ;
        RECT 65.200 113.600 66.000 113.700 ;
    END
  END sr[5]
  PIN sr[4]
    PORT
      LAYER metal1 ;
        RECT 1.200 92.400 2.000 99.800 ;
        RECT 1.200 90.200 1.800 92.400 ;
        RECT 1.200 82.200 2.000 90.200 ;
      LAYER via1 ;
        RECT 1.200 87.600 2.000 88.400 ;
      LAYER metal2 ;
        RECT 1.200 89.600 2.000 90.400 ;
        RECT 1.300 88.400 1.900 89.600 ;
        RECT 1.200 87.600 2.000 88.400 ;
      LAYER metal3 ;
        RECT 1.200 90.300 2.000 90.400 ;
        RECT -3.500 89.700 2.000 90.300 ;
        RECT 1.200 89.600 2.000 89.700 ;
    END
  END sr[4]
  PIN sr[3]
    PORT
      LAYER metal1 ;
        RECT 1.200 71.800 2.000 79.800 ;
        RECT 1.200 69.600 1.800 71.800 ;
        RECT 1.200 62.200 2.000 69.600 ;
      LAYER via1 ;
        RECT 1.200 73.600 2.000 74.400 ;
      LAYER metal2 ;
        RECT 1.200 73.600 2.000 74.400 ;
        RECT 1.300 72.400 1.900 73.600 ;
        RECT 1.200 71.600 2.000 72.400 ;
      LAYER metal3 ;
        RECT 1.200 72.300 2.000 72.400 ;
        RECT -3.500 71.700 2.000 72.300 ;
        RECT 1.200 71.600 2.000 71.700 ;
    END
  END sr[3]
  PIN sr[2]
    PORT
      LAYER metal1 ;
        RECT 1.200 52.400 2.000 59.800 ;
        RECT 1.200 50.200 1.800 52.400 ;
        RECT 1.200 42.200 2.000 50.200 ;
      LAYER via1 ;
        RECT 1.200 47.600 2.000 48.400 ;
      LAYER metal2 ;
        RECT 1.200 49.600 2.000 50.400 ;
        RECT 1.300 48.400 1.900 49.600 ;
        RECT 1.200 47.600 2.000 48.400 ;
      LAYER metal3 ;
        RECT 1.200 50.300 2.000 50.400 ;
        RECT -3.500 49.700 2.000 50.300 ;
        RECT 1.200 49.600 2.000 49.700 ;
    END
  END sr[2]
  PIN sr[1]
    PORT
      LAYER metal1 ;
        RECT 1.200 132.400 2.000 139.800 ;
        RECT 1.200 130.200 1.800 132.400 ;
        RECT 1.200 122.200 2.000 130.200 ;
      LAYER via1 ;
        RECT 1.200 127.600 2.000 128.400 ;
      LAYER metal2 ;
        RECT 1.200 129.600 2.000 130.400 ;
        RECT 1.300 128.400 1.900 129.600 ;
        RECT 1.200 127.600 2.000 128.400 ;
      LAYER metal3 ;
        RECT 1.200 130.300 2.000 130.400 ;
        RECT -3.500 129.700 2.000 130.300 ;
        RECT 1.200 129.600 2.000 129.700 ;
    END
  END sr[1]
  PIN sr[0]
    PORT
      LAYER metal1 ;
        RECT 1.200 151.800 2.000 159.800 ;
        RECT 1.200 149.600 1.800 151.800 ;
        RECT 1.200 142.200 2.000 149.600 ;
      LAYER via1 ;
        RECT 1.200 147.600 2.000 148.400 ;
      LAYER metal2 ;
        RECT 1.200 149.600 2.000 150.400 ;
        RECT 1.300 148.400 1.900 149.600 ;
        RECT 1.200 147.600 2.000 148.400 ;
      LAYER metal3 ;
        RECT 1.200 150.300 2.000 150.400 ;
        RECT -3.500 149.700 2.000 150.300 ;
        RECT 1.200 149.600 2.000 149.700 ;
    END
  END sr[0]
  PIN start
    PORT
      LAYER metal1 ;
        RECT 71.600 13.600 72.400 15.200 ;
      LAYER metal2 ;
        RECT 71.600 13.600 72.400 14.400 ;
        RECT 71.700 -1.700 72.300 13.600 ;
        RECT 71.700 -2.300 75.500 -1.700 ;
    END
  END start
  OBS
      LAYER metal1 ;
        RECT 4.400 175.200 5.200 179.800 ;
        RECT 7.600 176.000 8.400 179.800 ;
        RECT 3.000 174.600 5.200 175.200 ;
        RECT 7.400 175.200 8.400 176.000 ;
        RECT 3.000 171.600 3.600 174.600 ;
        RECT 4.400 172.300 5.200 173.200 ;
        RECT 7.400 172.300 8.200 175.200 ;
        RECT 9.200 174.600 10.000 179.800 ;
        RECT 15.600 176.600 16.400 179.800 ;
        RECT 17.200 177.000 18.000 179.800 ;
        RECT 18.800 177.000 19.600 179.800 ;
        RECT 20.400 177.000 21.200 179.800 ;
        RECT 22.000 177.000 22.800 179.800 ;
        RECT 25.200 177.000 26.000 179.800 ;
        RECT 28.400 177.000 29.200 179.800 ;
        RECT 30.000 177.000 30.800 179.800 ;
        RECT 31.600 177.000 32.400 179.800 ;
        RECT 14.000 175.800 16.400 176.600 ;
        RECT 33.200 176.600 34.000 179.800 ;
        RECT 14.000 175.200 14.800 175.800 ;
        RECT 4.400 171.700 8.200 172.300 ;
        RECT 4.400 171.600 5.200 171.700 ;
        RECT 2.400 170.800 3.600 171.600 ;
        RECT 3.000 170.200 3.600 170.800 ;
        RECT 7.400 170.800 8.200 171.700 ;
        RECT 8.800 174.000 10.000 174.600 ;
        RECT 13.000 174.600 14.800 175.200 ;
        RECT 18.800 175.600 19.800 176.400 ;
        RECT 22.800 175.600 24.400 176.400 ;
        RECT 25.200 175.800 29.800 176.400 ;
        RECT 33.200 175.800 35.800 176.600 ;
        RECT 25.200 175.600 26.000 175.800 ;
        RECT 8.800 172.000 9.400 174.000 ;
        RECT 13.000 173.400 13.800 174.600 ;
        RECT 10.000 172.600 13.800 173.400 ;
        RECT 18.800 172.800 19.600 175.600 ;
        RECT 25.200 174.800 26.000 175.000 ;
        RECT 21.600 174.200 26.000 174.800 ;
        RECT 21.600 174.000 22.400 174.200 ;
        RECT 26.800 173.600 27.600 175.200 ;
        RECT 29.000 173.400 29.800 175.800 ;
        RECT 35.000 175.200 35.800 175.800 ;
        RECT 35.000 174.400 38.000 175.200 ;
        RECT 39.600 173.800 40.400 179.800 ;
        RECT 42.800 177.800 43.600 179.800 ;
        RECT 41.200 175.600 42.000 177.200 ;
        RECT 43.000 176.300 43.600 177.800 ;
        RECT 46.200 176.400 47.000 177.200 ;
        RECT 46.000 176.300 46.800 176.400 ;
        RECT 42.900 175.700 46.800 176.300 ;
        RECT 47.600 175.800 48.400 179.800 ;
        RECT 43.000 174.400 43.600 175.700 ;
        RECT 46.000 175.600 46.800 175.700 ;
        RECT 22.000 172.600 25.200 173.400 ;
        RECT 29.000 172.600 31.000 173.400 ;
        RECT 31.600 173.000 40.400 173.800 ;
        RECT 42.800 173.600 43.600 174.400 ;
        RECT 15.600 172.000 16.400 172.600 ;
        RECT 33.200 172.000 34.000 172.400 ;
        RECT 34.800 172.000 35.600 172.400 ;
        RECT 38.200 172.000 39.000 172.200 ;
        RECT 8.800 171.400 9.600 172.000 ;
        RECT 15.600 171.400 39.000 172.000 ;
        RECT 3.000 169.600 5.200 170.200 ;
        RECT 7.400 170.000 8.400 170.800 ;
        RECT 4.400 162.200 5.200 169.600 ;
        RECT 7.600 162.200 8.400 170.000 ;
        RECT 9.000 169.600 9.600 171.400 ;
        RECT 9.000 169.000 18.000 169.600 ;
        RECT 9.000 167.400 9.600 169.000 ;
        RECT 17.200 168.800 18.000 169.000 ;
        RECT 20.400 169.000 29.000 169.600 ;
        RECT 20.400 168.800 21.200 169.000 ;
        RECT 12.200 167.600 14.800 168.400 ;
        RECT 9.000 166.800 11.600 167.400 ;
        RECT 10.800 162.200 11.600 166.800 ;
        RECT 14.000 162.200 14.800 167.600 ;
        RECT 15.400 166.800 19.600 167.600 ;
        RECT 17.200 162.200 18.000 165.000 ;
        RECT 18.800 162.200 19.600 165.000 ;
        RECT 20.400 162.200 21.200 165.000 ;
        RECT 22.000 162.200 22.800 168.400 ;
        RECT 25.200 167.600 27.800 168.400 ;
        RECT 28.400 168.200 29.000 169.000 ;
        RECT 30.000 169.400 30.800 169.600 ;
        RECT 30.000 169.000 35.400 169.400 ;
        RECT 30.000 168.800 36.200 169.000 ;
        RECT 34.800 168.200 36.200 168.800 ;
        RECT 28.400 167.600 34.200 168.200 ;
        RECT 37.200 168.000 38.800 168.800 ;
        RECT 37.200 167.600 37.800 168.000 ;
        RECT 25.200 162.200 26.000 167.000 ;
        RECT 28.400 162.200 29.200 167.000 ;
        RECT 33.600 166.800 37.800 167.600 ;
        RECT 39.600 167.400 40.400 173.000 ;
        RECT 43.000 170.200 43.600 173.600 ;
        RECT 44.400 170.800 45.200 172.400 ;
        RECT 46.000 172.200 46.800 172.400 ;
        RECT 47.800 172.200 48.400 175.800 ;
        RECT 55.600 175.200 56.400 179.800 ;
        RECT 54.200 174.600 56.400 175.200 ;
        RECT 49.200 172.800 50.000 174.400 ;
        RECT 50.800 172.200 51.600 172.400 ;
        RECT 46.000 171.600 48.400 172.200 ;
        RECT 50.000 171.600 51.600 172.200 ;
        RECT 54.200 171.600 54.800 174.600 ;
        RECT 63.600 173.800 64.400 179.800 ;
        RECT 70.000 176.600 70.800 179.800 ;
        RECT 71.600 177.000 72.400 179.800 ;
        RECT 73.200 177.000 74.000 179.800 ;
        RECT 74.800 177.000 75.600 179.800 ;
        RECT 78.000 177.000 78.800 179.800 ;
        RECT 81.200 177.000 82.000 179.800 ;
        RECT 82.800 177.000 83.600 179.800 ;
        RECT 84.400 177.000 85.200 179.800 ;
        RECT 86.000 177.000 86.800 179.800 ;
        RECT 68.200 175.800 70.800 176.600 ;
        RECT 87.600 176.600 88.400 179.800 ;
        RECT 74.200 175.800 78.800 176.400 ;
        RECT 68.200 175.200 69.000 175.800 ;
        RECT 66.000 174.400 69.000 175.200 ;
        RECT 55.600 171.600 56.400 173.200 ;
        RECT 63.600 173.000 72.400 173.800 ;
        RECT 74.200 173.400 75.000 175.800 ;
        RECT 78.000 175.600 78.800 175.800 ;
        RECT 79.600 175.600 81.200 176.400 ;
        RECT 84.200 175.600 85.200 176.400 ;
        RECT 87.600 175.800 90.000 176.600 ;
        RECT 76.400 173.600 77.200 175.200 ;
        RECT 78.000 174.800 78.800 175.000 ;
        RECT 78.000 174.200 82.400 174.800 ;
        RECT 81.600 174.000 82.400 174.200 ;
        RECT 46.200 170.200 46.800 171.600 ;
        RECT 50.000 171.200 50.800 171.600 ;
        RECT 53.600 170.800 54.800 171.600 ;
        RECT 54.200 170.200 54.800 170.800 ;
        RECT 42.800 169.400 44.600 170.200 ;
        RECT 38.400 166.800 40.400 167.400 ;
        RECT 30.000 162.200 30.800 165.000 ;
        RECT 31.600 162.200 32.400 165.000 ;
        RECT 34.800 162.200 35.600 166.800 ;
        RECT 38.400 166.200 39.000 166.800 ;
        RECT 38.000 165.600 39.000 166.200 ;
        RECT 38.000 162.200 38.800 165.600 ;
        RECT 43.800 162.200 44.600 169.400 ;
        RECT 46.000 162.200 46.800 170.200 ;
        RECT 47.600 169.600 51.600 170.200 ;
        RECT 54.200 169.600 56.400 170.200 ;
        RECT 47.600 162.200 48.400 169.600 ;
        RECT 50.800 162.200 51.600 169.600 ;
        RECT 55.600 162.200 56.400 169.600 ;
        RECT 63.600 167.400 64.400 173.000 ;
        RECT 73.000 172.600 75.000 173.400 ;
        RECT 78.800 172.600 82.000 173.400 ;
        RECT 84.400 172.800 85.200 175.600 ;
        RECT 89.200 175.200 90.000 175.800 ;
        RECT 89.200 174.600 91.000 175.200 ;
        RECT 90.200 173.400 91.000 174.600 ;
        RECT 94.000 174.600 94.800 179.800 ;
        RECT 95.600 176.000 96.400 179.800 ;
        RECT 95.600 175.200 96.600 176.000 ;
        RECT 94.000 174.000 95.200 174.600 ;
        RECT 90.200 172.600 94.000 173.400 ;
        RECT 65.000 172.000 65.800 172.200 ;
        RECT 66.800 172.000 67.600 172.400 ;
        RECT 70.000 172.000 70.800 172.400 ;
        RECT 87.600 172.000 88.400 172.600 ;
        RECT 94.600 172.000 95.200 174.000 ;
        RECT 65.000 171.400 88.400 172.000 ;
        RECT 94.400 171.400 95.200 172.000 ;
        RECT 95.800 172.300 96.600 175.200 ;
        RECT 98.800 175.200 99.600 179.800 ;
        RECT 106.800 175.200 107.600 179.800 ;
        RECT 110.000 176.000 110.800 179.800 ;
        RECT 98.800 174.600 101.000 175.200 ;
        RECT 98.800 172.300 99.600 173.200 ;
        RECT 95.800 171.700 99.600 172.300 ;
        RECT 94.400 169.600 95.000 171.400 ;
        RECT 95.800 170.800 96.600 171.700 ;
        RECT 98.800 171.600 99.600 171.700 ;
        RECT 100.400 171.600 101.000 174.600 ;
        RECT 105.400 174.600 107.600 175.200 ;
        RECT 109.800 175.200 110.800 176.000 ;
        RECT 105.400 171.600 106.000 174.600 ;
        RECT 106.800 172.300 107.600 173.200 ;
        RECT 109.800 172.300 110.600 175.200 ;
        RECT 111.600 174.600 112.400 179.800 ;
        RECT 118.000 176.600 118.800 179.800 ;
        RECT 119.600 177.000 120.400 179.800 ;
        RECT 121.200 177.000 122.000 179.800 ;
        RECT 122.800 177.000 123.600 179.800 ;
        RECT 124.400 177.000 125.200 179.800 ;
        RECT 127.600 177.000 128.400 179.800 ;
        RECT 130.800 177.000 131.600 179.800 ;
        RECT 132.400 177.000 133.200 179.800 ;
        RECT 134.000 177.000 134.800 179.800 ;
        RECT 116.400 175.800 118.800 176.600 ;
        RECT 135.600 176.600 136.400 179.800 ;
        RECT 116.400 175.200 117.200 175.800 ;
        RECT 106.800 171.700 110.600 172.300 ;
        RECT 106.800 171.600 107.600 171.700 ;
        RECT 73.200 169.400 74.000 169.600 ;
        RECT 68.600 169.000 74.000 169.400 ;
        RECT 67.800 168.800 74.000 169.000 ;
        RECT 75.000 169.000 83.600 169.600 ;
        RECT 65.200 168.000 66.800 168.800 ;
        RECT 67.800 168.200 69.200 168.800 ;
        RECT 75.000 168.200 75.600 169.000 ;
        RECT 82.800 168.800 83.600 169.000 ;
        RECT 86.000 169.000 95.000 169.600 ;
        RECT 86.000 168.800 86.800 169.000 ;
        RECT 66.200 167.600 66.800 168.000 ;
        RECT 69.800 167.600 75.600 168.200 ;
        RECT 76.200 167.600 78.800 168.400 ;
        RECT 63.600 166.800 65.600 167.400 ;
        RECT 66.200 166.800 70.400 167.600 ;
        RECT 65.000 166.200 65.600 166.800 ;
        RECT 65.000 165.600 66.000 166.200 ;
        RECT 65.200 162.200 66.000 165.600 ;
        RECT 68.400 162.200 69.200 166.800 ;
        RECT 71.600 162.200 72.400 165.000 ;
        RECT 73.200 162.200 74.000 165.000 ;
        RECT 74.800 162.200 75.600 167.000 ;
        RECT 78.000 162.200 78.800 167.000 ;
        RECT 81.200 162.200 82.000 168.400 ;
        RECT 89.200 167.600 91.800 168.400 ;
        RECT 84.400 166.800 88.600 167.600 ;
        RECT 82.800 162.200 83.600 165.000 ;
        RECT 84.400 162.200 85.200 165.000 ;
        RECT 86.000 162.200 86.800 165.000 ;
        RECT 89.200 162.200 90.000 167.600 ;
        RECT 94.400 167.400 95.000 169.000 ;
        RECT 92.400 166.800 95.000 167.400 ;
        RECT 95.600 170.000 96.600 170.800 ;
        RECT 100.400 170.800 101.600 171.600 ;
        RECT 104.800 170.800 106.000 171.600 ;
        RECT 100.400 170.200 101.000 170.800 ;
        RECT 92.400 162.200 93.200 166.800 ;
        RECT 95.600 162.200 96.400 170.000 ;
        RECT 98.800 169.600 101.000 170.200 ;
        RECT 105.400 170.200 106.000 170.800 ;
        RECT 109.800 170.800 110.600 171.700 ;
        RECT 111.200 174.000 112.400 174.600 ;
        RECT 115.400 174.600 117.200 175.200 ;
        RECT 121.200 175.600 122.200 176.400 ;
        RECT 125.200 175.600 126.800 176.400 ;
        RECT 127.600 175.800 132.200 176.400 ;
        RECT 135.600 175.800 138.200 176.600 ;
        RECT 127.600 175.600 128.400 175.800 ;
        RECT 111.200 172.000 111.800 174.000 ;
        RECT 115.400 173.400 116.200 174.600 ;
        RECT 112.400 172.600 116.200 173.400 ;
        RECT 121.200 172.800 122.000 175.600 ;
        RECT 127.600 174.800 128.400 175.000 ;
        RECT 124.000 174.200 128.400 174.800 ;
        RECT 124.000 174.000 124.800 174.200 ;
        RECT 129.200 173.600 130.000 175.200 ;
        RECT 131.400 173.400 132.200 175.800 ;
        RECT 137.400 175.200 138.200 175.800 ;
        RECT 137.400 174.400 140.400 175.200 ;
        RECT 142.000 173.800 142.800 179.800 ;
        RECT 143.600 175.200 144.400 179.800 ;
        RECT 148.400 175.200 149.200 179.800 ;
        RECT 143.600 174.600 145.800 175.200 ;
        RECT 148.400 174.600 150.600 175.200 ;
        RECT 124.400 172.600 127.600 173.400 ;
        RECT 131.400 172.600 133.400 173.400 ;
        RECT 134.000 173.000 142.800 173.800 ;
        RECT 118.000 172.000 118.800 172.600 ;
        RECT 135.600 172.000 136.400 172.400 ;
        RECT 138.800 172.000 139.600 172.400 ;
        RECT 140.600 172.000 141.400 172.200 ;
        RECT 111.200 171.400 112.000 172.000 ;
        RECT 118.000 171.400 141.400 172.000 ;
        RECT 105.400 169.600 107.600 170.200 ;
        RECT 109.800 170.000 110.800 170.800 ;
        RECT 98.800 162.200 99.600 169.600 ;
        RECT 106.800 162.200 107.600 169.600 ;
        RECT 110.000 162.200 110.800 170.000 ;
        RECT 111.400 169.600 112.000 171.400 ;
        RECT 111.400 169.000 120.400 169.600 ;
        RECT 111.400 167.400 112.000 169.000 ;
        RECT 119.600 168.800 120.400 169.000 ;
        RECT 122.800 169.000 131.400 169.600 ;
        RECT 122.800 168.800 123.600 169.000 ;
        RECT 114.600 167.600 117.200 168.400 ;
        RECT 111.400 166.800 114.000 167.400 ;
        RECT 113.200 162.200 114.000 166.800 ;
        RECT 116.400 162.200 117.200 167.600 ;
        RECT 117.800 166.800 122.000 167.600 ;
        RECT 119.600 162.200 120.400 165.000 ;
        RECT 121.200 162.200 122.000 165.000 ;
        RECT 122.800 162.200 123.600 165.000 ;
        RECT 124.400 162.200 125.200 168.400 ;
        RECT 127.600 167.600 130.200 168.400 ;
        RECT 130.800 168.200 131.400 169.000 ;
        RECT 132.400 169.400 133.200 169.600 ;
        RECT 132.400 169.000 137.800 169.400 ;
        RECT 132.400 168.800 138.600 169.000 ;
        RECT 137.200 168.200 138.600 168.800 ;
        RECT 130.800 167.600 136.600 168.200 ;
        RECT 139.600 168.000 141.200 168.800 ;
        RECT 139.600 167.600 140.200 168.000 ;
        RECT 127.600 162.200 128.400 167.000 ;
        RECT 130.800 162.200 131.600 167.000 ;
        RECT 136.000 166.800 140.200 167.600 ;
        RECT 142.000 167.400 142.800 173.000 ;
        RECT 143.600 171.600 144.400 173.200 ;
        RECT 145.200 171.600 145.800 174.600 ;
        RECT 148.400 171.600 149.200 173.200 ;
        RECT 150.000 171.600 150.600 174.600 ;
        RECT 153.200 173.800 154.000 179.800 ;
        RECT 159.600 176.600 160.400 179.800 ;
        RECT 161.200 177.000 162.000 179.800 ;
        RECT 162.800 177.000 163.600 179.800 ;
        RECT 164.400 177.000 165.200 179.800 ;
        RECT 167.600 177.000 168.400 179.800 ;
        RECT 170.800 177.000 171.600 179.800 ;
        RECT 172.400 177.000 173.200 179.800 ;
        RECT 174.000 177.000 174.800 179.800 ;
        RECT 175.600 177.000 176.400 179.800 ;
        RECT 157.800 175.800 160.400 176.600 ;
        RECT 177.200 176.600 178.000 179.800 ;
        RECT 163.800 175.800 168.400 176.400 ;
        RECT 157.800 175.200 158.600 175.800 ;
        RECT 155.600 174.400 158.600 175.200 ;
        RECT 153.200 173.000 162.000 173.800 ;
        RECT 163.800 173.400 164.600 175.800 ;
        RECT 167.600 175.600 168.400 175.800 ;
        RECT 169.200 175.600 170.800 176.400 ;
        RECT 173.800 175.600 174.800 176.400 ;
        RECT 177.200 175.800 179.600 176.600 ;
        RECT 166.000 173.600 166.800 175.200 ;
        RECT 167.600 174.800 168.400 175.000 ;
        RECT 167.600 174.200 172.000 174.800 ;
        RECT 171.200 174.000 172.000 174.200 ;
        RECT 145.200 170.800 146.400 171.600 ;
        RECT 150.000 170.800 151.200 171.600 ;
        RECT 145.200 170.200 145.800 170.800 ;
        RECT 150.000 170.200 150.600 170.800 ;
        RECT 140.800 166.800 142.800 167.400 ;
        RECT 143.600 169.600 145.800 170.200 ;
        RECT 148.400 169.600 150.600 170.200 ;
        RECT 132.400 162.200 133.200 165.000 ;
        RECT 134.000 162.200 134.800 165.000 ;
        RECT 137.200 162.200 138.000 166.800 ;
        RECT 140.800 166.200 141.400 166.800 ;
        RECT 140.400 165.600 141.400 166.200 ;
        RECT 140.400 162.200 141.200 165.600 ;
        RECT 143.600 162.200 144.400 169.600 ;
        RECT 148.400 162.200 149.200 169.600 ;
        RECT 153.200 167.400 154.000 173.000 ;
        RECT 162.600 172.600 164.600 173.400 ;
        RECT 168.400 172.600 171.600 173.400 ;
        RECT 174.000 172.800 174.800 175.600 ;
        RECT 178.800 175.200 179.600 175.800 ;
        RECT 178.800 174.600 180.600 175.200 ;
        RECT 179.800 173.400 180.600 174.600 ;
        RECT 183.600 174.600 184.400 179.800 ;
        RECT 185.200 176.000 186.000 179.800 ;
        RECT 185.200 175.200 186.200 176.000 ;
        RECT 183.600 174.000 184.800 174.600 ;
        RECT 179.800 172.600 183.600 173.400 ;
        RECT 154.600 172.000 155.400 172.200 ;
        RECT 159.600 172.000 160.400 172.400 ;
        RECT 166.000 172.000 166.800 172.400 ;
        RECT 177.200 172.000 178.000 172.600 ;
        RECT 184.200 172.000 184.800 174.000 ;
        RECT 154.600 171.400 178.000 172.000 ;
        RECT 184.000 171.400 184.800 172.000 ;
        RECT 185.400 172.300 186.200 175.200 ;
        RECT 194.800 175.200 195.600 179.800 ;
        RECT 194.800 174.600 197.000 175.200 ;
        RECT 194.800 172.300 195.600 173.200 ;
        RECT 185.400 171.700 195.600 172.300 ;
        RECT 184.000 169.600 184.600 171.400 ;
        RECT 185.400 170.800 186.200 171.700 ;
        RECT 194.800 171.600 195.600 171.700 ;
        RECT 196.400 171.600 197.000 174.600 ;
        RECT 199.600 173.800 200.400 179.800 ;
        RECT 206.000 176.600 206.800 179.800 ;
        RECT 207.600 177.000 208.400 179.800 ;
        RECT 209.200 177.000 210.000 179.800 ;
        RECT 210.800 177.000 211.600 179.800 ;
        RECT 214.000 177.000 214.800 179.800 ;
        RECT 217.200 177.000 218.000 179.800 ;
        RECT 218.800 177.000 219.600 179.800 ;
        RECT 220.400 177.000 221.200 179.800 ;
        RECT 222.000 177.000 222.800 179.800 ;
        RECT 204.200 175.800 206.800 176.600 ;
        RECT 223.600 176.600 224.400 179.800 ;
        RECT 210.200 175.800 214.800 176.400 ;
        RECT 204.200 175.200 205.000 175.800 ;
        RECT 202.000 174.400 205.000 175.200 ;
        RECT 199.600 173.000 208.400 173.800 ;
        RECT 210.200 173.400 211.000 175.800 ;
        RECT 214.000 175.600 214.800 175.800 ;
        RECT 215.600 175.600 217.200 176.400 ;
        RECT 220.200 175.600 221.200 176.400 ;
        RECT 223.600 175.800 226.000 176.600 ;
        RECT 212.400 173.600 213.200 175.200 ;
        RECT 214.000 174.800 214.800 175.000 ;
        RECT 214.000 174.200 218.400 174.800 ;
        RECT 217.600 174.000 218.400 174.200 ;
        RECT 162.800 169.400 163.600 169.600 ;
        RECT 158.200 169.000 163.600 169.400 ;
        RECT 157.400 168.800 163.600 169.000 ;
        RECT 164.600 169.000 173.200 169.600 ;
        RECT 154.800 168.000 156.400 168.800 ;
        RECT 157.400 168.200 158.800 168.800 ;
        RECT 164.600 168.200 165.200 169.000 ;
        RECT 172.400 168.800 173.200 169.000 ;
        RECT 175.600 169.000 184.600 169.600 ;
        RECT 175.600 168.800 176.400 169.000 ;
        RECT 155.800 167.600 156.400 168.000 ;
        RECT 159.400 167.600 165.200 168.200 ;
        RECT 165.800 167.600 168.400 168.400 ;
        RECT 153.200 166.800 155.200 167.400 ;
        RECT 155.800 166.800 160.000 167.600 ;
        RECT 154.600 166.200 155.200 166.800 ;
        RECT 154.600 165.600 155.600 166.200 ;
        RECT 154.800 162.200 155.600 165.600 ;
        RECT 158.000 162.200 158.800 166.800 ;
        RECT 161.200 162.200 162.000 165.000 ;
        RECT 162.800 162.200 163.600 165.000 ;
        RECT 164.400 162.200 165.200 167.000 ;
        RECT 167.600 162.200 168.400 167.000 ;
        RECT 170.800 162.200 171.600 168.400 ;
        RECT 178.800 167.600 181.400 168.400 ;
        RECT 174.000 166.800 178.200 167.600 ;
        RECT 172.400 162.200 173.200 165.000 ;
        RECT 174.000 162.200 174.800 165.000 ;
        RECT 175.600 162.200 176.400 165.000 ;
        RECT 178.800 162.200 179.600 167.600 ;
        RECT 184.000 167.400 184.600 169.000 ;
        RECT 182.000 166.800 184.600 167.400 ;
        RECT 185.200 170.000 186.200 170.800 ;
        RECT 196.400 170.800 197.600 171.600 ;
        RECT 196.400 170.200 197.000 170.800 ;
        RECT 182.000 162.200 182.800 166.800 ;
        RECT 185.200 162.200 186.000 170.000 ;
        RECT 194.800 169.600 197.000 170.200 ;
        RECT 194.800 162.200 195.600 169.600 ;
        RECT 199.600 167.400 200.400 173.000 ;
        RECT 209.000 172.600 211.000 173.400 ;
        RECT 214.800 172.600 218.000 173.400 ;
        RECT 220.400 172.800 221.200 175.600 ;
        RECT 225.200 175.200 226.000 175.800 ;
        RECT 225.200 174.600 227.000 175.200 ;
        RECT 226.200 173.400 227.000 174.600 ;
        RECT 230.000 174.600 230.800 179.800 ;
        RECT 231.600 176.000 232.400 179.800 ;
        RECT 231.600 175.200 232.600 176.000 ;
        RECT 230.000 174.000 231.200 174.600 ;
        RECT 226.200 172.600 230.000 173.400 ;
        RECT 201.000 172.000 201.800 172.200 ;
        RECT 202.800 172.000 203.600 172.400 ;
        RECT 206.000 172.000 206.800 172.400 ;
        RECT 223.600 172.000 224.400 172.600 ;
        RECT 230.600 172.000 231.200 174.000 ;
        RECT 201.000 171.400 224.400 172.000 ;
        RECT 230.400 171.400 231.200 172.000 ;
        RECT 231.800 172.300 232.600 175.200 ;
        RECT 234.800 175.200 235.600 179.800 ;
        RECT 241.200 177.800 242.000 179.800 ;
        RECT 234.800 174.600 237.000 175.200 ;
        RECT 234.800 172.300 235.600 173.200 ;
        RECT 231.800 171.700 235.600 172.300 ;
        RECT 230.400 169.600 231.000 171.400 ;
        RECT 231.800 170.800 232.600 171.700 ;
        RECT 234.800 171.600 235.600 171.700 ;
        RECT 236.400 171.600 237.000 174.600 ;
        RECT 241.400 174.400 242.000 177.800 ;
        RECT 245.000 176.400 245.800 179.800 ;
        RECT 245.000 175.800 246.800 176.400 ;
        RECT 241.200 173.600 242.000 174.400 ;
        RECT 242.800 174.300 243.600 174.400 ;
        RECT 246.000 174.300 246.800 175.800 ;
        RECT 249.200 175.200 250.000 179.800 ;
        RECT 249.200 174.600 251.400 175.200 ;
        RECT 242.800 173.700 246.800 174.300 ;
        RECT 242.800 173.600 243.600 173.700 ;
        RECT 209.200 169.400 210.000 169.600 ;
        RECT 204.600 169.000 210.000 169.400 ;
        RECT 203.800 168.800 210.000 169.000 ;
        RECT 211.000 169.000 219.600 169.600 ;
        RECT 201.200 168.000 202.800 168.800 ;
        RECT 203.800 168.200 205.200 168.800 ;
        RECT 211.000 168.200 211.600 169.000 ;
        RECT 218.800 168.800 219.600 169.000 ;
        RECT 222.000 169.000 231.000 169.600 ;
        RECT 222.000 168.800 222.800 169.000 ;
        RECT 202.200 167.600 202.800 168.000 ;
        RECT 205.800 167.600 211.600 168.200 ;
        RECT 212.200 167.600 214.800 168.400 ;
        RECT 199.600 166.800 201.600 167.400 ;
        RECT 202.200 166.800 206.400 167.600 ;
        RECT 201.000 166.200 201.600 166.800 ;
        RECT 201.000 165.600 202.000 166.200 ;
        RECT 201.200 162.200 202.000 165.600 ;
        RECT 204.400 162.200 205.200 166.800 ;
        RECT 207.600 162.200 208.400 165.000 ;
        RECT 209.200 162.200 210.000 165.000 ;
        RECT 210.800 162.200 211.600 167.000 ;
        RECT 214.000 162.200 214.800 167.000 ;
        RECT 217.200 162.200 218.000 168.400 ;
        RECT 225.200 167.600 227.800 168.400 ;
        RECT 220.400 166.800 224.600 167.600 ;
        RECT 218.800 162.200 219.600 165.000 ;
        RECT 220.400 162.200 221.200 165.000 ;
        RECT 222.000 162.200 222.800 165.000 ;
        RECT 225.200 162.200 226.000 167.600 ;
        RECT 230.400 167.400 231.000 169.000 ;
        RECT 228.400 166.800 231.000 167.400 ;
        RECT 231.600 170.000 232.600 170.800 ;
        RECT 236.400 170.800 237.600 171.600 ;
        RECT 236.400 170.200 237.000 170.800 ;
        RECT 241.400 170.200 242.000 173.600 ;
        RECT 228.400 162.200 229.200 166.800 ;
        RECT 231.600 162.200 232.400 170.000 ;
        RECT 234.800 169.600 237.000 170.200 ;
        RECT 234.800 162.200 235.600 169.600 ;
        RECT 241.200 169.400 243.000 170.200 ;
        RECT 242.200 164.400 243.000 169.400 ;
        RECT 241.200 163.600 243.000 164.400 ;
        RECT 242.200 162.200 243.000 163.600 ;
        RECT 246.000 162.200 246.800 173.700 ;
        RECT 249.200 171.600 250.000 173.200 ;
        RECT 250.800 171.600 251.400 174.600 ;
        RECT 250.800 170.800 252.000 171.600 ;
        RECT 250.800 170.200 251.400 170.800 ;
        RECT 249.200 169.600 251.400 170.200 ;
        RECT 249.200 162.200 250.000 169.600 ;
        RECT 4.400 152.400 5.200 159.800 ;
        RECT 3.000 151.800 5.200 152.400 ;
        RECT 7.600 152.000 8.400 159.800 ;
        RECT 10.800 155.200 11.600 159.800 ;
        RECT 3.000 151.200 3.600 151.800 ;
        RECT 2.400 150.400 3.600 151.200 ;
        RECT 7.400 151.200 8.400 152.000 ;
        RECT 9.000 154.600 11.600 155.200 ;
        RECT 9.000 153.000 9.600 154.600 ;
        RECT 14.000 154.400 14.800 159.800 ;
        RECT 17.200 157.000 18.000 159.800 ;
        RECT 18.800 157.000 19.600 159.800 ;
        RECT 20.400 157.000 21.200 159.800 ;
        RECT 15.400 154.400 19.600 155.200 ;
        RECT 12.200 153.600 14.800 154.400 ;
        RECT 22.000 153.600 22.800 159.800 ;
        RECT 25.200 155.000 26.000 159.800 ;
        RECT 28.400 155.000 29.200 159.800 ;
        RECT 30.000 157.000 30.800 159.800 ;
        RECT 31.600 157.000 32.400 159.800 ;
        RECT 34.800 155.200 35.600 159.800 ;
        RECT 38.000 156.400 38.800 159.800 ;
        RECT 38.000 155.800 39.000 156.400 ;
        RECT 38.400 155.200 39.000 155.800 ;
        RECT 33.600 154.400 37.800 155.200 ;
        RECT 38.400 154.600 40.400 155.200 ;
        RECT 25.200 153.600 27.800 154.400 ;
        RECT 28.400 153.800 34.200 154.400 ;
        RECT 37.200 154.000 37.800 154.400 ;
        RECT 17.200 153.000 18.000 153.200 ;
        RECT 9.000 152.400 18.000 153.000 ;
        RECT 20.400 153.000 21.200 153.200 ;
        RECT 28.400 153.000 29.000 153.800 ;
        RECT 34.800 153.200 36.200 153.800 ;
        RECT 37.200 153.200 38.800 154.000 ;
        RECT 20.400 152.400 29.000 153.000 ;
        RECT 30.000 153.000 36.200 153.200 ;
        RECT 30.000 152.600 35.400 153.000 ;
        RECT 30.000 152.400 30.800 152.600 ;
        RECT 3.000 147.400 3.600 150.400 ;
        RECT 4.400 150.300 5.200 150.400 ;
        RECT 7.400 150.300 8.200 151.200 ;
        RECT 9.000 150.600 9.600 152.400 ;
        RECT 4.400 149.700 8.200 150.300 ;
        RECT 4.400 148.800 5.200 149.700 ;
        RECT 3.000 146.800 5.200 147.400 ;
        RECT 4.400 142.200 5.200 146.800 ;
        RECT 7.400 146.800 8.200 149.700 ;
        RECT 8.800 150.000 9.600 150.600 ;
        RECT 15.600 150.000 39.000 150.600 ;
        RECT 8.800 148.000 9.400 150.000 ;
        RECT 15.600 149.400 16.400 150.000 ;
        RECT 33.200 149.600 34.000 150.000 ;
        RECT 34.800 149.600 35.600 150.000 ;
        RECT 38.200 149.800 39.000 150.000 ;
        RECT 10.000 148.600 13.800 149.400 ;
        RECT 8.800 147.400 10.000 148.000 ;
        RECT 7.400 146.000 8.400 146.800 ;
        RECT 7.600 142.200 8.400 146.000 ;
        RECT 9.200 142.200 10.000 147.400 ;
        RECT 13.000 147.400 13.800 148.600 ;
        RECT 13.000 146.800 14.800 147.400 ;
        RECT 14.000 146.200 14.800 146.800 ;
        RECT 18.800 146.400 19.600 149.200 ;
        RECT 22.000 148.600 25.200 149.400 ;
        RECT 29.000 148.600 31.000 149.400 ;
        RECT 39.600 149.000 40.400 154.600 ;
        RECT 21.600 147.800 22.400 148.000 ;
        RECT 21.600 147.200 26.000 147.800 ;
        RECT 25.200 147.000 26.000 147.200 ;
        RECT 26.800 146.800 27.600 148.400 ;
        RECT 14.000 145.400 16.400 146.200 ;
        RECT 18.800 145.600 19.800 146.400 ;
        RECT 22.800 145.600 24.400 146.400 ;
        RECT 25.200 146.200 26.000 146.400 ;
        RECT 29.000 146.200 29.800 148.600 ;
        RECT 31.600 148.200 40.400 149.000 ;
        RECT 35.000 146.800 38.000 147.600 ;
        RECT 35.000 146.200 35.800 146.800 ;
        RECT 25.200 145.600 29.800 146.200 ;
        RECT 15.600 142.200 16.400 145.400 ;
        RECT 33.200 145.400 35.800 146.200 ;
        RECT 17.200 142.200 18.000 145.000 ;
        RECT 18.800 142.200 19.600 145.000 ;
        RECT 20.400 142.200 21.200 145.000 ;
        RECT 22.000 142.200 22.800 145.000 ;
        RECT 25.200 142.200 26.000 145.000 ;
        RECT 28.400 142.200 29.200 145.000 ;
        RECT 30.000 142.200 30.800 145.000 ;
        RECT 31.600 142.200 32.400 145.000 ;
        RECT 33.200 142.200 34.000 145.400 ;
        RECT 39.600 142.200 40.400 148.200 ;
        RECT 41.200 144.800 42.000 146.400 ;
        RECT 42.800 142.200 43.600 159.800 ;
        RECT 46.000 156.400 46.800 159.800 ;
        RECT 45.800 155.800 46.800 156.400 ;
        RECT 45.800 155.200 46.400 155.800 ;
        RECT 49.200 155.200 50.000 159.800 ;
        RECT 52.400 157.000 53.200 159.800 ;
        RECT 54.000 157.000 54.800 159.800 ;
        RECT 44.400 154.600 46.400 155.200 ;
        RECT 44.400 149.000 45.200 154.600 ;
        RECT 47.000 154.400 51.200 155.200 ;
        RECT 55.600 155.000 56.400 159.800 ;
        RECT 58.800 155.000 59.600 159.800 ;
        RECT 47.000 154.000 47.600 154.400 ;
        RECT 46.000 153.200 47.600 154.000 ;
        RECT 50.600 153.800 56.400 154.400 ;
        RECT 48.600 153.200 50.000 153.800 ;
        RECT 48.600 153.000 54.800 153.200 ;
        RECT 49.400 152.600 54.800 153.000 ;
        RECT 54.000 152.400 54.800 152.600 ;
        RECT 55.800 153.000 56.400 153.800 ;
        RECT 57.000 153.600 59.600 154.400 ;
        RECT 62.000 153.600 62.800 159.800 ;
        RECT 63.600 157.000 64.400 159.800 ;
        RECT 65.200 157.000 66.000 159.800 ;
        RECT 66.800 157.000 67.600 159.800 ;
        RECT 65.200 154.400 69.400 155.200 ;
        RECT 70.000 154.400 70.800 159.800 ;
        RECT 73.200 155.200 74.000 159.800 ;
        RECT 73.200 154.600 75.800 155.200 ;
        RECT 70.000 153.600 72.600 154.400 ;
        RECT 63.600 153.000 64.400 153.200 ;
        RECT 55.800 152.400 64.400 153.000 ;
        RECT 66.800 153.000 67.600 153.200 ;
        RECT 75.200 153.000 75.800 154.600 ;
        RECT 66.800 152.400 75.800 153.000 ;
        RECT 75.200 150.600 75.800 152.400 ;
        RECT 76.400 152.000 77.200 159.800 ;
        RECT 86.000 152.400 86.800 159.800 ;
        RECT 89.200 152.400 90.000 159.800 ;
        RECT 76.400 151.200 77.400 152.000 ;
        RECT 86.000 151.800 90.000 152.400 ;
        RECT 90.800 151.800 91.600 159.800 ;
        RECT 95.000 152.600 95.800 159.800 ;
        RECT 94.000 151.800 95.800 152.600 ;
        RECT 97.200 152.400 98.000 159.800 ;
        RECT 100.400 152.400 101.200 159.800 ;
        RECT 97.200 151.800 101.200 152.400 ;
        RECT 102.000 151.800 102.800 159.800 ;
        RECT 103.600 152.400 104.400 159.800 ;
        RECT 103.600 151.800 105.800 152.400 ;
        RECT 106.800 151.800 107.600 159.800 ;
        RECT 109.000 152.600 109.800 159.800 ;
        RECT 109.000 151.800 110.800 152.600 ;
        RECT 113.200 152.400 114.000 159.800 ;
        RECT 120.600 152.600 121.400 159.800 ;
        RECT 113.200 151.800 115.400 152.400 ;
        RECT 119.600 151.800 121.400 152.600 ;
        RECT 122.800 151.800 123.600 159.800 ;
        RECT 124.400 152.400 125.200 159.800 ;
        RECT 127.600 152.400 128.400 159.800 ;
        RECT 124.400 151.800 128.400 152.400 ;
        RECT 45.800 150.000 69.200 150.600 ;
        RECT 75.200 150.000 76.000 150.600 ;
        RECT 45.800 149.800 46.600 150.000 ;
        RECT 47.600 149.600 48.400 150.000 ;
        RECT 50.800 149.600 51.600 150.000 ;
        RECT 68.400 149.400 69.200 150.000 ;
        RECT 44.400 148.200 53.200 149.000 ;
        RECT 53.800 148.600 55.800 149.400 ;
        RECT 59.600 148.600 62.800 149.400 ;
        RECT 44.400 142.200 45.200 148.200 ;
        RECT 46.800 146.800 49.800 147.600 ;
        RECT 49.000 146.200 49.800 146.800 ;
        RECT 55.000 146.200 55.800 148.600 ;
        RECT 57.200 146.800 58.000 148.400 ;
        RECT 62.400 147.800 63.200 148.000 ;
        RECT 58.800 147.200 63.200 147.800 ;
        RECT 58.800 147.000 59.600 147.200 ;
        RECT 65.200 146.400 66.000 149.200 ;
        RECT 71.000 148.600 74.800 149.400 ;
        RECT 71.000 147.400 71.800 148.600 ;
        RECT 75.400 148.000 76.000 150.000 ;
        RECT 58.800 146.200 59.600 146.400 ;
        RECT 49.000 145.400 51.600 146.200 ;
        RECT 55.000 145.600 59.600 146.200 ;
        RECT 60.400 145.600 62.000 146.400 ;
        RECT 65.000 145.600 66.000 146.400 ;
        RECT 70.000 146.800 71.800 147.400 ;
        RECT 74.800 147.400 76.000 148.000 ;
        RECT 70.000 146.200 70.800 146.800 ;
        RECT 50.800 142.200 51.600 145.400 ;
        RECT 68.400 145.400 70.800 146.200 ;
        RECT 52.400 142.200 53.200 145.000 ;
        RECT 54.000 142.200 54.800 145.000 ;
        RECT 55.600 142.200 56.400 145.000 ;
        RECT 58.800 142.200 59.600 145.000 ;
        RECT 62.000 142.200 62.800 145.000 ;
        RECT 63.600 142.200 64.400 145.000 ;
        RECT 65.200 142.200 66.000 145.000 ;
        RECT 66.800 142.200 67.600 145.000 ;
        RECT 68.400 142.200 69.200 145.400 ;
        RECT 74.800 142.200 75.600 147.400 ;
        RECT 76.600 146.800 77.400 151.200 ;
        RECT 86.800 150.400 87.600 150.800 ;
        RECT 90.800 150.400 91.400 151.800 ;
        RECT 86.000 149.800 87.600 150.400 ;
        RECT 89.200 149.800 91.600 150.400 ;
        RECT 86.000 149.600 86.800 149.800 ;
        RECT 78.000 148.300 78.800 148.400 ;
        RECT 87.600 148.300 88.400 149.200 ;
        RECT 78.000 147.700 88.400 148.300 ;
        RECT 78.000 147.600 78.800 147.700 ;
        RECT 87.600 147.600 88.400 147.700 ;
        RECT 76.400 146.000 77.400 146.800 ;
        RECT 89.200 146.200 89.800 149.800 ;
        RECT 90.800 149.600 91.600 149.800 ;
        RECT 94.200 148.400 94.800 151.800 ;
        RECT 95.600 149.600 96.400 151.200 ;
        RECT 98.000 150.400 98.800 150.800 ;
        RECT 102.000 150.400 102.600 151.800 ;
        RECT 105.200 151.200 105.800 151.800 ;
        RECT 105.200 150.400 106.400 151.200 ;
        RECT 97.200 149.800 98.800 150.400 ;
        RECT 100.400 149.800 102.800 150.400 ;
        RECT 97.200 149.600 98.000 149.800 ;
        RECT 94.000 148.300 94.800 148.400 ;
        RECT 90.900 147.700 94.800 148.300 ;
        RECT 95.700 148.300 96.300 149.600 ;
        RECT 98.800 148.300 99.600 149.200 ;
        RECT 95.700 147.700 99.600 148.300 ;
        RECT 90.900 146.400 91.500 147.700 ;
        RECT 94.000 147.600 94.800 147.700 ;
        RECT 98.800 147.600 99.600 147.700 ;
        RECT 76.400 142.200 77.200 146.000 ;
        RECT 89.200 142.200 90.000 146.200 ;
        RECT 90.800 145.600 91.600 146.400 ;
        RECT 90.600 144.800 91.400 145.600 ;
        RECT 92.400 144.800 93.200 146.400 ;
        RECT 94.200 144.200 94.800 147.600 ;
        RECT 94.000 142.200 94.800 144.200 ;
        RECT 100.400 146.200 101.000 149.800 ;
        RECT 102.000 149.600 102.800 149.800 ;
        RECT 103.600 148.800 104.400 150.400 ;
        RECT 105.200 147.400 105.800 150.400 ;
        RECT 107.000 149.600 107.600 151.800 ;
        RECT 108.400 149.600 109.200 151.200 ;
        RECT 103.600 146.800 105.800 147.400 ;
        RECT 106.800 148.300 107.600 149.600 ;
        RECT 108.500 148.300 109.100 149.600 ;
        RECT 106.800 147.700 109.100 148.300 ;
        RECT 110.000 148.400 110.600 151.800 ;
        RECT 114.800 151.200 115.400 151.800 ;
        RECT 114.800 150.400 116.000 151.200 ;
        RECT 111.600 150.300 112.400 150.400 ;
        RECT 113.200 150.300 114.000 150.400 ;
        RECT 111.600 149.700 114.000 150.300 ;
        RECT 111.600 149.600 112.400 149.700 ;
        RECT 113.200 148.800 114.000 149.700 ;
        RECT 100.400 142.200 101.200 146.200 ;
        RECT 102.000 145.600 102.800 146.400 ;
        RECT 101.800 144.800 102.600 145.600 ;
        RECT 103.600 142.200 104.400 146.800 ;
        RECT 106.800 142.200 107.600 147.700 ;
        RECT 110.000 147.600 110.800 148.400 ;
        RECT 108.400 146.300 109.200 146.400 ;
        RECT 110.000 146.300 110.600 147.600 ;
        RECT 114.800 147.400 115.400 150.400 ;
        RECT 119.800 148.400 120.400 151.800 ;
        RECT 121.200 149.600 122.000 151.200 ;
        RECT 123.000 150.400 123.600 151.800 ;
        RECT 126.800 150.400 127.600 150.800 ;
        RECT 122.800 149.800 125.200 150.400 ;
        RECT 126.800 150.300 128.400 150.400 ;
        RECT 129.200 150.300 130.000 159.800 ;
        RECT 132.400 152.400 133.200 159.800 ;
        RECT 132.400 151.800 134.600 152.400 ;
        RECT 134.000 151.200 134.600 151.800 ;
        RECT 134.000 150.400 135.200 151.200 ;
        RECT 126.800 149.800 130.000 150.300 ;
        RECT 122.800 149.600 123.600 149.800 ;
        RECT 119.600 147.600 120.400 148.400 ;
        RECT 113.200 146.800 115.400 147.400 ;
        RECT 108.400 145.700 110.700 146.300 ;
        RECT 108.400 145.600 109.200 145.700 ;
        RECT 110.000 144.200 110.600 145.700 ;
        RECT 111.600 144.800 112.400 146.400 ;
        RECT 110.000 142.200 110.800 144.200 ;
        RECT 113.200 142.200 114.000 146.800 ;
        RECT 118.000 144.800 118.800 146.400 ;
        RECT 119.800 146.300 120.400 147.600 ;
        RECT 122.800 146.300 123.600 146.400 ;
        RECT 119.700 145.700 123.600 146.300 ;
        RECT 124.600 146.200 125.200 149.800 ;
        RECT 127.600 149.700 130.000 149.800 ;
        RECT 127.600 149.600 128.400 149.700 ;
        RECT 126.000 147.600 126.800 149.200 ;
        RECT 119.800 144.200 120.400 145.700 ;
        RECT 122.800 145.600 123.600 145.700 ;
        RECT 123.000 144.800 123.800 145.600 ;
        RECT 119.600 142.200 120.400 144.200 ;
        RECT 124.400 142.200 125.200 146.200 ;
        RECT 129.200 142.200 130.000 149.700 ;
        RECT 132.400 148.800 133.200 150.400 ;
        RECT 134.000 147.400 134.600 150.400 ;
        RECT 132.400 146.800 134.600 147.400 ;
        RECT 137.200 146.800 138.000 148.400 ;
        RECT 130.800 144.800 131.600 146.400 ;
        RECT 132.400 142.200 133.200 146.800 ;
        RECT 138.800 146.200 139.600 159.800 ;
        RECT 143.600 156.400 144.400 159.800 ;
        RECT 143.400 155.800 144.400 156.400 ;
        RECT 143.400 155.200 144.000 155.800 ;
        RECT 146.800 155.200 147.600 159.800 ;
        RECT 150.000 157.000 150.800 159.800 ;
        RECT 151.600 157.000 152.400 159.800 ;
        RECT 142.000 154.600 144.000 155.200 ;
        RECT 140.400 151.600 141.200 153.200 ;
        RECT 142.000 149.000 142.800 154.600 ;
        RECT 144.600 154.400 148.800 155.200 ;
        RECT 153.200 155.000 154.000 159.800 ;
        RECT 156.400 155.000 157.200 159.800 ;
        RECT 144.600 154.000 145.200 154.400 ;
        RECT 143.600 153.200 145.200 154.000 ;
        RECT 148.200 153.800 154.000 154.400 ;
        RECT 146.200 153.200 147.600 153.800 ;
        RECT 146.200 153.000 152.400 153.200 ;
        RECT 147.000 152.600 152.400 153.000 ;
        RECT 151.600 152.400 152.400 152.600 ;
        RECT 153.400 153.000 154.000 153.800 ;
        RECT 154.600 153.600 157.200 154.400 ;
        RECT 159.600 153.600 160.400 159.800 ;
        RECT 161.200 157.000 162.000 159.800 ;
        RECT 162.800 157.000 163.600 159.800 ;
        RECT 164.400 157.000 165.200 159.800 ;
        RECT 162.800 154.400 167.000 155.200 ;
        RECT 167.600 154.400 168.400 159.800 ;
        RECT 170.800 155.200 171.600 159.800 ;
        RECT 170.800 154.600 173.400 155.200 ;
        RECT 167.600 153.600 170.200 154.400 ;
        RECT 161.200 153.000 162.000 153.200 ;
        RECT 153.400 152.400 162.000 153.000 ;
        RECT 164.400 153.000 165.200 153.200 ;
        RECT 172.800 153.000 173.400 154.600 ;
        RECT 164.400 152.400 173.400 153.000 ;
        RECT 172.800 150.600 173.400 152.400 ;
        RECT 174.000 152.000 174.800 159.800 ;
        RECT 180.400 152.400 181.200 159.800 ;
        RECT 184.600 158.400 185.400 159.800 ;
        RECT 183.600 157.600 185.400 158.400 ;
        RECT 174.000 151.200 175.000 152.000 ;
        RECT 179.000 151.800 181.200 152.400 ;
        RECT 184.600 152.400 185.400 157.600 ;
        RECT 186.000 153.600 186.800 154.400 ;
        RECT 186.200 152.400 186.800 153.600 ;
        RECT 184.600 151.800 185.600 152.400 ;
        RECT 186.200 151.800 187.600 152.400 ;
        RECT 179.000 151.200 179.600 151.800 ;
        RECT 143.400 150.000 166.800 150.600 ;
        RECT 172.800 150.000 173.600 150.600 ;
        RECT 143.400 149.800 144.200 150.000 ;
        RECT 146.800 149.600 147.600 150.000 ;
        RECT 148.400 149.600 149.200 150.000 ;
        RECT 166.000 149.400 166.800 150.000 ;
        RECT 142.000 148.200 150.800 149.000 ;
        RECT 151.400 148.600 153.400 149.400 ;
        RECT 157.200 148.600 160.400 149.400 ;
        RECT 138.800 145.600 140.600 146.200 ;
        RECT 139.800 144.400 140.600 145.600 ;
        RECT 138.800 143.600 140.600 144.400 ;
        RECT 139.800 142.200 140.600 143.600 ;
        RECT 142.000 142.200 142.800 148.200 ;
        RECT 144.400 146.800 147.400 147.600 ;
        RECT 146.600 146.200 147.400 146.800 ;
        RECT 152.600 146.200 153.400 148.600 ;
        RECT 154.800 146.800 155.600 148.400 ;
        RECT 160.000 147.800 160.800 148.000 ;
        RECT 156.400 147.200 160.800 147.800 ;
        RECT 156.400 147.000 157.200 147.200 ;
        RECT 162.800 146.400 163.600 149.200 ;
        RECT 168.600 148.600 172.400 149.400 ;
        RECT 168.600 147.400 169.400 148.600 ;
        RECT 173.000 148.000 173.600 150.000 ;
        RECT 156.400 146.200 157.200 146.400 ;
        RECT 146.600 145.400 149.200 146.200 ;
        RECT 152.600 145.600 157.200 146.200 ;
        RECT 158.000 145.600 159.600 146.400 ;
        RECT 162.600 145.600 163.600 146.400 ;
        RECT 167.600 146.800 169.400 147.400 ;
        RECT 172.400 147.400 173.600 148.000 ;
        RECT 167.600 146.200 168.400 146.800 ;
        RECT 148.400 142.200 149.200 145.400 ;
        RECT 166.000 145.400 168.400 146.200 ;
        RECT 150.000 142.200 150.800 145.000 ;
        RECT 151.600 142.200 152.400 145.000 ;
        RECT 153.200 142.200 154.000 145.000 ;
        RECT 156.400 142.200 157.200 145.000 ;
        RECT 159.600 142.200 160.400 145.000 ;
        RECT 161.200 142.200 162.000 145.000 ;
        RECT 162.800 142.200 163.600 145.000 ;
        RECT 164.400 142.200 165.200 145.000 ;
        RECT 166.000 142.200 166.800 145.400 ;
        RECT 172.400 142.200 173.200 147.400 ;
        RECT 174.200 146.800 175.000 151.200 ;
        RECT 178.400 150.400 179.600 151.200 ;
        RECT 179.000 147.400 179.600 150.400 ;
        RECT 180.400 148.800 181.200 150.400 ;
        RECT 183.600 148.800 184.400 150.400 ;
        RECT 185.000 148.400 185.600 151.800 ;
        RECT 186.800 151.600 187.600 151.800 ;
        RECT 194.800 151.600 195.600 153.200 ;
        RECT 186.900 150.300 187.500 151.600 ;
        RECT 196.400 150.300 197.200 159.800 ;
        RECT 202.200 152.600 203.000 159.800 ;
        RECT 201.200 151.800 203.000 152.600 ;
        RECT 186.900 149.700 197.200 150.300 ;
        RECT 182.000 148.200 182.800 148.400 ;
        RECT 182.000 147.600 183.600 148.200 ;
        RECT 185.000 147.600 187.600 148.400 ;
        RECT 179.000 146.800 181.200 147.400 ;
        RECT 182.800 147.200 183.600 147.600 ;
        RECT 174.000 146.000 175.000 146.800 ;
        RECT 174.000 142.200 174.800 146.000 ;
        RECT 180.400 142.200 181.200 146.800 ;
        RECT 182.200 146.200 185.800 146.600 ;
        RECT 186.800 146.200 187.400 147.600 ;
        RECT 196.400 146.200 197.200 149.700 ;
        RECT 201.400 148.400 202.000 151.800 ;
        RECT 204.400 151.600 205.200 153.200 ;
        RECT 202.800 149.600 203.600 151.200 ;
        RECT 198.000 148.300 198.800 148.400 ;
        RECT 198.000 147.700 200.300 148.300 ;
        RECT 198.000 146.800 198.800 147.700 ;
        RECT 199.700 146.400 200.300 147.700 ;
        RECT 201.200 147.600 202.000 148.400 ;
        RECT 182.000 146.000 186.000 146.200 ;
        RECT 182.000 142.200 182.800 146.000 ;
        RECT 185.200 142.200 186.000 146.000 ;
        RECT 186.800 142.200 187.600 146.200 ;
        RECT 195.400 145.600 197.200 146.200 ;
        RECT 195.400 142.200 196.200 145.600 ;
        RECT 199.600 144.800 200.400 146.400 ;
        RECT 201.400 146.300 202.000 147.600 ;
        RECT 202.800 146.300 203.600 146.400 ;
        RECT 201.300 145.700 203.600 146.300 ;
        RECT 206.000 146.200 206.800 159.800 ;
        RECT 211.800 152.400 212.600 159.800 ;
        RECT 213.200 153.600 214.000 154.400 ;
        RECT 213.400 152.400 214.000 153.600 ;
        RECT 211.800 151.800 212.800 152.400 ;
        RECT 213.400 151.800 214.800 152.400 ;
        RECT 212.200 150.400 212.800 151.800 ;
        RECT 214.000 151.600 214.800 151.800 ;
        RECT 215.600 151.600 216.400 153.200 ;
        RECT 210.800 148.800 211.600 150.400 ;
        RECT 212.200 149.600 213.200 150.400 ;
        RECT 214.100 150.300 214.700 151.600 ;
        RECT 217.200 150.300 218.000 159.800 ;
        RECT 220.400 152.400 221.200 159.800 ;
        RECT 221.800 152.400 222.600 152.600 ;
        RECT 220.400 151.800 222.600 152.400 ;
        RECT 224.800 152.400 226.400 159.800 ;
        RECT 228.400 152.400 229.200 152.600 ;
        RECT 230.000 152.400 230.800 159.800 ;
        RECT 224.800 151.800 226.800 152.400 ;
        RECT 228.400 151.800 230.800 152.400 ;
        RECT 234.200 152.400 235.000 159.800 ;
        RECT 235.600 153.600 236.400 154.400 ;
        RECT 235.800 152.400 236.400 153.600 ;
        RECT 240.600 152.400 241.400 159.800 ;
        RECT 234.200 151.800 235.200 152.400 ;
        RECT 235.800 151.800 237.200 152.400 ;
        RECT 222.000 151.200 222.600 151.800 ;
        RECT 222.000 150.600 225.400 151.200 ;
        RECT 224.600 150.400 225.400 150.600 ;
        RECT 226.200 150.400 226.800 151.800 ;
        RECT 214.100 149.700 218.000 150.300 ;
        RECT 212.200 148.400 212.800 149.600 ;
        RECT 207.600 146.800 208.400 148.400 ;
        RECT 209.200 148.200 210.000 148.400 ;
        RECT 209.200 147.600 210.800 148.200 ;
        RECT 212.200 147.600 214.800 148.400 ;
        RECT 210.000 147.200 210.800 147.600 ;
        RECT 209.400 146.200 213.000 146.600 ;
        RECT 214.000 146.200 214.600 147.600 ;
        RECT 217.200 146.200 218.000 149.700 ;
        RECT 222.400 149.800 223.200 150.000 ;
        RECT 226.200 149.800 227.600 150.400 ;
        RECT 222.400 149.200 225.000 149.800 ;
        RECT 224.400 148.600 225.000 149.200 ;
        RECT 225.800 149.600 227.600 149.800 ;
        RECT 225.800 149.200 226.800 149.600 ;
        RECT 218.800 146.800 219.600 148.400 ;
        RECT 220.400 148.200 222.000 148.400 ;
        RECT 220.400 147.600 223.800 148.200 ;
        RECT 224.400 147.800 225.200 148.600 ;
        RECT 223.200 147.200 223.800 147.600 ;
        RECT 221.800 146.800 222.600 147.000 ;
        RECT 201.400 144.200 202.000 145.700 ;
        RECT 202.800 145.600 203.600 145.700 ;
        RECT 205.000 145.600 206.800 146.200 ;
        RECT 209.200 146.000 213.200 146.200 ;
        RECT 201.200 142.200 202.000 144.200 ;
        RECT 205.000 144.400 205.800 145.600 ;
        RECT 205.000 143.600 206.800 144.400 ;
        RECT 205.000 142.200 205.800 143.600 ;
        RECT 209.200 142.200 210.000 146.000 ;
        RECT 212.400 142.200 213.200 146.000 ;
        RECT 214.000 142.200 214.800 146.200 ;
        RECT 216.200 145.600 218.000 146.200 ;
        RECT 220.400 146.200 222.600 146.800 ;
        RECT 223.200 146.600 225.200 147.200 ;
        RECT 223.600 146.400 225.200 146.600 ;
        RECT 216.200 142.200 217.000 145.600 ;
        RECT 220.400 142.200 221.200 146.200 ;
        RECT 225.800 145.800 226.400 149.200 ;
        RECT 233.200 148.800 234.000 150.400 ;
        RECT 234.600 148.400 235.200 151.800 ;
        RECT 236.400 151.600 237.200 151.800 ;
        RECT 239.600 151.600 241.600 152.400 ;
        RECT 236.400 150.300 237.200 150.400 ;
        RECT 239.600 150.300 240.400 150.400 ;
        RECT 236.400 149.700 240.400 150.300 ;
        RECT 236.400 149.600 237.200 149.700 ;
        RECT 239.600 148.800 240.400 149.700 ;
        RECT 241.000 148.400 241.600 151.600 ;
        RECT 227.200 147.600 228.000 148.400 ;
        RECT 231.600 148.200 232.400 148.400 ;
        RECT 231.600 147.600 233.200 148.200 ;
        RECT 234.600 147.600 237.200 148.400 ;
        RECT 241.000 147.600 243.600 148.400 ;
        RECT 227.200 147.200 227.800 147.600 ;
        RECT 232.400 147.200 233.200 147.600 ;
        RECT 227.000 146.400 227.800 147.200 ;
        RECT 228.400 146.800 229.200 147.000 ;
        RECT 228.400 146.200 230.800 146.800 ;
        RECT 231.800 146.200 235.400 146.600 ;
        RECT 236.400 146.200 237.000 147.600 ;
        RECT 238.200 146.200 241.800 146.600 ;
        RECT 242.800 146.200 243.400 147.600 ;
        RECT 224.800 144.400 226.400 145.800 ;
        RECT 223.600 143.600 226.400 144.400 ;
        RECT 224.800 142.200 226.400 143.600 ;
        RECT 230.000 142.200 230.800 146.200 ;
        RECT 231.600 146.000 235.600 146.200 ;
        RECT 231.600 142.200 232.400 146.000 ;
        RECT 234.800 142.200 235.600 146.000 ;
        RECT 236.400 142.200 237.200 146.200 ;
        RECT 238.000 146.000 242.000 146.200 ;
        RECT 238.000 142.200 238.800 146.000 ;
        RECT 241.200 142.200 242.000 146.000 ;
        RECT 242.800 142.200 243.600 146.200 ;
        RECT 244.400 142.200 245.200 159.800 ;
        RECT 250.200 152.600 251.000 159.800 ;
        RECT 249.200 151.800 251.000 152.600 ;
        RECT 249.400 148.400 250.000 151.800 ;
        RECT 249.200 148.300 250.000 148.400 ;
        RECT 246.100 147.700 250.000 148.300 ;
        RECT 246.100 146.400 246.700 147.700 ;
        RECT 249.200 147.600 250.000 147.700 ;
        RECT 246.000 144.800 246.800 146.400 ;
        RECT 249.400 144.400 250.000 147.600 ;
        RECT 249.200 142.200 250.000 144.400 ;
        RECT 4.400 135.200 5.200 139.800 ;
        RECT 7.600 136.000 8.400 139.800 ;
        RECT 3.000 134.600 5.200 135.200 ;
        RECT 7.400 135.200 8.400 136.000 ;
        RECT 3.000 131.600 3.600 134.600 ;
        RECT 4.400 132.300 5.200 133.200 ;
        RECT 7.400 132.300 8.200 135.200 ;
        RECT 9.200 134.600 10.000 139.800 ;
        RECT 15.600 136.600 16.400 139.800 ;
        RECT 17.200 137.000 18.000 139.800 ;
        RECT 18.800 137.000 19.600 139.800 ;
        RECT 20.400 137.000 21.200 139.800 ;
        RECT 22.000 137.000 22.800 139.800 ;
        RECT 25.200 137.000 26.000 139.800 ;
        RECT 28.400 137.000 29.200 139.800 ;
        RECT 30.000 137.000 30.800 139.800 ;
        RECT 31.600 137.000 32.400 139.800 ;
        RECT 14.000 135.800 16.400 136.600 ;
        RECT 33.200 136.600 34.000 139.800 ;
        RECT 14.000 135.200 14.800 135.800 ;
        RECT 4.400 131.700 8.200 132.300 ;
        RECT 4.400 131.600 5.200 131.700 ;
        RECT 2.400 130.800 3.600 131.600 ;
        RECT 3.000 130.200 3.600 130.800 ;
        RECT 7.400 130.800 8.200 131.700 ;
        RECT 8.800 134.000 10.000 134.600 ;
        RECT 13.000 134.600 14.800 135.200 ;
        RECT 18.800 135.600 19.800 136.400 ;
        RECT 22.800 135.600 24.400 136.400 ;
        RECT 25.200 135.800 29.800 136.400 ;
        RECT 33.200 135.800 35.800 136.600 ;
        RECT 25.200 135.600 26.000 135.800 ;
        RECT 8.800 132.000 9.400 134.000 ;
        RECT 13.000 133.400 13.800 134.600 ;
        RECT 10.000 132.600 13.800 133.400 ;
        RECT 18.800 132.800 19.600 135.600 ;
        RECT 25.200 134.800 26.000 135.000 ;
        RECT 21.600 134.200 26.000 134.800 ;
        RECT 21.600 134.000 22.400 134.200 ;
        RECT 26.800 133.600 27.600 135.200 ;
        RECT 29.000 133.400 29.800 135.800 ;
        RECT 35.000 135.200 35.800 135.800 ;
        RECT 35.000 134.400 38.000 135.200 ;
        RECT 39.600 133.800 40.400 139.800 ;
        RECT 41.200 135.600 42.000 137.200 ;
        RECT 22.000 132.600 25.200 133.400 ;
        RECT 29.000 132.600 31.000 133.400 ;
        RECT 31.600 133.000 40.400 133.800 ;
        RECT 15.600 132.000 16.400 132.600 ;
        RECT 33.200 132.000 34.000 132.400 ;
        RECT 34.800 132.000 35.600 132.400 ;
        RECT 38.200 132.000 39.000 132.200 ;
        RECT 8.800 131.400 9.600 132.000 ;
        RECT 15.600 131.400 39.000 132.000 ;
        RECT 3.000 129.600 5.200 130.200 ;
        RECT 7.400 130.000 8.400 130.800 ;
        RECT 4.400 122.200 5.200 129.600 ;
        RECT 7.600 122.200 8.400 130.000 ;
        RECT 9.000 129.600 9.600 131.400 ;
        RECT 9.000 129.000 18.000 129.600 ;
        RECT 9.000 127.400 9.600 129.000 ;
        RECT 17.200 128.800 18.000 129.000 ;
        RECT 20.400 129.000 29.000 129.600 ;
        RECT 20.400 128.800 21.200 129.000 ;
        RECT 12.200 127.600 14.800 128.400 ;
        RECT 9.000 126.800 11.600 127.400 ;
        RECT 10.800 122.200 11.600 126.800 ;
        RECT 14.000 122.200 14.800 127.600 ;
        RECT 15.400 126.800 19.600 127.600 ;
        RECT 17.200 122.200 18.000 125.000 ;
        RECT 18.800 122.200 19.600 125.000 ;
        RECT 20.400 122.200 21.200 125.000 ;
        RECT 22.000 122.200 22.800 128.400 ;
        RECT 25.200 127.600 27.800 128.400 ;
        RECT 28.400 128.200 29.000 129.000 ;
        RECT 30.000 129.400 30.800 129.600 ;
        RECT 30.000 129.000 35.400 129.400 ;
        RECT 30.000 128.800 36.200 129.000 ;
        RECT 34.800 128.200 36.200 128.800 ;
        RECT 28.400 127.600 34.200 128.200 ;
        RECT 37.200 128.000 38.800 128.800 ;
        RECT 37.200 127.600 37.800 128.000 ;
        RECT 25.200 122.200 26.000 127.000 ;
        RECT 28.400 122.200 29.200 127.000 ;
        RECT 33.600 126.800 37.800 127.600 ;
        RECT 39.600 127.400 40.400 133.000 ;
        RECT 38.400 126.800 40.400 127.400 ;
        RECT 42.800 134.300 43.600 139.800 ;
        RECT 44.400 136.000 45.200 139.800 ;
        RECT 47.600 139.200 51.600 139.800 ;
        RECT 47.600 136.000 48.400 139.200 ;
        RECT 44.400 135.800 48.400 136.000 ;
        RECT 49.200 135.800 50.000 138.600 ;
        RECT 50.800 135.800 51.600 139.200 ;
        RECT 52.400 136.000 53.200 139.800 ;
        RECT 55.600 139.200 59.600 139.800 ;
        RECT 55.600 136.000 56.400 139.200 ;
        RECT 52.400 135.800 56.400 136.000 ;
        RECT 57.200 135.800 58.000 138.600 ;
        RECT 58.800 135.800 59.600 139.200 ;
        RECT 44.600 135.400 48.200 135.800 ;
        RECT 45.200 134.400 46.000 134.800 ;
        RECT 49.400 134.400 50.000 135.800 ;
        RECT 52.600 135.400 56.200 135.800 ;
        RECT 53.200 134.400 54.000 134.800 ;
        RECT 57.400 134.400 58.000 135.800 ;
        RECT 44.400 134.300 46.000 134.400 ;
        RECT 42.800 133.800 46.000 134.300 ;
        RECT 47.600 133.800 50.000 134.400 ;
        RECT 50.800 134.300 51.600 134.400 ;
        RECT 52.400 134.300 54.000 134.400 ;
        RECT 50.800 133.800 54.000 134.300 ;
        RECT 55.600 133.800 58.000 134.400 ;
        RECT 42.800 133.700 45.200 133.800 ;
        RECT 30.000 122.200 30.800 125.000 ;
        RECT 31.600 122.200 32.400 125.000 ;
        RECT 34.800 122.200 35.600 126.800 ;
        RECT 38.400 126.200 39.000 126.800 ;
        RECT 38.000 125.600 39.000 126.200 ;
        RECT 38.000 122.200 38.800 125.600 ;
        RECT 42.800 122.200 43.600 133.700 ;
        RECT 44.400 133.600 45.200 133.700 ;
        RECT 47.600 133.600 48.400 133.800 ;
        RECT 50.800 133.700 53.200 133.800 ;
        RECT 46.000 131.600 46.800 133.200 ;
        RECT 47.600 130.200 48.200 133.600 ;
        RECT 49.200 131.600 50.000 133.200 ;
        RECT 50.800 132.800 51.600 133.700 ;
        RECT 52.400 133.600 53.200 133.700 ;
        RECT 55.600 133.600 56.400 133.800 ;
        RECT 54.000 131.600 54.800 133.200 ;
        RECT 55.600 130.200 56.200 133.600 ;
        RECT 57.200 131.600 58.000 133.200 ;
        RECT 58.800 132.800 59.600 134.400 ;
        RECT 60.400 134.300 61.200 139.800 ;
        RECT 62.000 136.300 62.800 137.200 ;
        RECT 68.400 136.300 69.200 136.400 ;
        RECT 62.000 135.700 69.200 136.300 ;
        RECT 70.000 136.000 70.800 139.800 ;
        RECT 73.200 139.200 77.200 139.800 ;
        RECT 73.200 136.000 74.000 139.200 ;
        RECT 70.000 135.800 74.000 136.000 ;
        RECT 74.800 135.800 75.600 138.600 ;
        RECT 76.400 135.800 77.200 139.200 ;
        RECT 62.000 135.600 62.800 135.700 ;
        RECT 68.400 135.600 69.200 135.700 ;
        RECT 70.200 135.400 73.800 135.800 ;
        RECT 70.800 134.400 71.600 134.800 ;
        RECT 75.000 134.400 75.600 135.800 ;
        RECT 70.000 134.300 71.600 134.400 ;
        RECT 60.400 133.800 71.600 134.300 ;
        RECT 73.200 133.800 75.600 134.400 ;
        RECT 60.400 133.700 70.800 133.800 ;
        RECT 47.000 122.200 49.000 130.200 ;
        RECT 55.000 122.200 57.000 130.200 ;
        RECT 60.400 122.200 61.200 133.700 ;
        RECT 70.000 133.600 70.800 133.700 ;
        RECT 73.200 133.600 74.000 133.800 ;
        RECT 62.000 132.300 62.800 132.400 ;
        RECT 71.600 132.300 72.400 133.200 ;
        RECT 62.000 131.700 72.400 132.300 ;
        RECT 62.000 131.600 62.800 131.700 ;
        RECT 71.600 131.600 72.400 131.700 ;
        RECT 73.200 130.200 73.800 133.600 ;
        RECT 74.800 131.600 75.600 133.200 ;
        RECT 76.400 132.800 77.200 134.400 ;
        RECT 78.000 132.400 78.800 139.800 ;
        RECT 81.200 135.200 82.000 139.800 ;
        RECT 79.800 134.600 82.000 135.200 ;
        RECT 78.000 130.200 78.600 132.400 ;
        RECT 79.800 131.600 80.400 134.600 ;
        RECT 82.800 133.800 83.600 139.800 ;
        RECT 89.200 136.600 90.000 139.800 ;
        RECT 90.800 137.000 91.600 139.800 ;
        RECT 92.400 137.000 93.200 139.800 ;
        RECT 94.000 137.000 94.800 139.800 ;
        RECT 97.200 137.000 98.000 139.800 ;
        RECT 100.400 137.000 101.200 139.800 ;
        RECT 102.000 137.000 102.800 139.800 ;
        RECT 103.600 137.000 104.400 139.800 ;
        RECT 105.200 137.000 106.000 139.800 ;
        RECT 87.400 135.800 90.000 136.600 ;
        RECT 106.800 136.600 107.600 139.800 ;
        RECT 93.400 135.800 98.000 136.400 ;
        RECT 87.400 135.200 88.200 135.800 ;
        RECT 85.200 134.400 88.200 135.200 ;
        RECT 81.200 131.600 82.000 133.200 ;
        RECT 82.800 133.000 91.600 133.800 ;
        RECT 93.400 133.400 94.200 135.800 ;
        RECT 97.200 135.600 98.000 135.800 ;
        RECT 98.800 135.600 100.400 136.400 ;
        RECT 103.400 135.600 104.400 136.400 ;
        RECT 106.800 135.800 109.200 136.600 ;
        RECT 95.600 133.600 96.400 135.200 ;
        RECT 97.200 134.800 98.000 135.000 ;
        RECT 97.200 134.200 101.600 134.800 ;
        RECT 100.800 134.000 101.600 134.200 ;
        RECT 79.200 130.800 80.400 131.600 ;
        RECT 79.800 130.200 80.400 130.800 ;
        RECT 72.600 122.200 74.600 130.200 ;
        RECT 78.000 122.200 78.800 130.200 ;
        RECT 79.800 129.600 82.000 130.200 ;
        RECT 81.200 122.200 82.000 129.600 ;
        RECT 82.800 127.400 83.600 133.000 ;
        RECT 92.200 132.600 94.200 133.400 ;
        RECT 98.000 132.600 101.200 133.400 ;
        RECT 103.600 132.800 104.400 135.600 ;
        RECT 108.400 135.200 109.200 135.800 ;
        RECT 108.400 134.600 110.200 135.200 ;
        RECT 109.400 133.400 110.200 134.600 ;
        RECT 113.200 134.600 114.000 139.800 ;
        RECT 114.800 136.000 115.600 139.800 ;
        RECT 119.600 136.000 120.400 139.800 ;
        RECT 114.800 135.200 115.800 136.000 ;
        RECT 113.200 134.000 114.400 134.600 ;
        RECT 109.400 132.600 113.200 133.400 ;
        RECT 84.200 132.000 85.000 132.200 ;
        RECT 89.200 132.000 90.000 132.400 ;
        RECT 106.800 132.000 107.600 132.600 ;
        RECT 113.800 132.000 114.400 134.000 ;
        RECT 84.200 131.400 107.600 132.000 ;
        RECT 113.600 131.400 114.400 132.000 ;
        RECT 113.600 129.600 114.200 131.400 ;
        RECT 115.000 130.800 115.800 135.200 ;
        RECT 92.400 129.400 93.200 129.600 ;
        RECT 87.800 129.000 93.200 129.400 ;
        RECT 87.000 128.800 93.200 129.000 ;
        RECT 94.200 129.000 102.800 129.600 ;
        RECT 84.400 128.000 86.000 128.800 ;
        RECT 87.000 128.200 88.400 128.800 ;
        RECT 94.200 128.200 94.800 129.000 ;
        RECT 102.000 128.800 102.800 129.000 ;
        RECT 105.200 129.000 114.200 129.600 ;
        RECT 105.200 128.800 106.000 129.000 ;
        RECT 85.400 127.600 86.000 128.000 ;
        RECT 89.000 127.600 94.800 128.200 ;
        RECT 95.400 127.600 98.000 128.400 ;
        RECT 82.800 126.800 84.800 127.400 ;
        RECT 85.400 126.800 89.600 127.600 ;
        RECT 84.200 126.200 84.800 126.800 ;
        RECT 84.200 125.600 85.200 126.200 ;
        RECT 84.400 122.200 85.200 125.600 ;
        RECT 87.600 122.200 88.400 126.800 ;
        RECT 90.800 122.200 91.600 125.000 ;
        RECT 92.400 122.200 93.200 125.000 ;
        RECT 94.000 122.200 94.800 127.000 ;
        RECT 97.200 122.200 98.000 127.000 ;
        RECT 100.400 122.200 101.200 128.400 ;
        RECT 108.400 127.600 111.000 128.400 ;
        RECT 103.600 126.800 107.800 127.600 ;
        RECT 102.000 122.200 102.800 125.000 ;
        RECT 103.600 122.200 104.400 125.000 ;
        RECT 105.200 122.200 106.000 125.000 ;
        RECT 108.400 122.200 109.200 127.600 ;
        RECT 113.600 127.400 114.200 129.000 ;
        RECT 111.600 126.800 114.200 127.400 ;
        RECT 114.800 130.000 115.800 130.800 ;
        RECT 119.400 135.200 120.400 136.000 ;
        RECT 119.400 130.800 120.200 135.200 ;
        RECT 121.200 134.600 122.000 139.800 ;
        RECT 127.600 136.600 128.400 139.800 ;
        RECT 129.200 137.000 130.000 139.800 ;
        RECT 130.800 137.000 131.600 139.800 ;
        RECT 132.400 137.000 133.200 139.800 ;
        RECT 134.000 137.000 134.800 139.800 ;
        RECT 137.200 137.000 138.000 139.800 ;
        RECT 140.400 137.000 141.200 139.800 ;
        RECT 142.000 137.000 142.800 139.800 ;
        RECT 143.600 137.000 144.400 139.800 ;
        RECT 126.000 135.800 128.400 136.600 ;
        RECT 145.200 136.600 146.000 139.800 ;
        RECT 126.000 135.200 126.800 135.800 ;
        RECT 120.800 134.000 122.000 134.600 ;
        RECT 125.000 134.600 126.800 135.200 ;
        RECT 130.800 135.600 131.800 136.400 ;
        RECT 134.800 135.600 136.400 136.400 ;
        RECT 137.200 135.800 141.800 136.400 ;
        RECT 145.200 135.800 147.800 136.600 ;
        RECT 137.200 135.600 138.000 135.800 ;
        RECT 120.800 132.000 121.400 134.000 ;
        RECT 125.000 133.400 125.800 134.600 ;
        RECT 122.000 132.600 125.800 133.400 ;
        RECT 130.800 132.800 131.600 135.600 ;
        RECT 137.200 134.800 138.000 135.000 ;
        RECT 133.600 134.200 138.000 134.800 ;
        RECT 133.600 134.000 134.400 134.200 ;
        RECT 138.800 133.600 139.600 135.200 ;
        RECT 141.000 133.400 141.800 135.800 ;
        RECT 147.000 135.200 147.800 135.800 ;
        RECT 147.000 134.400 150.000 135.200 ;
        RECT 151.600 133.800 152.400 139.800 ;
        RECT 134.000 132.600 137.200 133.400 ;
        RECT 141.000 132.600 143.000 133.400 ;
        RECT 143.600 133.000 152.400 133.800 ;
        RECT 127.600 132.000 128.400 132.600 ;
        RECT 145.200 132.000 146.000 132.400 ;
        RECT 146.800 132.000 147.600 132.400 ;
        RECT 150.200 132.000 151.000 132.200 ;
        RECT 120.800 131.400 121.600 132.000 ;
        RECT 127.600 131.400 151.000 132.000 ;
        RECT 119.400 130.000 120.400 130.800 ;
        RECT 111.600 122.200 112.400 126.800 ;
        RECT 114.800 122.200 115.600 130.000 ;
        RECT 119.600 122.200 120.400 130.000 ;
        RECT 121.000 129.600 121.600 131.400 ;
        RECT 121.000 129.000 130.000 129.600 ;
        RECT 121.000 127.400 121.600 129.000 ;
        RECT 129.200 128.800 130.000 129.000 ;
        RECT 132.400 129.000 141.000 129.600 ;
        RECT 132.400 128.800 133.200 129.000 ;
        RECT 124.200 127.600 126.800 128.400 ;
        RECT 121.000 126.800 123.600 127.400 ;
        RECT 122.800 122.200 123.600 126.800 ;
        RECT 126.000 122.200 126.800 127.600 ;
        RECT 127.400 126.800 131.600 127.600 ;
        RECT 129.200 122.200 130.000 125.000 ;
        RECT 130.800 122.200 131.600 125.000 ;
        RECT 132.400 122.200 133.200 125.000 ;
        RECT 134.000 122.200 134.800 128.400 ;
        RECT 137.200 127.600 139.800 128.400 ;
        RECT 140.400 128.200 141.000 129.000 ;
        RECT 142.000 129.400 142.800 129.600 ;
        RECT 142.000 129.000 147.400 129.400 ;
        RECT 142.000 128.800 148.200 129.000 ;
        RECT 146.800 128.200 148.200 128.800 ;
        RECT 140.400 127.600 146.200 128.200 ;
        RECT 149.200 128.000 150.800 128.800 ;
        RECT 149.200 127.600 149.800 128.000 ;
        RECT 137.200 122.200 138.000 127.000 ;
        RECT 140.400 122.200 141.200 127.000 ;
        RECT 145.600 126.800 149.800 127.600 ;
        RECT 151.600 127.400 152.400 133.000 ;
        RECT 150.400 126.800 152.400 127.400 ;
        RECT 142.000 122.200 142.800 125.000 ;
        RECT 143.600 122.200 144.400 125.000 ;
        RECT 146.800 122.200 147.600 126.800 ;
        RECT 150.400 126.200 151.000 126.800 ;
        RECT 150.000 125.600 151.000 126.200 ;
        RECT 150.000 122.200 150.800 125.600 ;
        RECT 154.800 122.200 155.600 139.800 ;
        RECT 161.200 135.800 162.000 139.800 ;
        RECT 164.400 139.200 168.400 139.800 ;
        RECT 162.600 136.400 163.400 137.200 ;
        RECT 156.400 134.300 157.200 135.200 ;
        RECT 159.600 134.300 160.400 134.400 ;
        RECT 156.400 133.700 160.400 134.300 ;
        RECT 156.400 133.600 157.200 133.700 ;
        RECT 159.600 132.800 160.400 133.700 ;
        RECT 158.000 132.200 158.800 132.400 ;
        RECT 161.200 132.200 161.800 135.800 ;
        RECT 162.800 135.600 163.600 136.400 ;
        RECT 164.400 135.800 165.200 139.200 ;
        RECT 166.000 135.600 166.800 138.600 ;
        RECT 167.600 136.000 168.400 139.200 ;
        RECT 170.800 136.000 171.600 139.800 ;
        RECT 167.600 135.800 171.600 136.000 ;
        RECT 166.000 134.400 166.600 135.600 ;
        RECT 167.800 135.400 171.400 135.800 ;
        RECT 170.000 134.400 170.800 134.800 ;
        RECT 164.400 132.800 165.200 134.400 ;
        RECT 166.000 133.800 168.400 134.400 ;
        RECT 170.000 133.800 171.600 134.400 ;
        RECT 167.600 133.600 168.400 133.800 ;
        RECT 170.800 133.600 171.600 133.800 ;
        RECT 162.800 132.200 163.600 132.400 ;
        RECT 158.000 131.600 159.600 132.200 ;
        RECT 161.200 131.600 163.600 132.200 ;
        RECT 166.000 131.600 166.800 133.200 ;
        RECT 158.800 131.200 159.600 131.600 ;
        RECT 162.800 130.200 163.400 131.600 ;
        RECT 167.800 130.200 168.400 133.600 ;
        RECT 169.200 132.300 170.000 133.200 ;
        RECT 174.000 132.300 174.800 139.800 ;
        RECT 177.200 136.000 178.000 139.800 ;
        RECT 180.400 136.000 181.200 139.800 ;
        RECT 177.200 135.800 181.200 136.000 ;
        RECT 182.000 135.800 182.800 139.800 ;
        RECT 193.200 135.800 194.000 139.800 ;
        RECT 198.000 137.800 198.800 139.800 ;
        RECT 194.600 136.400 195.400 137.200 ;
        RECT 177.400 135.400 181.000 135.800 ;
        RECT 175.600 133.600 176.400 135.200 ;
        RECT 178.000 134.400 178.800 134.800 ;
        RECT 182.000 134.400 182.600 135.800 ;
        RECT 177.200 133.800 178.800 134.400 ;
        RECT 177.200 133.600 178.000 133.800 ;
        RECT 180.200 133.600 182.800 134.400 ;
        RECT 169.200 131.700 174.800 132.300 ;
        RECT 169.200 131.600 170.000 131.700 ;
        RECT 158.000 129.600 162.000 130.200 ;
        RECT 158.000 122.200 158.800 129.600 ;
        RECT 161.200 122.200 162.000 129.600 ;
        RECT 162.800 122.200 163.600 130.200 ;
        RECT 167.000 122.200 169.000 130.200 ;
        RECT 174.000 122.200 174.800 131.700 ;
        RECT 177.200 132.300 178.000 132.400 ;
        RECT 178.800 132.300 179.600 133.200 ;
        RECT 177.200 131.700 179.600 132.300 ;
        RECT 177.200 131.600 178.000 131.700 ;
        RECT 178.800 131.600 179.600 131.700 ;
        RECT 180.200 130.200 180.800 133.600 ;
        RECT 191.600 132.800 192.400 134.400 ;
        RECT 182.000 132.300 182.800 132.400 ;
        RECT 190.000 132.300 190.800 132.400 ;
        RECT 182.000 132.200 190.800 132.300 ;
        RECT 193.200 132.200 193.800 135.800 ;
        RECT 194.800 135.600 195.600 136.400 ;
        RECT 196.400 135.600 197.200 137.200 ;
        RECT 198.200 134.400 198.800 137.800 ;
        RECT 201.200 136.000 202.000 139.800 ;
        RECT 204.400 136.000 205.200 139.800 ;
        RECT 201.200 135.800 205.200 136.000 ;
        RECT 206.000 135.800 206.800 139.800 ;
        RECT 207.600 135.800 208.400 139.800 ;
        RECT 209.200 136.000 210.000 139.800 ;
        RECT 212.400 136.000 213.200 139.800 ;
        RECT 209.200 135.800 213.200 136.000 ;
        RECT 201.400 135.400 205.000 135.800 ;
        RECT 202.000 134.400 202.800 134.800 ;
        RECT 206.000 134.400 206.600 135.800 ;
        RECT 207.800 134.400 208.400 135.800 ;
        RECT 209.400 135.400 213.000 135.800 ;
        RECT 211.600 134.400 212.400 134.800 ;
        RECT 198.000 133.600 198.800 134.400 ;
        RECT 199.600 134.300 200.400 134.400 ;
        RECT 201.200 134.300 202.800 134.400 ;
        RECT 199.600 133.800 202.800 134.300 ;
        RECT 199.600 133.700 202.000 133.800 ;
        RECT 199.600 133.600 200.400 133.700 ;
        RECT 201.200 133.600 202.000 133.700 ;
        RECT 204.200 133.600 206.800 134.400 ;
        RECT 207.600 133.600 210.200 134.400 ;
        RECT 211.600 133.800 213.200 134.400 ;
        RECT 212.400 133.600 213.200 133.800 ;
        RECT 194.800 132.200 195.600 132.400 ;
        RECT 182.000 131.700 191.600 132.200 ;
        RECT 182.000 131.600 182.800 131.700 ;
        RECT 190.000 131.600 191.600 131.700 ;
        RECT 193.200 131.600 195.600 132.200 ;
        RECT 190.800 131.200 191.600 131.600 ;
        RECT 182.000 130.300 182.800 130.400 ;
        RECT 186.800 130.300 187.600 130.400 ;
        RECT 182.000 130.200 187.600 130.300 ;
        RECT 194.800 130.200 195.400 131.600 ;
        RECT 198.200 130.200 198.800 133.600 ;
        RECT 199.600 130.800 200.400 132.400 ;
        RECT 201.200 132.300 202.000 132.400 ;
        RECT 202.800 132.300 203.600 133.200 ;
        RECT 201.200 131.700 203.600 132.300 ;
        RECT 201.200 131.600 202.000 131.700 ;
        RECT 202.800 131.600 203.600 131.700 ;
        RECT 204.200 130.200 204.800 133.600 ;
        RECT 206.000 132.300 206.800 132.400 ;
        RECT 206.000 131.700 208.300 132.300 ;
        RECT 206.000 131.600 206.800 131.700 ;
        RECT 207.700 130.400 208.300 131.700 ;
        RECT 206.000 130.200 206.800 130.400 ;
        RECT 179.800 129.600 180.800 130.200 ;
        RECT 181.400 129.700 187.600 130.200 ;
        RECT 181.400 129.600 182.800 129.700 ;
        RECT 186.800 129.600 187.600 129.700 ;
        RECT 190.000 129.600 194.000 130.200 ;
        RECT 179.800 122.200 180.600 129.600 ;
        RECT 181.400 128.400 182.000 129.600 ;
        RECT 181.200 127.600 182.000 128.400 ;
        RECT 190.000 122.200 190.800 129.600 ;
        RECT 193.200 122.200 194.000 129.600 ;
        RECT 194.800 122.200 195.600 130.200 ;
        RECT 198.000 129.400 199.800 130.200 ;
        RECT 199.000 128.400 199.800 129.400 ;
        RECT 203.800 129.600 204.800 130.200 ;
        RECT 205.400 129.600 206.800 130.200 ;
        RECT 207.600 130.200 208.400 130.400 ;
        RECT 209.600 130.200 210.200 133.600 ;
        RECT 207.600 129.600 209.000 130.200 ;
        RECT 209.600 129.600 210.600 130.200 ;
        RECT 199.000 127.600 200.400 128.400 ;
        RECT 199.000 122.200 199.800 127.600 ;
        RECT 203.800 124.400 204.600 129.600 ;
        RECT 205.400 128.400 206.000 129.600 ;
        RECT 205.200 127.600 206.000 128.400 ;
        RECT 208.400 128.400 209.000 129.600 ;
        RECT 208.400 127.600 209.200 128.400 ;
        RECT 202.800 123.600 204.600 124.400 ;
        RECT 203.800 122.200 204.600 123.600 ;
        RECT 209.800 122.200 210.600 129.600 ;
        RECT 214.000 122.200 214.800 139.800 ;
        RECT 215.600 135.600 216.400 137.200 ;
        RECT 217.400 136.400 218.200 137.200 ;
        RECT 217.200 135.600 218.000 136.400 ;
        RECT 218.800 135.800 219.600 139.800 ;
        RECT 217.200 132.200 218.000 132.400 ;
        RECT 219.000 132.200 219.600 135.800 ;
        RECT 220.400 132.800 221.200 134.400 ;
        RECT 225.200 134.300 226.000 139.800 ;
        RECT 229.400 136.400 230.200 139.800 ;
        RECT 228.400 135.800 230.200 136.400 ;
        RECT 231.600 136.000 232.400 139.800 ;
        RECT 234.800 136.000 235.600 139.800 ;
        RECT 231.600 135.800 235.600 136.000 ;
        RECT 236.400 135.800 237.200 139.800 ;
        RECT 226.800 134.300 227.600 135.200 ;
        RECT 225.200 133.700 227.600 134.300 ;
        RECT 222.000 132.200 222.800 132.400 ;
        RECT 217.200 131.600 219.600 132.200 ;
        RECT 221.200 131.600 222.800 132.200 ;
        RECT 217.400 130.200 218.000 131.600 ;
        RECT 221.200 131.200 222.000 131.600 ;
        RECT 217.200 122.200 218.000 130.200 ;
        RECT 218.800 129.600 222.800 130.200 ;
        RECT 218.800 122.200 219.600 129.600 ;
        RECT 222.000 122.200 222.800 129.600 ;
        RECT 225.200 122.200 226.000 133.700 ;
        RECT 226.800 133.600 227.600 133.700 ;
        RECT 226.800 132.300 227.600 132.400 ;
        RECT 228.400 132.300 229.200 135.800 ;
        RECT 231.800 135.400 235.400 135.800 ;
        RECT 232.400 134.400 233.200 134.800 ;
        RECT 236.400 134.400 237.000 135.800 ;
        RECT 231.600 133.800 233.200 134.400 ;
        RECT 231.600 133.600 232.400 133.800 ;
        RECT 234.600 133.600 237.200 134.400 ;
        RECT 233.200 132.300 234.000 133.200 ;
        RECT 226.800 131.700 229.200 132.300 ;
        RECT 226.800 131.600 227.600 131.700 ;
        RECT 228.400 122.200 229.200 131.700 ;
        RECT 230.100 131.700 234.000 132.300 ;
        RECT 230.100 130.400 230.700 131.700 ;
        RECT 233.200 131.600 234.000 131.700 ;
        RECT 230.000 128.800 230.800 130.400 ;
        RECT 234.600 130.200 235.200 133.600 ;
        RECT 238.000 132.300 238.800 132.400 ;
        RECT 239.600 132.300 240.400 139.800 ;
        RECT 241.200 135.600 242.000 137.200 ;
        RECT 238.000 131.700 240.400 132.300 ;
        RECT 238.000 131.600 238.800 131.700 ;
        RECT 236.400 130.200 237.200 130.400 ;
        RECT 234.200 129.600 235.200 130.200 ;
        RECT 235.800 129.600 237.200 130.200 ;
        RECT 234.200 122.200 235.000 129.600 ;
        RECT 235.800 128.400 236.400 129.600 ;
        RECT 235.600 127.600 236.400 128.400 ;
        RECT 239.600 122.200 240.400 131.700 ;
        RECT 242.800 122.200 243.600 139.800 ;
        RECT 248.000 134.200 248.800 139.800 ;
        RECT 248.000 133.800 249.800 134.200 ;
        RECT 248.200 133.600 249.800 133.800 ;
        RECT 246.000 131.600 247.600 132.400 ;
        RECT 244.400 129.600 245.200 131.200 ;
        RECT 249.200 130.400 249.800 133.600 ;
        RECT 249.200 129.600 250.000 130.400 ;
        RECT 247.600 127.600 248.400 129.200 ;
        RECT 249.200 127.000 249.800 129.600 ;
        RECT 246.200 126.400 249.800 127.000 ;
        RECT 246.200 126.200 246.800 126.400 ;
        RECT 246.000 122.200 246.800 126.200 ;
        RECT 249.200 126.200 249.800 126.400 ;
        RECT 249.200 122.200 250.000 126.200 ;
        RECT 4.400 112.400 5.200 119.800 ;
        RECT 3.000 111.800 5.200 112.400 ;
        RECT 7.600 112.000 8.400 119.800 ;
        RECT 10.800 115.200 11.600 119.800 ;
        RECT 3.000 111.200 3.600 111.800 ;
        RECT 2.400 110.400 3.600 111.200 ;
        RECT 7.400 111.200 8.400 112.000 ;
        RECT 9.000 114.600 11.600 115.200 ;
        RECT 9.000 113.000 9.600 114.600 ;
        RECT 14.000 114.400 14.800 119.800 ;
        RECT 17.200 117.000 18.000 119.800 ;
        RECT 18.800 117.000 19.600 119.800 ;
        RECT 20.400 117.000 21.200 119.800 ;
        RECT 15.400 114.400 19.600 115.200 ;
        RECT 12.200 113.600 14.800 114.400 ;
        RECT 22.000 113.600 22.800 119.800 ;
        RECT 25.200 115.000 26.000 119.800 ;
        RECT 28.400 115.000 29.200 119.800 ;
        RECT 30.000 117.000 30.800 119.800 ;
        RECT 31.600 117.000 32.400 119.800 ;
        RECT 34.800 115.200 35.600 119.800 ;
        RECT 38.000 116.400 38.800 119.800 ;
        RECT 38.000 115.800 39.000 116.400 ;
        RECT 38.400 115.200 39.000 115.800 ;
        RECT 33.600 114.400 37.800 115.200 ;
        RECT 38.400 114.600 40.400 115.200 ;
        RECT 25.200 113.600 27.800 114.400 ;
        RECT 28.400 113.800 34.200 114.400 ;
        RECT 37.200 114.000 37.800 114.400 ;
        RECT 17.200 113.000 18.000 113.200 ;
        RECT 9.000 112.400 18.000 113.000 ;
        RECT 20.400 113.000 21.200 113.200 ;
        RECT 28.400 113.000 29.000 113.800 ;
        RECT 34.800 113.200 36.200 113.800 ;
        RECT 37.200 113.200 38.800 114.000 ;
        RECT 20.400 112.400 29.000 113.000 ;
        RECT 30.000 113.000 36.200 113.200 ;
        RECT 30.000 112.600 35.400 113.000 ;
        RECT 30.000 112.400 30.800 112.600 ;
        RECT 3.000 107.400 3.600 110.400 ;
        RECT 4.400 110.300 5.200 110.400 ;
        RECT 7.400 110.300 8.200 111.200 ;
        RECT 9.000 110.600 9.600 112.400 ;
        RECT 4.400 109.700 8.200 110.300 ;
        RECT 4.400 108.800 5.200 109.700 ;
        RECT 3.000 106.800 5.200 107.400 ;
        RECT 4.400 102.200 5.200 106.800 ;
        RECT 7.400 106.800 8.200 109.700 ;
        RECT 8.800 110.000 9.600 110.600 ;
        RECT 15.600 110.000 39.000 110.600 ;
        RECT 8.800 108.000 9.400 110.000 ;
        RECT 15.600 109.400 16.400 110.000 ;
        RECT 33.200 109.600 34.000 110.000 ;
        RECT 34.800 109.600 35.600 110.000 ;
        RECT 36.400 109.600 37.200 110.000 ;
        RECT 38.200 109.800 39.000 110.000 ;
        RECT 10.000 108.600 13.800 109.400 ;
        RECT 8.800 107.400 10.000 108.000 ;
        RECT 7.400 106.000 8.400 106.800 ;
        RECT 7.600 102.200 8.400 106.000 ;
        RECT 9.200 102.200 10.000 107.400 ;
        RECT 13.000 107.400 13.800 108.600 ;
        RECT 13.000 106.800 14.800 107.400 ;
        RECT 14.000 106.200 14.800 106.800 ;
        RECT 18.800 106.400 19.600 109.200 ;
        RECT 22.000 108.600 25.200 109.400 ;
        RECT 29.000 108.600 31.000 109.400 ;
        RECT 39.600 109.000 40.400 114.600 ;
        RECT 41.200 112.400 42.000 119.800 ;
        RECT 44.400 112.400 45.200 119.800 ;
        RECT 41.200 111.800 45.200 112.400 ;
        RECT 46.000 111.800 46.800 119.800 ;
        RECT 50.200 112.600 51.000 119.800 ;
        RECT 49.200 111.800 51.000 112.600 ;
        RECT 55.000 112.400 55.800 119.800 ;
        RECT 60.400 115.800 61.200 119.800 ;
        RECT 56.400 113.600 57.200 114.400 ;
        RECT 56.600 112.400 57.200 113.600 ;
        RECT 55.000 111.800 56.000 112.400 ;
        RECT 56.600 111.800 58.000 112.400 ;
        RECT 42.000 110.400 42.800 110.800 ;
        RECT 46.000 110.400 46.600 111.800 ;
        RECT 41.200 109.800 42.800 110.400 ;
        RECT 44.400 109.800 46.800 110.400 ;
        RECT 41.200 109.600 42.000 109.800 ;
        RECT 21.600 107.800 22.400 108.000 ;
        RECT 21.600 107.200 26.000 107.800 ;
        RECT 25.200 107.000 26.000 107.200 ;
        RECT 26.800 106.800 27.600 108.400 ;
        RECT 14.000 105.400 16.400 106.200 ;
        RECT 18.800 105.600 19.800 106.400 ;
        RECT 22.800 105.600 24.400 106.400 ;
        RECT 25.200 106.200 26.000 106.400 ;
        RECT 29.000 106.200 29.800 108.600 ;
        RECT 31.600 108.200 40.400 109.000 ;
        RECT 35.000 106.800 38.000 107.600 ;
        RECT 35.000 106.200 35.800 106.800 ;
        RECT 25.200 105.600 29.800 106.200 ;
        RECT 15.600 102.200 16.400 105.400 ;
        RECT 33.200 105.400 35.800 106.200 ;
        RECT 17.200 102.200 18.000 105.000 ;
        RECT 18.800 102.200 19.600 105.000 ;
        RECT 20.400 102.200 21.200 105.000 ;
        RECT 22.000 102.200 22.800 105.000 ;
        RECT 25.200 102.200 26.000 105.000 ;
        RECT 28.400 102.200 29.200 105.000 ;
        RECT 30.000 102.200 30.800 105.000 ;
        RECT 31.600 102.200 32.400 105.000 ;
        RECT 33.200 102.200 34.000 105.400 ;
        RECT 39.600 102.200 40.400 108.200 ;
        RECT 42.800 107.600 43.600 109.200 ;
        RECT 44.400 106.200 45.000 109.800 ;
        RECT 46.000 109.600 46.800 109.800 ;
        RECT 49.400 108.400 50.000 111.800 ;
        RECT 50.800 109.600 51.600 111.200 ;
        RECT 55.400 110.400 56.000 111.800 ;
        RECT 57.200 111.600 58.000 111.800 ;
        RECT 60.600 111.600 61.200 115.800 ;
        RECT 63.600 111.800 64.400 119.800 ;
        RECT 74.800 112.400 75.600 119.800 ;
        RECT 60.600 111.000 63.000 111.600 ;
        RECT 54.000 108.800 54.800 110.400 ;
        RECT 55.400 109.600 56.400 110.400 ;
        RECT 60.400 109.600 61.200 110.400 ;
        RECT 55.400 108.400 56.000 109.600 ;
        RECT 49.200 108.300 50.000 108.400 ;
        RECT 46.100 107.700 50.000 108.300 ;
        RECT 46.100 106.400 46.700 107.700 ;
        RECT 49.200 107.600 50.000 107.700 ;
        RECT 52.400 108.200 53.200 108.400 ;
        RECT 52.400 107.600 54.000 108.200 ;
        RECT 55.400 107.600 58.000 108.400 ;
        RECT 58.800 107.600 59.600 109.200 ;
        RECT 60.600 108.800 61.200 109.600 ;
        RECT 60.600 108.200 61.600 108.800 ;
        RECT 60.800 108.000 61.600 108.200 ;
        RECT 62.400 107.600 63.000 111.000 ;
        RECT 63.800 110.400 64.400 111.800 ;
        RECT 73.400 111.800 75.600 112.400 ;
        RECT 76.400 112.400 77.200 119.800 ;
        RECT 78.000 112.400 78.800 112.600 ;
        RECT 80.800 112.400 82.400 119.800 ;
        RECT 76.400 111.800 78.800 112.400 ;
        RECT 79.600 111.800 82.400 112.400 ;
        RECT 84.600 112.400 85.400 112.600 ;
        RECT 86.000 112.400 86.800 119.800 ;
        RECT 84.600 111.800 86.800 112.400 ;
        RECT 90.200 111.800 92.200 119.800 ;
        RECT 97.200 116.400 98.000 119.800 ;
        RECT 97.000 115.800 98.000 116.400 ;
        RECT 97.000 115.200 97.600 115.800 ;
        RECT 100.400 115.200 101.200 119.800 ;
        RECT 103.600 117.000 104.400 119.800 ;
        RECT 105.200 117.000 106.000 119.800 ;
        RECT 95.600 114.600 97.600 115.200 ;
        RECT 73.400 111.200 74.000 111.800 ;
        RECT 79.600 111.600 81.000 111.800 ;
        RECT 72.800 110.400 74.000 111.200 ;
        RECT 80.400 110.400 81.000 111.600 ;
        RECT 84.600 111.200 85.200 111.800 ;
        RECT 81.800 110.600 85.200 111.200 ;
        RECT 81.800 110.400 82.600 110.600 ;
        RECT 63.600 109.600 64.400 110.400 ;
        RECT 44.400 102.200 45.200 106.200 ;
        RECT 46.000 105.600 46.800 106.400 ;
        RECT 45.800 104.800 46.600 105.600 ;
        RECT 47.600 104.800 48.400 106.400 ;
        RECT 49.400 104.200 50.000 107.600 ;
        RECT 53.200 107.200 54.000 107.600 ;
        RECT 52.600 106.200 56.200 106.600 ;
        RECT 57.200 106.200 57.800 107.600 ;
        RECT 62.400 107.400 63.200 107.600 ;
        RECT 60.200 107.000 63.200 107.400 ;
        RECT 59.000 106.800 63.200 107.000 ;
        RECT 59.000 106.400 60.800 106.800 ;
        RECT 59.000 106.200 59.600 106.400 ;
        RECT 63.800 106.200 64.400 109.600 ;
        RECT 73.400 107.400 74.000 110.400 ;
        RECT 74.800 110.300 75.600 110.400 ;
        RECT 74.800 109.700 77.100 110.300 ;
        RECT 74.800 108.800 75.600 109.700 ;
        RECT 76.500 108.400 77.100 109.700 ;
        RECT 79.600 109.800 81.000 110.400 ;
        RECT 84.000 109.800 84.800 110.000 ;
        RECT 79.600 109.600 81.400 109.800 ;
        RECT 80.400 109.200 81.400 109.600 ;
        RECT 76.400 107.600 78.000 108.400 ;
        RECT 79.200 107.600 80.000 108.400 ;
        RECT 73.400 106.800 75.600 107.400 ;
        RECT 79.400 107.200 80.000 107.600 ;
        RECT 78.000 106.800 78.800 107.000 ;
        RECT 49.200 102.200 50.000 104.200 ;
        RECT 52.400 106.000 56.400 106.200 ;
        RECT 52.400 102.200 53.200 106.000 ;
        RECT 55.600 102.200 56.400 106.000 ;
        RECT 57.200 102.200 58.000 106.200 ;
        RECT 58.800 102.200 59.600 106.200 ;
        RECT 63.000 105.200 64.400 106.200 ;
        RECT 63.000 102.200 63.800 105.200 ;
        RECT 74.800 102.200 75.600 106.800 ;
        RECT 76.400 106.200 78.800 106.800 ;
        RECT 79.400 106.400 80.200 107.200 ;
        RECT 76.400 102.200 77.200 106.200 ;
        RECT 80.800 105.800 81.400 109.200 ;
        RECT 82.200 109.200 84.800 109.800 ;
        RECT 82.200 108.600 82.800 109.200 ;
        RECT 82.000 107.800 82.800 108.600 ;
        RECT 85.200 108.200 86.800 108.400 ;
        RECT 83.400 107.600 86.800 108.200 ;
        RECT 87.600 107.600 88.400 109.200 ;
        RECT 89.200 108.800 90.000 110.400 ;
        RECT 91.000 108.400 91.600 111.800 ;
        RECT 92.400 108.800 93.200 110.400 ;
        RECT 95.600 109.000 96.400 114.600 ;
        RECT 98.200 114.400 102.400 115.200 ;
        RECT 106.800 115.000 107.600 119.800 ;
        RECT 110.000 115.000 110.800 119.800 ;
        RECT 98.200 114.000 98.800 114.400 ;
        RECT 97.200 113.200 98.800 114.000 ;
        RECT 101.800 113.800 107.600 114.400 ;
        RECT 99.800 113.200 101.200 113.800 ;
        RECT 99.800 113.000 106.000 113.200 ;
        RECT 100.600 112.600 106.000 113.000 ;
        RECT 105.200 112.400 106.000 112.600 ;
        RECT 107.000 113.000 107.600 113.800 ;
        RECT 108.200 113.600 110.800 114.400 ;
        RECT 113.200 113.600 114.000 119.800 ;
        RECT 114.800 117.000 115.600 119.800 ;
        RECT 116.400 117.000 117.200 119.800 ;
        RECT 118.000 117.000 118.800 119.800 ;
        RECT 116.400 114.400 120.600 115.200 ;
        RECT 121.200 114.400 122.000 119.800 ;
        RECT 124.400 115.200 125.200 119.800 ;
        RECT 124.400 114.600 127.000 115.200 ;
        RECT 121.200 113.600 123.800 114.400 ;
        RECT 114.800 113.000 115.600 113.200 ;
        RECT 107.000 112.400 115.600 113.000 ;
        RECT 118.000 113.000 118.800 113.200 ;
        RECT 126.400 113.000 127.000 114.600 ;
        RECT 118.000 112.400 127.000 113.000 ;
        RECT 126.400 110.600 127.000 112.400 ;
        RECT 127.600 112.000 128.400 119.800 ;
        RECT 127.600 111.200 128.600 112.000 ;
        RECT 97.000 110.000 120.400 110.600 ;
        RECT 126.400 110.000 127.200 110.600 ;
        RECT 97.000 109.800 97.800 110.000 ;
        RECT 102.000 109.600 102.800 110.000 ;
        RECT 108.400 109.600 109.200 110.000 ;
        RECT 119.600 109.400 120.400 110.000 ;
        RECT 90.800 108.200 91.600 108.400 ;
        RECT 94.000 108.200 94.800 108.400 ;
        RECT 89.200 107.600 91.600 108.200 ;
        RECT 93.200 107.600 94.800 108.200 ;
        RECT 95.600 108.200 104.400 109.000 ;
        RECT 105.000 108.600 107.000 109.400 ;
        RECT 110.800 108.600 114.000 109.400 ;
        RECT 83.400 107.200 84.000 107.600 ;
        RECT 82.000 106.600 84.000 107.200 ;
        RECT 84.600 106.800 85.400 107.000 ;
        RECT 82.000 106.400 83.600 106.600 ;
        RECT 84.600 106.200 86.800 106.800 ;
        RECT 89.200 106.200 89.800 107.600 ;
        RECT 93.200 107.200 94.000 107.600 ;
        RECT 91.000 106.200 94.600 106.600 ;
        RECT 80.800 102.200 82.400 105.800 ;
        RECT 86.000 102.200 86.800 106.200 ;
        RECT 87.600 102.800 88.400 106.200 ;
        RECT 89.200 103.400 90.000 106.200 ;
        RECT 90.800 106.000 94.800 106.200 ;
        RECT 90.800 102.800 91.600 106.000 ;
        RECT 87.600 102.200 91.600 102.800 ;
        RECT 94.000 102.200 94.800 106.000 ;
        RECT 95.600 102.200 96.400 108.200 ;
        RECT 98.000 106.800 101.000 107.600 ;
        RECT 100.200 106.200 101.000 106.800 ;
        RECT 106.200 106.200 107.000 108.600 ;
        RECT 108.400 106.800 109.200 108.400 ;
        RECT 113.600 107.800 114.400 108.000 ;
        RECT 110.000 107.200 114.400 107.800 ;
        RECT 110.000 107.000 110.800 107.200 ;
        RECT 116.400 106.400 117.200 109.200 ;
        RECT 122.200 108.600 126.000 109.400 ;
        RECT 122.200 107.400 123.000 108.600 ;
        RECT 126.600 108.000 127.200 110.000 ;
        RECT 110.000 106.200 110.800 106.400 ;
        RECT 100.200 105.400 102.800 106.200 ;
        RECT 106.200 105.600 110.800 106.200 ;
        RECT 111.600 105.600 113.200 106.400 ;
        RECT 116.200 105.600 117.200 106.400 ;
        RECT 121.200 106.800 123.000 107.400 ;
        RECT 126.000 107.400 127.200 108.000 ;
        RECT 121.200 106.200 122.000 106.800 ;
        RECT 102.000 102.200 102.800 105.400 ;
        RECT 119.600 105.400 122.000 106.200 ;
        RECT 103.600 102.200 104.400 105.000 ;
        RECT 105.200 102.200 106.000 105.000 ;
        RECT 106.800 102.200 107.600 105.000 ;
        RECT 110.000 102.200 110.800 105.000 ;
        RECT 113.200 102.200 114.000 105.000 ;
        RECT 114.800 102.200 115.600 105.000 ;
        RECT 116.400 102.200 117.200 105.000 ;
        RECT 118.000 102.200 118.800 105.000 ;
        RECT 119.600 102.200 120.400 105.400 ;
        RECT 126.000 102.200 126.800 107.400 ;
        RECT 127.800 106.800 128.600 111.200 ;
        RECT 127.600 106.000 128.600 106.800 ;
        RECT 130.800 111.800 131.600 119.800 ;
        RECT 134.000 115.800 134.800 119.800 ;
        RECT 130.800 110.400 131.400 111.800 ;
        RECT 134.000 111.600 134.600 115.800 ;
        RECT 138.000 113.600 138.800 114.400 ;
        RECT 138.000 112.400 138.600 113.600 ;
        RECT 139.400 112.400 140.200 119.800 ;
        RECT 135.600 112.300 136.400 112.400 ;
        RECT 137.200 112.300 138.600 112.400 ;
        RECT 135.600 111.800 138.600 112.300 ;
        RECT 139.200 111.800 140.200 112.400 ;
        RECT 146.200 112.400 147.000 119.800 ;
        RECT 147.600 113.600 148.400 114.400 ;
        RECT 147.800 112.400 148.400 113.600 ;
        RECT 146.200 111.800 147.200 112.400 ;
        RECT 147.800 111.800 149.200 112.400 ;
        RECT 152.600 111.800 154.600 119.800 ;
        RECT 158.000 111.800 158.800 119.800 ;
        RECT 159.600 112.400 160.400 119.800 ;
        RECT 162.800 112.400 163.600 119.800 ;
        RECT 165.200 113.600 166.000 114.400 ;
        RECT 165.200 112.400 165.800 113.600 ;
        RECT 166.600 112.400 167.400 119.800 ;
        RECT 173.400 114.300 174.200 119.800 ;
        RECT 175.600 114.300 176.400 114.400 ;
        RECT 173.400 113.700 176.400 114.300 ;
        RECT 173.400 112.600 174.200 113.700 ;
        RECT 175.600 113.600 176.400 113.700 ;
        RECT 159.600 111.800 163.600 112.400 ;
        RECT 164.400 111.800 165.800 112.400 ;
        RECT 166.400 111.800 167.400 112.400 ;
        RECT 172.400 111.800 174.200 112.600 ;
        RECT 135.600 111.700 138.000 111.800 ;
        RECT 135.600 111.600 136.400 111.700 ;
        RECT 137.200 111.600 138.000 111.700 ;
        RECT 132.200 111.000 134.600 111.600 ;
        RECT 130.800 109.600 131.600 110.400 ;
        RECT 130.800 106.200 131.400 109.600 ;
        RECT 132.200 107.600 132.800 111.000 ;
        RECT 139.200 110.400 139.800 111.800 ;
        RECT 134.000 109.600 134.800 110.400 ;
        RECT 138.800 109.600 139.800 110.400 ;
        RECT 134.000 108.800 134.600 109.600 ;
        RECT 133.600 108.200 134.600 108.800 ;
        RECT 133.600 108.000 134.400 108.200 ;
        RECT 135.600 107.600 136.400 109.200 ;
        RECT 139.200 108.400 139.800 109.600 ;
        RECT 140.400 108.800 141.200 110.400 ;
        RECT 145.200 108.800 146.000 110.400 ;
        RECT 146.600 110.300 147.200 111.800 ;
        RECT 148.400 111.600 149.200 111.800 ;
        RECT 148.400 110.300 149.200 110.400 ;
        RECT 146.600 109.700 149.200 110.300 ;
        RECT 146.600 108.400 147.200 109.700 ;
        RECT 148.400 109.600 149.200 109.700 ;
        RECT 137.200 107.600 139.800 108.400 ;
        RECT 142.000 108.200 142.800 108.400 ;
        RECT 141.200 107.600 142.800 108.200 ;
        RECT 143.600 108.200 144.400 108.400 ;
        RECT 143.600 107.600 145.200 108.200 ;
        RECT 146.600 107.600 149.200 108.400 ;
        RECT 150.000 107.600 150.800 109.200 ;
        RECT 151.600 108.800 152.400 110.400 ;
        RECT 153.400 108.400 154.000 111.800 ;
        RECT 158.200 110.400 158.800 111.800 ;
        RECT 164.400 111.600 165.200 111.800 ;
        RECT 162.000 110.400 162.800 110.800 ;
        RECT 166.400 110.400 167.000 111.800 ;
        RECT 154.800 108.800 155.600 110.400 ;
        RECT 158.000 109.800 160.400 110.400 ;
        RECT 162.000 109.800 163.600 110.400 ;
        RECT 158.000 109.600 158.800 109.800 ;
        RECT 153.200 108.200 154.000 108.400 ;
        RECT 156.400 108.200 157.200 108.400 ;
        RECT 151.600 107.600 154.000 108.200 ;
        RECT 155.600 107.600 157.200 108.200 ;
        RECT 132.000 107.400 132.800 107.600 ;
        RECT 132.000 107.000 135.000 107.400 ;
        RECT 132.000 106.800 136.200 107.000 ;
        RECT 134.400 106.400 136.200 106.800 ;
        RECT 135.600 106.200 136.200 106.400 ;
        RECT 137.400 106.200 138.000 107.600 ;
        RECT 141.200 107.200 142.000 107.600 ;
        RECT 144.400 107.200 145.200 107.600 ;
        RECT 139.000 106.200 142.600 106.600 ;
        RECT 143.800 106.200 147.400 106.600 ;
        RECT 148.400 106.200 149.000 107.600 ;
        RECT 151.600 106.200 152.200 107.600 ;
        RECT 155.600 107.200 156.400 107.600 ;
        RECT 153.400 106.200 157.000 106.600 ;
        RECT 127.600 102.200 128.400 106.000 ;
        RECT 130.800 105.200 132.200 106.200 ;
        RECT 131.400 102.200 132.200 105.200 ;
        RECT 135.600 102.200 136.400 106.200 ;
        RECT 137.200 102.200 138.000 106.200 ;
        RECT 138.800 106.000 142.800 106.200 ;
        RECT 138.800 102.200 139.600 106.000 ;
        RECT 142.000 102.200 142.800 106.000 ;
        RECT 143.600 106.000 147.600 106.200 ;
        RECT 143.600 102.200 144.400 106.000 ;
        RECT 146.800 102.200 147.600 106.000 ;
        RECT 148.400 102.200 149.200 106.200 ;
        RECT 150.000 102.800 150.800 106.200 ;
        RECT 151.600 103.400 152.400 106.200 ;
        RECT 153.200 106.000 157.200 106.200 ;
        RECT 153.200 102.800 154.000 106.000 ;
        RECT 150.000 102.200 154.000 102.800 ;
        RECT 156.400 102.200 157.200 106.000 ;
        RECT 158.000 105.600 158.800 106.400 ;
        RECT 159.800 106.200 160.400 109.800 ;
        RECT 162.800 109.600 163.600 109.800 ;
        RECT 166.000 109.600 167.000 110.400 ;
        RECT 161.200 107.600 162.000 109.200 ;
        RECT 166.400 108.400 167.000 109.600 ;
        RECT 167.600 108.800 168.400 110.400 ;
        RECT 172.600 108.400 173.200 111.800 ;
        RECT 174.000 109.600 174.800 111.200 ;
        RECT 177.200 110.300 178.000 119.800 ;
        RECT 179.400 118.400 180.200 119.800 ;
        RECT 178.800 117.600 180.200 118.400 ;
        RECT 179.400 112.600 180.200 117.600 ;
        RECT 179.400 111.800 181.200 112.600 ;
        RECT 190.000 112.400 190.800 119.800 ;
        RECT 193.200 119.200 197.200 119.800 ;
        RECT 193.200 112.400 194.000 119.200 ;
        RECT 190.000 111.800 194.000 112.400 ;
        RECT 194.800 111.800 195.600 118.600 ;
        RECT 196.400 111.800 197.200 119.200 ;
        RECT 200.600 112.600 201.400 119.800 ;
        RECT 199.600 111.800 201.400 112.600 ;
        RECT 203.600 113.600 204.400 114.400 ;
        RECT 203.600 112.400 204.200 113.600 ;
        RECT 205.000 112.400 205.800 119.800 ;
        RECT 210.800 116.400 211.600 119.800 ;
        RECT 210.600 115.800 211.600 116.400 ;
        RECT 210.600 115.200 211.200 115.800 ;
        RECT 214.000 115.200 214.800 119.800 ;
        RECT 217.200 117.000 218.000 119.800 ;
        RECT 218.800 117.000 219.600 119.800 ;
        RECT 202.800 111.800 204.200 112.400 ;
        RECT 204.800 111.800 205.800 112.400 ;
        RECT 209.200 114.600 211.200 115.200 ;
        RECT 178.800 110.300 179.600 111.200 ;
        RECT 177.200 109.700 179.600 110.300 ;
        RECT 164.400 107.600 167.000 108.400 ;
        RECT 169.200 108.200 170.000 108.400 ;
        RECT 168.400 107.600 170.000 108.200 ;
        RECT 172.400 107.600 173.200 108.400 ;
        RECT 164.600 106.200 165.200 107.600 ;
        RECT 168.400 107.200 169.200 107.600 ;
        RECT 166.200 106.200 169.800 106.600 ;
        RECT 158.200 104.800 159.000 105.600 ;
        RECT 159.600 102.200 160.400 106.200 ;
        RECT 164.400 102.200 165.200 106.200 ;
        RECT 166.000 106.000 170.000 106.200 ;
        RECT 166.000 102.200 166.800 106.000 ;
        RECT 169.200 102.200 170.000 106.000 ;
        RECT 170.800 104.800 171.600 106.400 ;
        RECT 172.600 104.200 173.200 107.600 ;
        RECT 177.200 108.300 178.000 109.700 ;
        RECT 178.800 109.600 179.600 109.700 ;
        RECT 180.400 108.400 181.000 111.800 ;
        RECT 194.800 111.200 195.400 111.800 ;
        RECT 190.800 110.400 191.600 110.800 ;
        RECT 193.400 110.600 195.400 111.200 ;
        RECT 193.400 110.400 194.000 110.600 ;
        RECT 190.000 109.800 191.600 110.400 ;
        RECT 190.000 109.600 190.800 109.800 ;
        RECT 193.200 109.600 194.000 110.400 ;
        RECT 196.400 109.600 197.200 111.200 ;
        RECT 178.800 108.300 179.600 108.400 ;
        RECT 177.200 107.700 179.600 108.300 ;
        RECT 175.600 104.800 176.400 106.400 ;
        RECT 172.400 102.200 173.200 104.200 ;
        RECT 177.200 102.200 178.000 107.700 ;
        RECT 178.800 107.600 179.600 107.700 ;
        RECT 180.400 107.600 181.200 108.400 ;
        RECT 183.600 108.300 184.400 108.400 ;
        RECT 191.600 108.300 192.400 109.200 ;
        RECT 183.600 107.700 192.400 108.300 ;
        RECT 183.600 107.600 184.400 107.700 ;
        RECT 191.600 107.600 192.400 107.700 ;
        RECT 180.400 104.200 181.000 107.600 ;
        RECT 182.000 104.800 182.800 106.400 ;
        RECT 193.400 106.200 194.000 109.600 ;
        RECT 194.600 108.800 195.400 109.600 ;
        RECT 194.800 108.400 195.400 108.800 ;
        RECT 199.800 108.400 200.400 111.800 ;
        RECT 202.800 111.600 203.600 111.800 ;
        RECT 201.200 109.600 202.000 111.200 ;
        RECT 204.800 108.400 205.400 111.800 ;
        RECT 206.000 108.800 206.800 110.400 ;
        RECT 209.200 109.000 210.000 114.600 ;
        RECT 211.800 114.400 216.000 115.200 ;
        RECT 220.400 115.000 221.200 119.800 ;
        RECT 223.600 115.000 224.400 119.800 ;
        RECT 211.800 114.000 212.400 114.400 ;
        RECT 210.800 113.200 212.400 114.000 ;
        RECT 215.400 113.800 221.200 114.400 ;
        RECT 213.400 113.200 214.800 113.800 ;
        RECT 213.400 113.000 219.600 113.200 ;
        RECT 214.200 112.600 219.600 113.000 ;
        RECT 218.800 112.400 219.600 112.600 ;
        RECT 220.600 113.000 221.200 113.800 ;
        RECT 221.800 113.600 224.400 114.400 ;
        RECT 226.800 113.600 227.600 119.800 ;
        RECT 228.400 117.000 229.200 119.800 ;
        RECT 230.000 117.000 230.800 119.800 ;
        RECT 231.600 117.000 232.400 119.800 ;
        RECT 230.000 114.400 234.200 115.200 ;
        RECT 234.800 114.400 235.600 119.800 ;
        RECT 238.000 115.200 238.800 119.800 ;
        RECT 238.000 114.600 240.600 115.200 ;
        RECT 234.800 113.600 237.400 114.400 ;
        RECT 228.400 113.000 229.200 113.200 ;
        RECT 220.600 112.400 229.200 113.000 ;
        RECT 231.600 113.000 232.400 113.200 ;
        RECT 240.000 113.000 240.600 114.600 ;
        RECT 231.600 112.400 240.600 113.000 ;
        RECT 240.000 110.600 240.600 112.400 ;
        RECT 241.200 112.000 242.000 119.800 ;
        RECT 247.000 112.400 247.800 119.800 ;
        RECT 241.200 111.200 242.200 112.000 ;
        RECT 247.000 111.800 248.000 112.400 ;
        RECT 210.600 110.000 234.000 110.600 ;
        RECT 240.000 110.000 240.800 110.600 ;
        RECT 210.600 109.800 211.400 110.000 ;
        RECT 212.400 109.600 213.200 110.000 ;
        RECT 215.600 109.600 216.400 110.000 ;
        RECT 233.200 109.400 234.000 110.000 ;
        RECT 194.800 108.300 195.600 108.400 ;
        RECT 199.600 108.300 200.400 108.400 ;
        RECT 194.800 107.700 200.400 108.300 ;
        RECT 194.800 107.600 195.600 107.700 ;
        RECT 199.600 107.600 200.400 107.700 ;
        RECT 202.800 107.600 205.400 108.400 ;
        RECT 207.600 108.200 208.400 108.400 ;
        RECT 206.800 107.600 208.400 108.200 ;
        RECT 209.200 108.200 218.000 109.000 ;
        RECT 218.600 108.600 220.600 109.400 ;
        RECT 224.400 108.600 227.600 109.400 ;
        RECT 193.000 104.400 194.600 106.200 ;
        RECT 198.000 104.800 198.800 106.400 ;
        RECT 180.400 102.200 181.200 104.200 ;
        RECT 193.000 103.600 195.600 104.400 ;
        RECT 199.800 104.200 200.400 107.600 ;
        RECT 203.000 106.200 203.600 107.600 ;
        RECT 206.800 107.200 207.600 107.600 ;
        RECT 204.600 106.200 208.200 106.600 ;
        RECT 193.000 102.200 194.600 103.600 ;
        RECT 199.600 102.200 200.400 104.200 ;
        RECT 202.800 102.200 203.600 106.200 ;
        RECT 204.400 106.000 208.400 106.200 ;
        RECT 204.400 102.200 205.200 106.000 ;
        RECT 207.600 102.200 208.400 106.000 ;
        RECT 209.200 102.200 210.000 108.200 ;
        RECT 211.600 106.800 214.600 107.600 ;
        RECT 213.800 106.200 214.600 106.800 ;
        RECT 219.800 106.200 220.600 108.600 ;
        RECT 222.000 106.800 222.800 108.400 ;
        RECT 227.200 107.800 228.000 108.000 ;
        RECT 223.600 107.200 228.000 107.800 ;
        RECT 223.600 107.000 224.400 107.200 ;
        RECT 230.000 106.400 230.800 109.200 ;
        RECT 235.800 108.600 239.600 109.400 ;
        RECT 235.800 107.400 236.600 108.600 ;
        RECT 240.200 108.000 240.800 110.000 ;
        RECT 223.600 106.200 224.400 106.400 ;
        RECT 213.800 105.400 216.400 106.200 ;
        RECT 219.800 105.600 224.400 106.200 ;
        RECT 225.200 105.600 226.800 106.400 ;
        RECT 229.800 105.600 230.800 106.400 ;
        RECT 234.800 106.800 236.600 107.400 ;
        RECT 239.600 107.400 240.800 108.000 ;
        RECT 234.800 106.200 235.600 106.800 ;
        RECT 215.600 102.200 216.400 105.400 ;
        RECT 233.200 105.400 235.600 106.200 ;
        RECT 217.200 102.200 218.000 105.000 ;
        RECT 218.800 102.200 219.600 105.000 ;
        RECT 220.400 102.200 221.200 105.000 ;
        RECT 223.600 102.200 224.400 105.000 ;
        RECT 226.800 102.200 227.600 105.000 ;
        RECT 228.400 102.200 229.200 105.000 ;
        RECT 230.000 102.200 230.800 105.000 ;
        RECT 231.600 102.200 232.400 105.000 ;
        RECT 233.200 102.200 234.000 105.400 ;
        RECT 239.600 102.200 240.400 107.400 ;
        RECT 241.400 106.800 242.200 111.200 ;
        RECT 247.400 110.400 248.000 111.800 ;
        RECT 242.800 110.300 243.600 110.400 ;
        RECT 246.000 110.300 246.800 110.400 ;
        RECT 242.800 109.700 246.800 110.300 ;
        RECT 242.800 109.600 243.600 109.700 ;
        RECT 246.000 108.800 246.800 109.700 ;
        RECT 247.400 109.600 248.400 110.400 ;
        RECT 247.400 108.400 248.000 109.600 ;
        RECT 247.400 107.600 250.000 108.400 ;
        RECT 241.200 106.000 242.200 106.800 ;
        RECT 244.600 106.200 248.200 106.600 ;
        RECT 249.200 106.200 249.800 107.600 ;
        RECT 244.400 106.000 248.400 106.200 ;
        RECT 241.200 102.200 242.000 106.000 ;
        RECT 244.400 102.200 245.200 106.000 ;
        RECT 247.600 102.200 248.400 106.000 ;
        RECT 249.200 102.200 250.000 106.200 ;
        RECT 4.400 95.200 5.200 99.800 ;
        RECT 7.600 96.000 8.400 99.800 ;
        RECT 3.000 94.600 5.200 95.200 ;
        RECT 7.400 95.200 8.400 96.000 ;
        RECT 3.000 91.600 3.600 94.600 ;
        RECT 4.400 92.300 5.200 93.200 ;
        RECT 7.400 92.300 8.200 95.200 ;
        RECT 9.200 94.600 10.000 99.800 ;
        RECT 15.600 96.600 16.400 99.800 ;
        RECT 17.200 97.000 18.000 99.800 ;
        RECT 18.800 97.000 19.600 99.800 ;
        RECT 20.400 97.000 21.200 99.800 ;
        RECT 22.000 97.000 22.800 99.800 ;
        RECT 25.200 97.000 26.000 99.800 ;
        RECT 28.400 97.000 29.200 99.800 ;
        RECT 30.000 97.000 30.800 99.800 ;
        RECT 31.600 97.000 32.400 99.800 ;
        RECT 14.000 95.800 16.400 96.600 ;
        RECT 33.200 96.600 34.000 99.800 ;
        RECT 14.000 95.200 14.800 95.800 ;
        RECT 4.400 91.700 8.200 92.300 ;
        RECT 4.400 91.600 5.200 91.700 ;
        RECT 2.400 90.800 3.600 91.600 ;
        RECT 3.000 90.200 3.600 90.800 ;
        RECT 7.400 90.800 8.200 91.700 ;
        RECT 8.800 94.000 10.000 94.600 ;
        RECT 13.000 94.600 14.800 95.200 ;
        RECT 18.800 95.600 19.800 96.400 ;
        RECT 22.800 95.600 24.400 96.400 ;
        RECT 25.200 95.800 29.800 96.400 ;
        RECT 33.200 95.800 35.800 96.600 ;
        RECT 25.200 95.600 26.000 95.800 ;
        RECT 8.800 92.000 9.400 94.000 ;
        RECT 13.000 93.400 13.800 94.600 ;
        RECT 10.000 92.600 13.800 93.400 ;
        RECT 18.800 92.800 19.600 95.600 ;
        RECT 25.200 94.800 26.000 95.000 ;
        RECT 21.600 94.200 26.000 94.800 ;
        RECT 21.600 94.000 22.400 94.200 ;
        RECT 26.800 93.600 27.600 95.200 ;
        RECT 29.000 93.400 29.800 95.800 ;
        RECT 35.000 95.200 35.800 95.800 ;
        RECT 35.000 94.400 38.000 95.200 ;
        RECT 39.600 93.800 40.400 99.800 ;
        RECT 41.200 99.200 45.200 99.800 ;
        RECT 41.200 95.800 42.000 99.200 ;
        RECT 42.800 95.600 43.600 98.600 ;
        RECT 44.400 96.000 45.200 99.200 ;
        RECT 47.600 96.000 48.400 99.800 ;
        RECT 44.400 95.800 48.400 96.000 ;
        RECT 49.200 95.800 50.000 99.800 ;
        RECT 53.600 96.200 55.200 99.800 ;
        RECT 42.800 94.400 43.400 95.600 ;
        RECT 44.600 95.400 48.200 95.800 ;
        RECT 49.200 95.200 51.600 95.800 ;
        RECT 50.800 95.000 51.600 95.200 ;
        RECT 52.200 94.800 53.000 95.600 ;
        RECT 46.800 94.400 47.600 94.800 ;
        RECT 52.200 94.400 52.800 94.800 ;
        RECT 22.000 92.600 25.200 93.400 ;
        RECT 29.000 92.600 31.000 93.400 ;
        RECT 31.600 93.000 40.400 93.800 ;
        RECT 15.600 92.000 16.400 92.600 ;
        RECT 33.200 92.000 34.000 92.400 ;
        RECT 36.400 92.000 37.200 92.400 ;
        RECT 38.200 92.000 39.000 92.200 ;
        RECT 8.800 91.400 9.600 92.000 ;
        RECT 15.600 91.400 39.000 92.000 ;
        RECT 3.000 89.600 5.200 90.200 ;
        RECT 7.400 90.000 8.400 90.800 ;
        RECT 4.400 82.200 5.200 89.600 ;
        RECT 7.600 82.200 8.400 90.000 ;
        RECT 9.000 89.600 9.600 91.400 ;
        RECT 9.000 89.000 18.000 89.600 ;
        RECT 9.000 87.400 9.600 89.000 ;
        RECT 17.200 88.800 18.000 89.000 ;
        RECT 20.400 89.000 29.000 89.600 ;
        RECT 20.400 88.800 21.200 89.000 ;
        RECT 12.200 87.600 14.800 88.400 ;
        RECT 9.000 86.800 11.600 87.400 ;
        RECT 10.800 82.200 11.600 86.800 ;
        RECT 14.000 82.200 14.800 87.600 ;
        RECT 15.400 86.800 19.600 87.600 ;
        RECT 17.200 82.200 18.000 85.000 ;
        RECT 18.800 82.200 19.600 85.000 ;
        RECT 20.400 82.200 21.200 85.000 ;
        RECT 22.000 82.200 22.800 88.400 ;
        RECT 25.200 87.600 27.800 88.400 ;
        RECT 28.400 88.200 29.000 89.000 ;
        RECT 30.000 89.400 30.800 89.600 ;
        RECT 30.000 89.000 35.400 89.400 ;
        RECT 30.000 88.800 36.200 89.000 ;
        RECT 34.800 88.200 36.200 88.800 ;
        RECT 28.400 87.600 34.200 88.200 ;
        RECT 37.200 88.000 38.800 88.800 ;
        RECT 37.200 87.600 37.800 88.000 ;
        RECT 25.200 82.200 26.000 87.000 ;
        RECT 28.400 82.200 29.200 87.000 ;
        RECT 33.600 86.800 37.800 87.600 ;
        RECT 39.600 87.400 40.400 93.000 ;
        RECT 41.200 92.800 42.000 94.400 ;
        RECT 42.800 93.800 45.200 94.400 ;
        RECT 46.800 93.800 48.400 94.400 ;
        RECT 44.400 93.600 45.200 93.800 ;
        RECT 47.600 93.600 48.400 93.800 ;
        RECT 49.200 93.600 50.800 94.400 ;
        RECT 52.000 93.600 52.800 94.400 ;
        RECT 53.600 94.200 54.200 96.200 ;
        RECT 58.800 95.800 59.600 99.800 ;
        RECT 54.800 94.800 56.400 95.600 ;
        RECT 57.000 95.200 59.600 95.800 ;
        RECT 60.400 95.600 61.200 97.200 ;
        RECT 57.000 95.000 57.800 95.200 ;
        RECT 58.000 94.300 59.600 94.400 ;
        RECT 60.500 94.300 61.100 95.600 ;
        RECT 58.000 94.200 61.100 94.300 ;
        RECT 53.600 93.600 54.600 94.200 ;
        RECT 57.400 94.000 61.100 94.200 ;
        RECT 42.800 91.600 43.600 93.200 ;
        RECT 44.600 90.200 45.200 93.600 ;
        RECT 46.000 92.300 46.800 93.200 ;
        RECT 54.000 92.400 54.600 93.600 ;
        RECT 55.200 93.700 61.100 94.000 ;
        RECT 62.000 94.300 62.800 99.800 ;
        RECT 70.000 99.200 74.000 99.800 ;
        RECT 70.000 95.800 70.800 99.200 ;
        RECT 71.600 95.800 72.400 98.600 ;
        RECT 73.200 96.000 74.000 99.200 ;
        RECT 76.400 96.000 77.200 99.800 ;
        RECT 73.200 95.800 77.200 96.000 ;
        RECT 71.600 94.400 72.200 95.800 ;
        RECT 73.400 95.400 77.000 95.800 ;
        RECT 75.600 94.400 76.400 94.800 ;
        RECT 70.000 94.300 70.800 94.400 ;
        RECT 62.000 93.700 70.800 94.300 ;
        RECT 71.600 93.800 74.000 94.400 ;
        RECT 75.600 94.300 77.200 94.400 ;
        RECT 78.000 94.300 78.800 99.800 ;
        RECT 79.600 96.300 80.400 97.200 ;
        RECT 82.800 96.300 83.600 99.800 ;
        RECT 79.600 95.700 83.600 96.300 ;
        RECT 79.600 95.600 80.400 95.700 ;
        RECT 75.600 93.800 78.800 94.300 ;
        RECT 55.200 93.600 59.600 93.700 ;
        RECT 55.200 93.400 58.000 93.600 ;
        RECT 55.200 93.200 56.000 93.400 ;
        RECT 52.400 92.300 53.200 92.400 ;
        RECT 46.000 91.700 53.200 92.300 ;
        RECT 46.000 91.600 46.800 91.700 ;
        RECT 52.400 91.600 53.200 91.700 ;
        RECT 54.000 91.600 54.800 92.400 ;
        RECT 56.600 92.200 57.400 92.400 ;
        RECT 55.800 91.600 57.400 92.200 ;
        RECT 54.000 90.200 54.600 91.600 ;
        RECT 55.800 91.400 56.600 91.600 ;
        RECT 38.400 86.800 40.400 87.400 ;
        RECT 30.000 82.200 30.800 85.000 ;
        RECT 31.600 82.200 32.400 85.000 ;
        RECT 34.800 82.200 35.600 86.800 ;
        RECT 38.400 86.200 39.000 86.800 ;
        RECT 38.000 85.600 39.000 86.200 ;
        RECT 38.000 82.200 38.800 85.600 ;
        RECT 43.800 82.200 45.800 90.200 ;
        RECT 49.200 89.600 51.600 90.200 ;
        RECT 49.200 82.200 50.000 89.600 ;
        RECT 50.800 89.400 51.600 89.600 ;
        RECT 53.600 82.200 55.200 90.200 ;
        RECT 57.000 89.600 59.600 90.200 ;
        RECT 57.000 89.400 57.800 89.600 ;
        RECT 58.800 82.200 59.600 89.600 ;
        RECT 62.000 82.200 62.800 93.700 ;
        RECT 70.000 92.800 70.800 93.700 ;
        RECT 73.200 93.600 74.000 93.800 ;
        RECT 76.400 93.700 78.800 93.800 ;
        RECT 76.400 93.600 77.200 93.700 ;
        RECT 71.600 91.600 72.400 93.200 ;
        RECT 73.400 90.200 74.000 93.600 ;
        RECT 74.800 91.600 75.600 93.200 ;
        RECT 72.600 82.200 74.600 90.200 ;
        RECT 78.000 82.200 78.800 93.700 ;
        RECT 82.600 95.200 83.600 95.700 ;
        RECT 82.600 90.800 83.400 95.200 ;
        RECT 84.400 94.600 85.200 99.800 ;
        RECT 90.800 96.600 91.600 99.800 ;
        RECT 92.400 97.000 93.200 99.800 ;
        RECT 94.000 97.000 94.800 99.800 ;
        RECT 95.600 97.000 96.400 99.800 ;
        RECT 97.200 97.000 98.000 99.800 ;
        RECT 100.400 97.000 101.200 99.800 ;
        RECT 103.600 97.000 104.400 99.800 ;
        RECT 105.200 97.000 106.000 99.800 ;
        RECT 106.800 97.000 107.600 99.800 ;
        RECT 89.200 95.800 91.600 96.600 ;
        RECT 108.400 96.600 109.200 99.800 ;
        RECT 89.200 95.200 90.000 95.800 ;
        RECT 84.000 94.000 85.200 94.600 ;
        RECT 88.200 94.600 90.000 95.200 ;
        RECT 94.000 95.600 95.000 96.400 ;
        RECT 98.000 95.600 99.600 96.400 ;
        RECT 100.400 95.800 105.000 96.400 ;
        RECT 108.400 95.800 111.000 96.600 ;
        RECT 100.400 95.600 101.200 95.800 ;
        RECT 84.000 92.000 84.600 94.000 ;
        RECT 88.200 93.400 89.000 94.600 ;
        RECT 85.200 92.600 89.000 93.400 ;
        RECT 94.000 92.800 94.800 95.600 ;
        RECT 100.400 94.800 101.200 95.000 ;
        RECT 96.800 94.200 101.200 94.800 ;
        RECT 96.800 94.000 97.600 94.200 ;
        RECT 102.000 93.600 102.800 95.200 ;
        RECT 104.200 93.400 105.000 95.800 ;
        RECT 110.200 95.200 111.000 95.800 ;
        RECT 110.200 94.400 113.200 95.200 ;
        RECT 114.800 93.800 115.600 99.800 ;
        RECT 97.200 92.600 100.400 93.400 ;
        RECT 104.200 92.600 106.200 93.400 ;
        RECT 106.800 93.000 115.600 93.800 ;
        RECT 90.800 92.000 91.600 92.600 ;
        RECT 108.400 92.000 109.200 92.400 ;
        RECT 113.200 92.200 114.000 92.400 ;
        RECT 113.200 92.000 114.200 92.200 ;
        RECT 84.000 91.400 84.800 92.000 ;
        RECT 90.800 91.400 114.200 92.000 ;
        RECT 82.600 90.000 83.600 90.800 ;
        RECT 82.800 82.200 83.600 90.000 ;
        RECT 84.200 89.600 84.800 91.400 ;
        RECT 84.200 89.000 93.200 89.600 ;
        RECT 84.200 87.400 84.800 89.000 ;
        RECT 92.400 88.800 93.200 89.000 ;
        RECT 95.600 89.000 104.200 89.600 ;
        RECT 95.600 88.800 96.400 89.000 ;
        RECT 87.400 87.600 90.000 88.400 ;
        RECT 84.200 86.800 86.800 87.400 ;
        RECT 86.000 82.200 86.800 86.800 ;
        RECT 89.200 82.200 90.000 87.600 ;
        RECT 90.600 86.800 94.800 87.600 ;
        RECT 92.400 82.200 93.200 85.000 ;
        RECT 94.000 82.200 94.800 85.000 ;
        RECT 95.600 82.200 96.400 85.000 ;
        RECT 97.200 82.200 98.000 88.400 ;
        RECT 100.400 87.600 103.000 88.400 ;
        RECT 103.600 88.200 104.200 89.000 ;
        RECT 105.200 89.400 106.000 89.600 ;
        RECT 105.200 89.000 110.600 89.400 ;
        RECT 105.200 88.800 111.400 89.000 ;
        RECT 110.000 88.200 111.400 88.800 ;
        RECT 103.600 87.600 109.400 88.200 ;
        RECT 112.400 88.000 114.000 88.800 ;
        RECT 112.400 87.600 113.000 88.000 ;
        RECT 100.400 82.200 101.200 87.000 ;
        RECT 103.600 82.200 104.400 87.000 ;
        RECT 108.800 86.800 113.000 87.600 ;
        RECT 114.800 87.400 115.600 93.000 ;
        RECT 113.600 86.800 115.600 87.400 ;
        RECT 116.400 93.800 117.200 99.800 ;
        RECT 122.800 96.600 123.600 99.800 ;
        RECT 124.400 97.000 125.200 99.800 ;
        RECT 126.000 97.000 126.800 99.800 ;
        RECT 127.600 97.000 128.400 99.800 ;
        RECT 130.800 97.000 131.600 99.800 ;
        RECT 134.000 97.000 134.800 99.800 ;
        RECT 135.600 97.000 136.400 99.800 ;
        RECT 137.200 97.000 138.000 99.800 ;
        RECT 138.800 97.000 139.600 99.800 ;
        RECT 121.000 95.800 123.600 96.600 ;
        RECT 140.400 96.600 141.200 99.800 ;
        RECT 127.000 95.800 131.600 96.400 ;
        RECT 121.000 95.200 121.800 95.800 ;
        RECT 118.800 94.400 121.800 95.200 ;
        RECT 116.400 93.000 125.200 93.800 ;
        RECT 127.000 93.400 127.800 95.800 ;
        RECT 130.800 95.600 131.600 95.800 ;
        RECT 132.400 95.600 134.000 96.400 ;
        RECT 137.000 95.600 138.000 96.400 ;
        RECT 140.400 95.800 142.800 96.600 ;
        RECT 129.200 93.600 130.000 95.200 ;
        RECT 130.800 94.800 131.600 95.000 ;
        RECT 130.800 94.200 135.200 94.800 ;
        RECT 134.400 94.000 135.200 94.200 ;
        RECT 116.400 87.400 117.200 93.000 ;
        RECT 125.800 92.600 127.800 93.400 ;
        RECT 131.600 92.600 134.800 93.400 ;
        RECT 137.200 92.800 138.000 95.600 ;
        RECT 142.000 95.200 142.800 95.800 ;
        RECT 142.000 94.600 143.800 95.200 ;
        RECT 143.000 93.400 143.800 94.600 ;
        RECT 146.800 94.600 147.600 99.800 ;
        RECT 148.400 96.000 149.200 99.800 ;
        RECT 148.400 95.200 149.400 96.000 ;
        RECT 151.600 95.800 152.400 99.800 ;
        RECT 153.200 96.000 154.000 99.800 ;
        RECT 156.400 96.000 157.200 99.800 ;
        RECT 153.200 95.800 157.200 96.000 ;
        RECT 146.800 94.000 148.000 94.600 ;
        RECT 143.000 92.600 146.800 93.400 ;
        RECT 117.800 92.000 118.600 92.200 ;
        RECT 119.600 92.000 120.400 92.400 ;
        RECT 122.800 92.000 123.600 92.400 ;
        RECT 140.400 92.000 141.200 92.600 ;
        RECT 147.400 92.000 148.000 94.000 ;
        RECT 117.800 91.400 141.200 92.000 ;
        RECT 147.200 91.400 148.000 92.000 ;
        RECT 147.200 89.600 147.800 91.400 ;
        RECT 148.600 90.800 149.400 95.200 ;
        RECT 151.800 94.400 152.400 95.800 ;
        RECT 153.400 95.400 157.000 95.800 ;
        RECT 158.000 95.600 158.800 97.200 ;
        RECT 155.600 94.400 156.400 94.800 ;
        RECT 151.600 93.600 154.200 94.400 ;
        RECT 155.600 94.300 157.200 94.400 ;
        RECT 159.600 94.300 160.400 99.800 ;
        RECT 155.600 93.800 160.400 94.300 ;
        RECT 156.400 93.700 160.400 93.800 ;
        RECT 156.400 93.600 157.200 93.700 ;
        RECT 151.600 92.300 152.400 92.400 ;
        RECT 153.600 92.300 154.200 93.600 ;
        RECT 151.600 91.700 154.200 92.300 ;
        RECT 151.600 91.600 152.400 91.700 ;
        RECT 126.000 89.400 126.800 89.600 ;
        RECT 121.400 89.000 126.800 89.400 ;
        RECT 120.600 88.800 126.800 89.000 ;
        RECT 127.800 89.000 136.400 89.600 ;
        RECT 118.000 88.000 119.600 88.800 ;
        RECT 120.600 88.200 122.000 88.800 ;
        RECT 127.800 88.200 128.400 89.000 ;
        RECT 135.600 88.800 136.400 89.000 ;
        RECT 138.800 89.000 147.800 89.600 ;
        RECT 138.800 88.800 139.600 89.000 ;
        RECT 119.000 87.600 119.600 88.000 ;
        RECT 122.600 87.600 128.400 88.200 ;
        RECT 129.000 87.600 131.600 88.400 ;
        RECT 116.400 86.800 118.400 87.400 ;
        RECT 119.000 86.800 123.200 87.600 ;
        RECT 105.200 82.200 106.000 85.000 ;
        RECT 106.800 82.200 107.600 85.000 ;
        RECT 110.000 82.200 110.800 86.800 ;
        RECT 113.600 86.200 114.200 86.800 ;
        RECT 113.200 85.600 114.200 86.200 ;
        RECT 117.800 86.200 118.400 86.800 ;
        RECT 117.800 85.600 118.800 86.200 ;
        RECT 113.200 82.200 114.000 85.600 ;
        RECT 118.000 82.200 118.800 85.600 ;
        RECT 121.200 82.200 122.000 86.800 ;
        RECT 124.400 82.200 125.200 85.000 ;
        RECT 126.000 82.200 126.800 85.000 ;
        RECT 127.600 82.200 128.400 87.000 ;
        RECT 130.800 82.200 131.600 87.000 ;
        RECT 134.000 82.200 134.800 88.400 ;
        RECT 142.000 87.600 144.600 88.400 ;
        RECT 137.200 86.800 141.400 87.600 ;
        RECT 135.600 82.200 136.400 85.000 ;
        RECT 137.200 82.200 138.000 85.000 ;
        RECT 138.800 82.200 139.600 85.000 ;
        RECT 142.000 82.200 142.800 87.600 ;
        RECT 147.200 87.400 147.800 89.000 ;
        RECT 145.200 86.800 147.800 87.400 ;
        RECT 148.400 90.000 149.400 90.800 ;
        RECT 150.000 90.300 150.800 90.400 ;
        RECT 151.600 90.300 152.400 90.400 ;
        RECT 150.000 90.200 152.400 90.300 ;
        RECT 153.600 90.200 154.200 91.700 ;
        RECT 154.800 91.600 155.600 93.200 ;
        RECT 159.600 92.300 160.400 93.700 ;
        RECT 162.800 97.600 163.600 99.800 ;
        RECT 167.600 97.800 168.400 99.800 ;
        RECT 172.400 97.800 173.200 99.800 ;
        RECT 162.800 94.400 163.400 97.600 ;
        RECT 164.400 95.600 165.200 97.200 ;
        RECT 166.000 95.600 166.800 97.200 ;
        RECT 167.800 94.400 168.400 97.800 ;
        RECT 170.800 95.600 171.600 97.200 ;
        RECT 172.600 94.400 173.200 97.800 ;
        RECT 176.200 96.400 177.000 99.800 ;
        RECT 176.200 95.800 178.000 96.400 ;
        RECT 162.800 93.600 163.600 94.400 ;
        RECT 167.600 93.600 168.400 94.400 ;
        RECT 172.400 93.600 173.200 94.400 ;
        RECT 161.200 92.300 162.000 92.400 ;
        RECT 159.600 91.700 162.000 92.300 ;
        RECT 145.200 82.200 146.000 86.800 ;
        RECT 148.400 82.200 149.200 90.000 ;
        RECT 150.000 89.700 153.000 90.200 ;
        RECT 150.000 89.600 150.800 89.700 ;
        RECT 151.600 89.600 153.000 89.700 ;
        RECT 153.600 89.600 154.600 90.200 ;
        RECT 152.400 88.400 153.000 89.600 ;
        RECT 152.400 87.600 153.200 88.400 ;
        RECT 153.800 82.200 154.600 89.600 ;
        RECT 159.600 82.200 160.400 91.700 ;
        RECT 161.200 90.800 162.000 91.700 ;
        RECT 162.800 90.200 163.400 93.600 ;
        RECT 167.800 90.200 168.400 93.600 ;
        RECT 169.200 90.800 170.000 92.400 ;
        RECT 172.600 90.200 173.200 93.600 ;
        RECT 174.000 92.300 174.800 92.400 ;
        RECT 177.200 92.300 178.000 95.800 ;
        RECT 180.400 95.600 181.200 97.200 ;
        RECT 178.800 93.600 179.600 95.200 ;
        RECT 174.000 91.700 178.000 92.300 ;
        RECT 174.000 90.800 174.800 91.700 ;
        RECT 161.800 89.400 163.600 90.200 ;
        RECT 167.600 89.400 169.400 90.200 ;
        RECT 172.400 89.400 174.200 90.200 ;
        RECT 161.800 84.400 162.600 89.400 ;
        RECT 161.200 83.600 162.600 84.400 ;
        RECT 161.800 82.200 162.600 83.600 ;
        RECT 168.600 88.400 169.400 89.400 ;
        RECT 168.600 87.600 170.000 88.400 ;
        RECT 168.600 82.200 169.400 87.600 ;
        RECT 173.400 84.400 174.200 89.400 ;
        RECT 175.600 88.800 176.400 90.400 ;
        RECT 172.400 83.600 174.200 84.400 ;
        RECT 173.400 82.200 174.200 83.600 ;
        RECT 177.200 82.200 178.000 91.700 ;
        RECT 182.000 90.300 182.800 99.800 ;
        RECT 193.600 94.200 194.400 99.800 ;
        RECT 197.000 98.400 197.800 99.800 ;
        RECT 196.400 97.600 197.800 98.400 ;
        RECT 197.000 96.400 197.800 97.600 ;
        RECT 197.000 95.800 198.800 96.400 ;
        RECT 201.200 96.000 202.000 99.800 ;
        RECT 204.400 96.000 205.200 99.800 ;
        RECT 201.200 95.800 205.200 96.000 ;
        RECT 206.000 95.800 206.800 99.800 ;
        RECT 207.600 95.800 208.400 99.800 ;
        RECT 209.200 96.000 210.000 99.800 ;
        RECT 212.400 96.000 213.200 99.800 ;
        RECT 214.600 96.400 215.400 99.800 ;
        RECT 220.400 97.800 221.200 99.800 ;
        RECT 209.200 95.800 213.200 96.000 ;
        RECT 193.600 93.800 195.400 94.200 ;
        RECT 193.800 93.600 195.400 93.800 ;
        RECT 191.600 91.600 193.200 92.400 ;
        RECT 190.000 90.300 190.800 91.200 ;
        RECT 182.000 89.700 190.800 90.300 ;
        RECT 182.000 82.200 182.800 89.700 ;
        RECT 190.000 89.600 190.800 89.700 ;
        RECT 194.800 90.400 195.400 93.600 ;
        RECT 194.800 89.600 195.600 90.400 ;
        RECT 193.200 87.600 194.000 89.200 ;
        RECT 194.800 87.000 195.400 89.600 ;
        RECT 196.400 88.800 197.200 90.400 ;
        RECT 191.800 86.400 195.400 87.000 ;
        RECT 191.800 86.200 192.400 86.400 ;
        RECT 191.600 82.200 192.400 86.200 ;
        RECT 194.800 86.200 195.400 86.400 ;
        RECT 194.800 82.200 195.600 86.200 ;
        RECT 198.000 82.200 198.800 95.800 ;
        RECT 201.400 95.400 205.000 95.800 ;
        RECT 199.600 93.600 200.400 95.200 ;
        RECT 202.000 94.400 202.800 94.800 ;
        RECT 206.000 94.400 206.600 95.800 ;
        RECT 207.800 94.400 208.400 95.800 ;
        RECT 209.400 95.400 213.000 95.800 ;
        RECT 214.000 95.600 216.400 96.400 ;
        RECT 211.600 94.400 212.400 94.800 ;
        RECT 201.200 93.800 202.800 94.400 ;
        RECT 201.200 93.600 202.000 93.800 ;
        RECT 204.200 93.600 206.800 94.400 ;
        RECT 207.600 93.600 210.200 94.400 ;
        RECT 211.600 93.800 213.200 94.400 ;
        RECT 212.400 93.600 213.200 93.800 ;
        RECT 202.800 91.600 203.600 93.200 ;
        RECT 204.200 90.200 204.800 93.600 ;
        RECT 206.000 90.200 206.800 90.400 ;
        RECT 203.800 89.600 204.800 90.200 ;
        RECT 205.400 89.600 206.800 90.200 ;
        RECT 207.600 90.200 208.400 90.400 ;
        RECT 209.600 90.200 210.200 93.600 ;
        RECT 210.800 91.600 211.600 93.200 ;
        RECT 207.600 89.600 209.000 90.200 ;
        RECT 209.600 89.600 210.600 90.200 ;
        RECT 203.800 84.400 204.600 89.600 ;
        RECT 205.400 88.400 206.000 89.600 ;
        RECT 205.200 87.600 206.000 88.400 ;
        RECT 208.400 88.400 209.000 89.600 ;
        RECT 209.800 88.400 210.600 89.600 ;
        RECT 214.000 88.800 214.800 90.400 ;
        RECT 208.400 87.600 209.200 88.400 ;
        RECT 209.800 87.600 211.600 88.400 ;
        RECT 202.800 83.600 204.600 84.400 ;
        RECT 203.800 82.200 204.600 83.600 ;
        RECT 209.800 82.200 210.600 87.600 ;
        RECT 215.600 82.200 216.400 95.600 ;
        RECT 217.200 93.600 218.000 95.200 ;
        RECT 220.400 94.400 221.000 97.800 ;
        RECT 222.000 95.600 222.800 97.200 ;
        RECT 226.800 95.800 227.600 99.800 ;
        RECT 228.200 96.400 229.000 97.200 ;
        RECT 230.600 96.800 231.400 99.800 ;
        RECT 220.400 93.600 221.200 94.400 ;
        RECT 218.800 90.800 219.600 92.400 ;
        RECT 220.400 90.200 221.000 93.600 ;
        RECT 225.200 92.800 226.000 94.400 ;
        RECT 223.600 92.200 224.400 92.400 ;
        RECT 226.800 92.200 227.400 95.800 ;
        RECT 228.400 95.600 229.200 96.400 ;
        RECT 230.000 95.800 231.400 96.800 ;
        RECT 234.800 95.800 235.600 99.800 ;
        RECT 230.000 92.400 230.600 95.800 ;
        RECT 234.800 95.600 235.400 95.800 ;
        RECT 233.600 95.200 235.400 95.600 ;
        RECT 231.200 95.000 235.400 95.200 ;
        RECT 231.200 94.600 234.200 95.000 ;
        RECT 231.200 94.400 232.000 94.600 ;
        RECT 228.400 92.200 229.200 92.400 ;
        RECT 223.600 91.600 225.200 92.200 ;
        RECT 226.800 91.600 229.200 92.200 ;
        RECT 230.000 91.600 230.800 92.400 ;
        RECT 224.400 91.200 225.200 91.600 ;
        RECT 228.400 90.200 229.000 91.600 ;
        RECT 230.000 90.200 230.600 91.600 ;
        RECT 231.400 91.000 232.000 94.400 ;
        RECT 232.800 93.800 233.600 94.000 ;
        RECT 232.800 93.200 233.800 93.800 ;
        RECT 233.200 92.400 233.800 93.200 ;
        RECT 234.800 92.800 235.600 94.400 ;
        RECT 233.200 91.600 234.000 92.400 ;
        RECT 231.400 90.400 233.800 91.000 ;
        RECT 219.400 89.400 221.200 90.200 ;
        RECT 223.600 89.600 227.600 90.200 ;
        RECT 217.200 88.300 218.000 88.400 ;
        RECT 219.400 88.300 220.200 89.400 ;
        RECT 217.200 87.700 220.200 88.300 ;
        RECT 217.200 87.600 218.000 87.700 ;
        RECT 219.400 82.200 220.200 87.700 ;
        RECT 223.600 82.200 224.400 89.600 ;
        RECT 226.800 82.200 227.600 89.600 ;
        RECT 228.400 82.200 229.200 90.200 ;
        RECT 230.000 82.200 230.800 90.200 ;
        RECT 233.200 86.200 233.800 90.400 ;
        RECT 234.800 90.300 235.600 90.400 ;
        RECT 236.400 90.300 237.200 99.800 ;
        RECT 238.000 95.600 238.800 97.200 ;
        RECT 239.600 95.800 240.400 99.800 ;
        RECT 241.200 96.000 242.000 99.800 ;
        RECT 244.400 96.000 245.200 99.800 ;
        RECT 246.200 96.400 247.000 97.200 ;
        RECT 241.200 95.800 245.200 96.000 ;
        RECT 239.800 94.400 240.400 95.800 ;
        RECT 241.400 95.400 245.000 95.800 ;
        RECT 246.000 95.600 246.800 96.400 ;
        RECT 247.600 95.800 248.400 99.800 ;
        RECT 239.600 93.600 242.200 94.400 ;
        RECT 234.800 89.700 237.200 90.300 ;
        RECT 234.800 89.600 235.600 89.700 ;
        RECT 233.200 82.200 234.000 86.200 ;
        RECT 236.400 82.200 237.200 89.700 ;
        RECT 239.600 90.200 240.400 90.400 ;
        RECT 241.600 90.200 242.200 93.600 ;
        RECT 242.800 91.600 243.600 93.200 ;
        RECT 246.000 92.200 246.800 92.400 ;
        RECT 247.800 92.200 248.400 95.800 ;
        RECT 249.200 92.800 250.000 94.400 ;
        RECT 246.000 91.600 248.400 92.200 ;
        RECT 246.200 90.200 246.800 91.600 ;
        RECT 239.600 89.600 241.000 90.200 ;
        RECT 241.600 89.600 242.600 90.200 ;
        RECT 240.400 88.400 241.000 89.600 ;
        RECT 240.400 87.600 241.200 88.400 ;
        RECT 241.800 82.200 242.600 89.600 ;
        RECT 246.000 82.200 246.800 90.200 ;
        RECT 247.600 89.600 251.600 90.200 ;
        RECT 247.600 82.200 248.400 89.600 ;
        RECT 250.800 82.200 251.600 89.600 ;
        RECT 4.400 72.400 5.200 79.800 ;
        RECT 3.000 71.800 5.200 72.400 ;
        RECT 3.000 71.200 3.600 71.800 ;
        RECT 2.400 70.400 3.600 71.200 ;
        RECT 7.600 71.200 8.400 79.800 ;
        RECT 10.800 71.200 11.600 79.800 ;
        RECT 14.000 71.200 14.800 79.800 ;
        RECT 17.200 71.200 18.000 79.800 ;
        RECT 22.000 71.200 22.800 79.800 ;
        RECT 25.200 71.200 26.000 79.800 ;
        RECT 28.400 71.200 29.200 79.800 ;
        RECT 31.600 71.200 32.400 79.800 ;
        RECT 7.600 70.400 9.400 71.200 ;
        RECT 10.800 70.400 13.000 71.200 ;
        RECT 14.000 70.400 16.200 71.200 ;
        RECT 17.200 70.400 19.600 71.200 ;
        RECT 22.000 70.400 23.800 71.200 ;
        RECT 25.200 70.400 27.400 71.200 ;
        RECT 28.400 70.400 30.600 71.200 ;
        RECT 31.600 70.400 34.000 71.200 ;
        RECT 3.000 67.400 3.600 70.400 ;
        RECT 4.400 68.800 5.200 70.400 ;
        RECT 8.600 69.000 9.400 70.400 ;
        RECT 12.200 69.000 13.000 70.400 ;
        RECT 15.400 69.000 16.200 70.400 ;
        RECT 8.600 68.200 11.200 69.000 ;
        RECT 12.200 68.200 14.600 69.000 ;
        RECT 15.400 68.200 18.000 69.000 ;
        RECT 8.600 67.600 9.400 68.200 ;
        RECT 12.200 67.600 13.000 68.200 ;
        RECT 15.400 67.600 16.200 68.200 ;
        RECT 18.800 67.600 19.600 70.400 ;
        RECT 23.000 69.000 23.800 70.400 ;
        RECT 26.600 69.000 27.400 70.400 ;
        RECT 29.800 69.000 30.600 70.400 ;
        RECT 23.000 68.200 25.600 69.000 ;
        RECT 26.600 68.200 29.000 69.000 ;
        RECT 29.800 68.200 32.400 69.000 ;
        RECT 23.000 67.600 23.800 68.200 ;
        RECT 26.600 67.600 27.400 68.200 ;
        RECT 29.800 67.600 30.600 68.200 ;
        RECT 33.200 67.600 34.000 70.400 ;
        RECT 3.000 66.800 5.200 67.400 ;
        RECT 4.400 62.200 5.200 66.800 ;
        RECT 7.600 66.800 9.400 67.600 ;
        RECT 10.800 66.800 13.000 67.600 ;
        RECT 14.000 66.800 16.200 67.600 ;
        RECT 17.200 66.800 19.600 67.600 ;
        RECT 22.000 66.800 23.800 67.600 ;
        RECT 25.200 66.800 27.400 67.600 ;
        RECT 28.400 66.800 30.600 67.600 ;
        RECT 31.600 66.800 34.000 67.600 ;
        RECT 7.600 62.200 8.400 66.800 ;
        RECT 10.800 62.200 11.600 66.800 ;
        RECT 14.000 62.200 14.800 66.800 ;
        RECT 17.200 62.200 18.000 66.800 ;
        RECT 22.000 62.200 22.800 66.800 ;
        RECT 25.200 62.200 26.000 66.800 ;
        RECT 28.400 62.200 29.200 66.800 ;
        RECT 31.600 62.200 32.400 66.800 ;
        RECT 34.800 64.800 35.600 66.400 ;
        RECT 36.400 62.200 37.200 79.800 ;
        RECT 40.600 71.800 42.600 79.800 ;
        RECT 48.600 71.800 50.600 79.800 ;
        RECT 39.600 68.800 40.400 70.400 ;
        RECT 41.200 68.400 41.800 71.800 ;
        RECT 42.800 68.800 43.600 70.400 ;
        RECT 38.000 68.200 38.800 68.400 ;
        RECT 41.200 68.200 42.000 68.400 ;
        RECT 38.000 67.600 39.600 68.200 ;
        RECT 41.200 67.600 43.600 68.200 ;
        RECT 44.400 67.600 45.200 69.200 ;
        RECT 46.000 67.600 46.800 70.400 ;
        RECT 47.600 68.800 48.400 70.400 ;
        RECT 49.400 68.400 50.000 71.800 ;
        RECT 50.800 70.300 51.600 70.400 ;
        RECT 52.400 70.300 53.200 70.400 ;
        RECT 50.800 69.700 53.200 70.300 ;
        RECT 50.800 68.800 51.600 69.700 ;
        RECT 52.400 69.600 53.200 69.700 ;
        RECT 49.200 68.200 50.000 68.400 ;
        RECT 52.400 68.200 53.200 68.400 ;
        RECT 47.600 67.600 50.000 68.200 ;
        RECT 51.600 67.600 53.200 68.200 ;
        RECT 38.800 67.200 39.600 67.600 ;
        RECT 38.200 66.200 41.800 66.600 ;
        RECT 43.000 66.200 43.600 67.600 ;
        RECT 47.600 66.200 48.200 67.600 ;
        RECT 51.600 67.200 52.400 67.600 ;
        RECT 49.400 66.200 53.000 66.600 ;
        RECT 38.000 66.000 42.000 66.200 ;
        RECT 38.000 62.200 38.800 66.000 ;
        RECT 41.200 62.800 42.000 66.000 ;
        RECT 42.800 63.400 43.600 66.200 ;
        RECT 44.400 62.800 45.200 66.200 ;
        RECT 41.200 62.200 45.200 62.800 ;
        RECT 46.000 62.800 46.800 66.200 ;
        RECT 47.600 63.400 48.400 66.200 ;
        RECT 49.200 66.000 53.200 66.200 ;
        RECT 49.200 62.800 50.000 66.000 ;
        RECT 46.000 62.200 50.000 62.800 ;
        RECT 52.400 62.200 53.200 66.000 ;
        RECT 55.600 62.200 56.400 79.800 ;
        RECT 66.800 71.200 67.600 79.800 ;
        RECT 70.000 71.200 70.800 79.800 ;
        RECT 73.200 71.200 74.000 79.800 ;
        RECT 76.400 71.200 77.200 79.800 ;
        RECT 79.600 71.800 80.400 79.800 ;
        RECT 82.800 72.400 83.600 79.800 ;
        RECT 86.000 76.400 86.800 79.800 ;
        RECT 85.800 75.800 86.800 76.400 ;
        RECT 85.800 75.200 86.400 75.800 ;
        RECT 89.200 75.200 90.000 79.800 ;
        RECT 92.400 77.000 93.200 79.800 ;
        RECT 94.000 77.000 94.800 79.800 ;
        RECT 81.400 71.800 83.600 72.400 ;
        RECT 84.400 74.600 86.400 75.200 ;
        RECT 66.800 70.400 68.600 71.200 ;
        RECT 70.000 70.400 72.200 71.200 ;
        RECT 73.200 70.400 75.400 71.200 ;
        RECT 76.400 70.400 78.800 71.200 ;
        RECT 67.800 69.000 68.600 70.400 ;
        RECT 71.400 69.000 72.200 70.400 ;
        RECT 74.600 69.000 75.400 70.400 ;
        RECT 57.200 66.800 58.000 68.400 ;
        RECT 67.800 68.200 70.400 69.000 ;
        RECT 71.400 68.200 73.800 69.000 ;
        RECT 74.600 68.200 77.200 69.000 ;
        RECT 67.800 67.600 68.600 68.200 ;
        RECT 71.400 67.600 72.200 68.200 ;
        RECT 74.600 67.600 75.400 68.200 ;
        RECT 78.000 67.600 78.800 70.400 ;
        RECT 66.800 66.800 68.600 67.600 ;
        RECT 70.000 66.800 72.200 67.600 ;
        RECT 73.200 66.800 75.400 67.600 ;
        RECT 76.400 66.800 78.800 67.600 ;
        RECT 79.600 69.600 80.200 71.800 ;
        RECT 81.400 71.200 82.000 71.800 ;
        RECT 80.800 70.400 82.000 71.200 ;
        RECT 66.800 62.200 67.600 66.800 ;
        RECT 70.000 62.200 70.800 66.800 ;
        RECT 73.200 62.200 74.000 66.800 ;
        RECT 76.400 62.200 77.200 66.800 ;
        RECT 79.600 62.200 80.400 69.600 ;
        RECT 81.400 67.400 82.000 70.400 ;
        RECT 82.800 68.800 83.600 70.400 ;
        RECT 84.400 69.000 85.200 74.600 ;
        RECT 87.000 74.400 91.200 75.200 ;
        RECT 95.600 75.000 96.400 79.800 ;
        RECT 98.800 75.000 99.600 79.800 ;
        RECT 87.000 74.000 87.600 74.400 ;
        RECT 86.000 73.200 87.600 74.000 ;
        RECT 90.600 73.800 96.400 74.400 ;
        RECT 88.600 73.200 90.000 73.800 ;
        RECT 88.600 73.000 94.800 73.200 ;
        RECT 89.400 72.600 94.800 73.000 ;
        RECT 94.000 72.400 94.800 72.600 ;
        RECT 95.800 73.000 96.400 73.800 ;
        RECT 97.000 73.600 99.600 74.400 ;
        RECT 102.000 73.600 102.800 79.800 ;
        RECT 103.600 77.000 104.400 79.800 ;
        RECT 105.200 77.000 106.000 79.800 ;
        RECT 106.800 77.000 107.600 79.800 ;
        RECT 105.200 74.400 109.400 75.200 ;
        RECT 110.000 74.400 110.800 79.800 ;
        RECT 113.200 75.200 114.000 79.800 ;
        RECT 113.200 74.600 115.800 75.200 ;
        RECT 110.000 73.600 112.600 74.400 ;
        RECT 103.600 73.000 104.400 73.200 ;
        RECT 95.800 72.400 104.400 73.000 ;
        RECT 106.800 73.000 107.600 73.200 ;
        RECT 115.200 73.000 115.800 74.600 ;
        RECT 106.800 72.400 115.800 73.000 ;
        RECT 115.200 70.600 115.800 72.400 ;
        RECT 116.400 72.000 117.200 79.800 ;
        RECT 116.400 71.200 117.400 72.000 ;
        RECT 85.800 70.000 109.200 70.600 ;
        RECT 115.200 70.000 116.000 70.600 ;
        RECT 85.800 69.800 86.600 70.000 ;
        RECT 90.800 69.600 91.600 70.000 ;
        RECT 108.400 69.400 109.200 70.000 ;
        RECT 84.400 68.200 93.200 69.000 ;
        RECT 93.800 68.600 95.800 69.400 ;
        RECT 99.600 68.600 102.800 69.400 ;
        RECT 81.400 66.800 83.600 67.400 ;
        RECT 82.800 62.200 83.600 66.800 ;
        RECT 84.400 62.200 85.200 68.200 ;
        RECT 86.800 66.800 89.800 67.600 ;
        RECT 89.000 66.200 89.800 66.800 ;
        RECT 95.000 66.200 95.800 68.600 ;
        RECT 97.200 66.800 98.000 68.400 ;
        RECT 102.400 67.800 103.200 68.000 ;
        RECT 98.800 67.200 103.200 67.800 ;
        RECT 98.800 67.000 99.600 67.200 ;
        RECT 105.200 66.400 106.000 69.200 ;
        RECT 111.000 68.600 114.800 69.400 ;
        RECT 111.000 67.400 111.800 68.600 ;
        RECT 115.400 68.000 116.000 70.000 ;
        RECT 98.800 66.200 99.600 66.400 ;
        RECT 89.000 65.400 91.600 66.200 ;
        RECT 95.000 65.600 99.600 66.200 ;
        RECT 100.400 65.600 102.000 66.400 ;
        RECT 105.000 65.600 106.000 66.400 ;
        RECT 110.000 66.800 111.800 67.400 ;
        RECT 114.800 67.400 116.000 68.000 ;
        RECT 110.000 66.200 110.800 66.800 ;
        RECT 90.800 62.200 91.600 65.400 ;
        RECT 108.400 65.400 110.800 66.200 ;
        RECT 92.400 62.200 93.200 65.000 ;
        RECT 94.000 62.200 94.800 65.000 ;
        RECT 95.600 62.200 96.400 65.000 ;
        RECT 98.800 62.200 99.600 65.000 ;
        RECT 102.000 62.200 102.800 65.000 ;
        RECT 103.600 62.200 104.400 65.000 ;
        RECT 105.200 62.200 106.000 65.000 ;
        RECT 106.800 62.200 107.600 65.000 ;
        RECT 108.400 62.200 109.200 65.400 ;
        RECT 114.800 62.200 115.600 67.400 ;
        RECT 116.600 66.800 117.400 71.200 ;
        RECT 119.600 71.800 120.400 79.800 ;
        RECT 122.800 75.800 123.600 79.800 ;
        RECT 119.600 70.400 120.200 71.800 ;
        RECT 122.800 71.600 123.400 75.800 ;
        RECT 126.000 72.400 126.800 79.800 ;
        RECT 126.000 71.800 128.200 72.400 ;
        RECT 129.200 71.800 130.000 79.800 ;
        RECT 131.000 79.200 134.600 79.800 ;
        RECT 131.000 79.000 131.600 79.200 ;
        RECT 130.800 73.000 131.600 79.000 ;
        RECT 134.000 79.000 134.600 79.200 ;
        RECT 135.600 79.200 139.600 79.800 ;
        RECT 132.400 73.000 133.200 78.600 ;
        RECT 134.000 73.400 134.800 79.000 ;
        RECT 135.600 74.000 136.400 79.200 ;
        RECT 137.200 73.800 138.000 78.600 ;
        RECT 138.800 73.800 139.600 79.200 ;
        RECT 137.200 73.400 137.800 73.800 ;
        RECT 134.000 73.000 137.800 73.400 ;
        RECT 132.600 72.400 133.200 73.000 ;
        RECT 134.200 72.800 137.800 73.000 ;
        RECT 139.000 73.200 139.600 73.800 ;
        RECT 142.000 73.800 142.800 79.800 ;
        RECT 142.000 73.200 142.600 73.800 ;
        RECT 139.000 72.600 142.600 73.200 ;
        RECT 121.000 71.000 123.400 71.600 ;
        RECT 127.600 71.200 128.200 71.800 ;
        RECT 118.000 70.300 118.800 70.400 ;
        RECT 119.600 70.300 120.400 70.400 ;
        RECT 118.000 69.700 120.400 70.300 ;
        RECT 118.000 69.600 118.800 69.700 ;
        RECT 119.600 69.600 120.400 69.700 ;
        RECT 116.400 66.000 117.400 66.800 ;
        RECT 119.600 66.200 120.200 69.600 ;
        RECT 121.000 67.600 121.600 71.000 ;
        RECT 127.600 70.400 128.800 71.200 ;
        RECT 122.800 69.600 123.600 70.400 ;
        RECT 122.800 68.800 123.400 69.600 ;
        RECT 122.400 68.200 123.400 68.800 ;
        RECT 122.400 68.000 123.200 68.200 ;
        RECT 124.400 67.600 125.200 69.200 ;
        RECT 126.000 68.800 126.800 70.400 ;
        RECT 120.800 67.400 121.600 67.600 ;
        RECT 127.600 67.400 128.200 70.400 ;
        RECT 129.400 69.600 130.000 71.800 ;
        RECT 132.400 72.200 133.200 72.400 ;
        RECT 146.200 72.400 147.000 79.800 ;
        RECT 147.600 73.600 148.400 74.400 ;
        RECT 147.800 72.400 148.400 73.600 ;
        RECT 152.600 72.400 153.400 79.800 ;
        RECT 154.000 73.600 154.800 74.400 ;
        RECT 154.200 72.400 154.800 73.600 ;
        RECT 159.000 72.400 159.800 79.800 ;
        RECT 160.400 73.600 161.200 74.400 ;
        RECT 160.600 72.400 161.200 73.600 ;
        RECT 132.400 71.600 135.800 72.200 ;
        RECT 146.200 71.800 147.200 72.400 ;
        RECT 147.800 71.800 149.200 72.400 ;
        RECT 152.600 71.800 153.600 72.400 ;
        RECT 154.200 71.800 155.600 72.400 ;
        RECT 159.000 71.800 160.000 72.400 ;
        RECT 160.600 71.800 162.000 72.400 ;
        RECT 120.800 67.000 123.800 67.400 ;
        RECT 120.800 66.800 125.000 67.000 ;
        RECT 123.200 66.400 125.000 66.800 ;
        RECT 124.400 66.200 125.000 66.400 ;
        RECT 126.000 66.800 128.200 67.400 ;
        RECT 116.400 62.200 117.200 66.000 ;
        RECT 119.600 65.200 121.000 66.200 ;
        RECT 120.200 62.200 121.000 65.200 ;
        RECT 124.400 62.200 125.200 66.200 ;
        RECT 126.000 62.200 126.800 66.800 ;
        RECT 129.200 62.200 130.000 69.600 ;
        RECT 135.200 68.400 135.800 71.600 ;
        RECT 136.400 70.300 138.000 70.400 ;
        RECT 145.200 70.300 146.000 70.400 ;
        RECT 136.400 69.700 146.000 70.300 ;
        RECT 136.400 69.600 138.000 69.700 ;
        RECT 145.200 68.800 146.000 69.700 ;
        RECT 146.600 68.400 147.200 71.800 ;
        RECT 148.400 71.600 149.200 71.800 ;
        RECT 151.600 68.800 152.400 70.400 ;
        RECT 153.000 68.400 153.600 71.800 ;
        RECT 154.800 71.600 155.600 71.800 ;
        RECT 154.800 70.300 155.600 70.400 ;
        RECT 158.000 70.300 158.800 70.400 ;
        RECT 154.800 69.700 158.800 70.300 ;
        RECT 154.800 69.600 155.600 69.700 ;
        RECT 158.000 68.800 158.800 69.700 ;
        RECT 159.400 68.400 160.000 71.800 ;
        RECT 161.200 71.600 162.000 71.800 ;
        RECT 162.800 71.600 163.600 73.200 ;
        RECT 135.200 67.600 136.400 68.400 ;
        RECT 138.000 67.600 139.600 68.400 ;
        RECT 142.000 68.300 142.800 68.400 ;
        RECT 143.600 68.300 144.400 68.400 ;
        RECT 142.000 68.200 144.400 68.300 ;
        RECT 142.000 67.700 145.200 68.200 ;
        RECT 142.000 67.600 142.800 67.700 ;
        RECT 143.600 67.600 145.200 67.700 ;
        RECT 146.600 67.600 149.200 68.400 ;
        RECT 150.000 68.200 150.800 68.400 ;
        RECT 150.000 67.600 151.600 68.200 ;
        RECT 153.000 67.600 155.600 68.400 ;
        RECT 156.400 68.200 157.200 68.400 ;
        RECT 156.400 67.600 158.000 68.200 ;
        RECT 159.400 67.600 162.000 68.400 ;
        RECT 162.800 68.300 163.600 68.400 ;
        RECT 164.400 68.300 165.200 79.800 ;
        RECT 167.600 71.800 168.400 79.800 ;
        RECT 169.200 72.400 170.000 79.800 ;
        RECT 172.400 72.400 173.200 79.800 ;
        RECT 176.600 78.300 177.400 79.800 ;
        RECT 178.800 78.300 179.600 78.400 ;
        RECT 176.600 77.700 179.600 78.300 ;
        RECT 176.600 72.600 177.400 77.700 ;
        RECT 178.800 77.600 179.600 77.700 ;
        RECT 186.800 76.400 187.600 79.800 ;
        RECT 186.600 75.800 187.600 76.400 ;
        RECT 186.600 75.200 187.200 75.800 ;
        RECT 190.000 75.200 190.800 79.800 ;
        RECT 193.200 77.000 194.000 79.800 ;
        RECT 194.800 77.000 195.600 79.800 ;
        RECT 169.200 71.800 173.200 72.400 ;
        RECT 175.600 71.800 177.400 72.600 ;
        RECT 185.200 74.600 187.200 75.200 ;
        RECT 167.800 70.400 168.400 71.800 ;
        RECT 171.600 70.400 172.400 70.800 ;
        RECT 167.600 69.800 170.000 70.400 ;
        RECT 171.600 70.300 173.200 70.400 ;
        RECT 174.000 70.300 174.800 70.400 ;
        RECT 171.600 69.800 174.800 70.300 ;
        RECT 167.600 69.600 168.400 69.800 ;
        RECT 162.800 67.700 165.200 68.300 ;
        RECT 162.800 67.600 163.600 67.700 ;
        RECT 135.200 65.000 135.800 67.600 ;
        RECT 139.400 66.300 141.200 66.400 ;
        RECT 142.100 66.300 142.700 67.600 ;
        RECT 144.400 67.200 145.200 67.600 ;
        RECT 139.400 65.700 142.700 66.300 ;
        RECT 143.800 66.200 147.400 66.600 ;
        RECT 148.400 66.200 149.000 67.600 ;
        RECT 150.800 67.200 151.600 67.600 ;
        RECT 150.200 66.200 153.800 66.600 ;
        RECT 154.800 66.200 155.400 67.600 ;
        RECT 157.200 67.200 158.000 67.600 ;
        RECT 156.600 66.200 160.200 66.600 ;
        RECT 161.200 66.400 161.800 67.600 ;
        RECT 143.600 66.000 147.600 66.200 ;
        RECT 139.400 65.600 141.200 65.700 ;
        RECT 135.200 64.400 139.200 65.000 ;
        RECT 135.200 64.200 136.400 64.400 ;
        RECT 135.600 62.200 136.400 64.200 ;
        RECT 138.600 64.200 139.200 64.400 ;
        RECT 138.600 63.600 139.600 64.200 ;
        RECT 138.800 62.200 139.600 63.600 ;
        RECT 143.600 62.200 144.400 66.000 ;
        RECT 146.800 62.200 147.600 66.000 ;
        RECT 148.400 62.200 149.200 66.200 ;
        RECT 150.000 66.000 154.000 66.200 ;
        RECT 150.000 62.200 150.800 66.000 ;
        RECT 153.200 62.200 154.000 66.000 ;
        RECT 154.800 62.200 155.600 66.200 ;
        RECT 156.400 66.000 160.400 66.200 ;
        RECT 156.400 62.200 157.200 66.000 ;
        RECT 159.600 62.200 160.400 66.000 ;
        RECT 161.200 62.200 162.000 66.400 ;
        RECT 164.400 66.200 165.200 67.700 ;
        RECT 166.000 66.800 166.800 68.400 ;
        RECT 169.400 66.400 170.000 69.800 ;
        RECT 172.400 69.700 174.800 69.800 ;
        RECT 172.400 69.600 173.200 69.700 ;
        RECT 174.000 69.600 174.800 69.700 ;
        RECT 170.800 68.300 171.600 69.200 ;
        RECT 175.800 68.400 176.400 71.800 ;
        RECT 177.200 69.600 178.000 71.200 ;
        RECT 172.400 68.300 173.200 68.400 ;
        RECT 170.800 67.700 173.200 68.300 ;
        RECT 170.800 67.600 171.600 67.700 ;
        RECT 172.400 67.600 173.200 67.700 ;
        RECT 175.600 67.600 176.400 68.400 ;
        RECT 163.400 65.600 165.200 66.200 ;
        RECT 167.600 65.600 168.400 66.400 ;
        RECT 163.400 62.200 164.200 65.600 ;
        RECT 167.800 64.800 168.600 65.600 ;
        RECT 169.200 62.200 170.000 66.400 ;
        RECT 174.000 64.800 174.800 66.400 ;
        RECT 175.800 64.200 176.400 67.600 ;
        RECT 175.600 62.200 176.400 64.200 ;
        RECT 185.200 69.000 186.000 74.600 ;
        RECT 187.800 74.400 192.000 75.200 ;
        RECT 196.400 75.000 197.200 79.800 ;
        RECT 199.600 75.000 200.400 79.800 ;
        RECT 187.800 74.000 188.400 74.400 ;
        RECT 186.800 73.200 188.400 74.000 ;
        RECT 191.400 73.800 197.200 74.400 ;
        RECT 189.400 73.200 190.800 73.800 ;
        RECT 189.400 73.000 195.600 73.200 ;
        RECT 190.200 72.600 195.600 73.000 ;
        RECT 194.800 72.400 195.600 72.600 ;
        RECT 196.600 73.000 197.200 73.800 ;
        RECT 197.800 73.600 200.400 74.400 ;
        RECT 202.800 73.600 203.600 79.800 ;
        RECT 204.400 77.000 205.200 79.800 ;
        RECT 206.000 77.000 206.800 79.800 ;
        RECT 207.600 77.000 208.400 79.800 ;
        RECT 206.000 74.400 210.200 75.200 ;
        RECT 210.800 74.400 211.600 79.800 ;
        RECT 214.000 75.200 214.800 79.800 ;
        RECT 214.000 74.600 216.600 75.200 ;
        RECT 210.800 73.600 213.400 74.400 ;
        RECT 204.400 73.000 205.200 73.200 ;
        RECT 196.600 72.400 205.200 73.000 ;
        RECT 207.600 73.000 208.400 73.200 ;
        RECT 216.000 73.000 216.600 74.600 ;
        RECT 207.600 72.400 216.600 73.000 ;
        RECT 216.000 70.600 216.600 72.400 ;
        RECT 217.200 72.000 218.000 79.800 ;
        RECT 220.400 72.400 221.200 79.800 ;
        RECT 223.600 79.200 227.600 79.800 ;
        RECT 223.600 72.400 224.400 79.200 ;
        RECT 217.200 71.200 218.200 72.000 ;
        RECT 220.400 71.800 224.400 72.400 ;
        RECT 225.200 71.800 226.000 78.600 ;
        RECT 226.800 71.800 227.600 79.200 ;
        RECT 225.200 71.200 225.800 71.800 ;
        RECT 186.600 70.000 210.000 70.600 ;
        RECT 216.000 70.000 216.800 70.600 ;
        RECT 186.600 69.800 187.400 70.000 ;
        RECT 188.400 69.600 189.200 70.000 ;
        RECT 191.600 69.600 192.400 70.000 ;
        RECT 209.200 69.400 210.000 70.000 ;
        RECT 185.200 68.200 194.000 69.000 ;
        RECT 194.600 68.600 196.600 69.400 ;
        RECT 200.400 68.600 203.600 69.400 ;
        RECT 185.200 62.200 186.000 68.200 ;
        RECT 187.600 66.800 190.600 67.600 ;
        RECT 189.800 66.200 190.600 66.800 ;
        RECT 195.800 66.200 196.600 68.600 ;
        RECT 198.000 66.800 198.800 68.400 ;
        RECT 203.200 67.800 204.000 68.000 ;
        RECT 199.600 67.200 204.000 67.800 ;
        RECT 199.600 67.000 200.400 67.200 ;
        RECT 206.000 66.400 206.800 69.200 ;
        RECT 211.800 68.600 215.600 69.400 ;
        RECT 211.800 67.400 212.600 68.600 ;
        RECT 216.200 68.000 216.800 70.000 ;
        RECT 199.600 66.200 200.400 66.400 ;
        RECT 189.800 65.400 192.400 66.200 ;
        RECT 195.800 65.600 200.400 66.200 ;
        RECT 201.200 65.600 202.800 66.400 ;
        RECT 205.800 65.600 206.800 66.400 ;
        RECT 210.800 66.800 212.600 67.400 ;
        RECT 215.600 67.400 216.800 68.000 ;
        RECT 210.800 66.200 211.600 66.800 ;
        RECT 191.600 62.200 192.400 65.400 ;
        RECT 209.200 65.400 211.600 66.200 ;
        RECT 193.200 62.200 194.000 65.000 ;
        RECT 194.800 62.200 195.600 65.000 ;
        RECT 196.400 62.200 197.200 65.000 ;
        RECT 199.600 62.200 200.400 65.000 ;
        RECT 202.800 62.200 203.600 65.000 ;
        RECT 204.400 62.200 205.200 65.000 ;
        RECT 206.000 62.200 206.800 65.000 ;
        RECT 207.600 62.200 208.400 65.000 ;
        RECT 209.200 62.200 210.000 65.400 ;
        RECT 215.600 62.200 216.400 67.400 ;
        RECT 217.400 66.800 218.200 71.200 ;
        RECT 221.200 70.400 222.000 70.800 ;
        RECT 223.800 70.600 225.800 71.200 ;
        RECT 223.800 70.400 224.400 70.600 ;
        RECT 220.400 69.800 222.000 70.400 ;
        RECT 220.400 69.600 221.200 69.800 ;
        RECT 223.600 69.600 224.400 70.400 ;
        RECT 226.800 69.600 227.600 71.200 ;
        RECT 222.000 67.600 222.800 69.200 ;
        RECT 217.200 66.000 218.200 66.800 ;
        RECT 223.800 66.200 224.400 69.600 ;
        RECT 225.000 68.800 225.800 69.600 ;
        RECT 225.200 68.400 225.800 68.800 ;
        RECT 225.200 67.600 226.000 68.400 ;
        RECT 217.200 62.200 218.000 66.000 ;
        RECT 223.400 62.200 225.000 66.200 ;
        RECT 228.400 62.200 229.200 79.800 ;
        RECT 231.600 72.400 232.400 79.800 ;
        RECT 233.400 72.400 234.200 72.600 ;
        RECT 231.600 71.800 234.200 72.400 ;
        RECT 236.000 71.800 237.600 79.800 ;
        RECT 239.600 72.400 240.400 72.600 ;
        RECT 241.200 72.400 242.000 79.800 ;
        RECT 244.400 75.600 245.200 79.800 ;
        RECT 247.600 75.800 248.400 79.800 ;
        RECT 247.600 75.600 248.200 75.800 ;
        RECT 244.600 75.000 248.200 75.600 ;
        RECT 246.000 72.800 246.800 74.400 ;
        RECT 247.600 72.400 248.200 75.000 ;
        RECT 249.800 72.600 250.600 79.800 ;
        RECT 239.600 71.800 242.000 72.400 ;
        RECT 234.600 70.400 235.400 70.600 ;
        RECT 236.600 70.400 237.200 71.800 ;
        RECT 242.800 70.800 243.600 72.400 ;
        RECT 247.600 71.600 248.400 72.400 ;
        RECT 249.800 71.800 251.600 72.600 ;
        RECT 233.800 69.800 235.400 70.400 ;
        RECT 233.800 69.600 234.600 69.800 ;
        RECT 236.400 69.600 237.200 70.400 ;
        RECT 244.400 69.600 246.000 70.400 ;
        RECT 235.200 68.600 236.000 68.800 ;
        RECT 233.200 68.400 236.000 68.600 ;
        RECT 231.600 68.000 236.000 68.400 ;
        RECT 236.600 68.400 237.200 69.600 ;
        RECT 247.600 68.400 248.200 71.600 ;
        RECT 249.200 69.600 250.000 71.200 ;
        RECT 231.600 67.800 233.800 68.000 ;
        RECT 236.600 67.800 237.600 68.400 ;
        RECT 231.600 67.600 233.200 67.800 ;
        RECT 233.400 66.800 234.200 67.000 ;
        RECT 230.000 64.800 230.800 66.400 ;
        RECT 231.600 66.200 234.200 66.800 ;
        RECT 234.800 66.400 236.400 67.200 ;
        RECT 231.600 62.200 232.400 66.200 ;
        RECT 237.000 65.800 237.600 67.800 ;
        RECT 238.400 67.600 239.200 68.400 ;
        RECT 246.600 68.200 248.200 68.400 ;
        RECT 246.400 67.800 248.200 68.200 ;
        RECT 250.800 68.400 251.400 71.800 ;
        RECT 238.400 67.200 239.000 67.600 ;
        RECT 238.200 66.400 239.000 67.200 ;
        RECT 239.600 66.800 240.400 67.000 ;
        RECT 239.600 66.200 242.000 66.800 ;
        RECT 236.000 64.400 237.600 65.800 ;
        RECT 234.800 63.600 237.600 64.400 ;
        RECT 236.000 62.200 237.600 63.600 ;
        RECT 241.200 62.200 242.000 66.200 ;
        RECT 246.400 62.200 247.200 67.800 ;
        RECT 250.800 67.600 251.600 68.400 ;
        RECT 249.200 66.300 250.000 66.400 ;
        RECT 250.800 66.300 251.400 67.600 ;
        RECT 249.200 65.700 251.500 66.300 ;
        RECT 249.200 65.600 250.000 65.700 ;
        RECT 250.800 64.200 251.400 65.700 ;
        RECT 250.800 62.200 251.600 64.200 ;
        RECT 4.400 55.200 5.200 59.800 ;
        RECT 6.000 55.600 6.800 57.200 ;
        RECT 3.000 54.600 5.200 55.200 ;
        RECT 3.000 51.600 3.600 54.600 ;
        RECT 4.400 52.300 5.200 53.200 ;
        RECT 6.000 52.300 6.800 52.400 ;
        RECT 4.400 51.700 6.800 52.300 ;
        RECT 4.400 51.600 5.200 51.700 ;
        RECT 6.000 51.600 6.800 51.700 ;
        RECT 2.400 50.800 3.600 51.600 ;
        RECT 3.000 50.200 3.600 50.800 ;
        RECT 3.000 49.600 5.200 50.200 ;
        RECT 4.400 42.200 5.200 49.600 ;
        RECT 7.600 42.200 8.400 59.800 ;
        RECT 9.200 56.300 10.000 56.400 ;
        RECT 10.800 56.300 11.600 59.800 ;
        RECT 9.200 55.700 11.600 56.300 ;
        RECT 9.200 55.600 10.000 55.700 ;
        RECT 10.600 55.200 11.600 55.700 ;
        RECT 10.600 50.800 11.400 55.200 ;
        RECT 12.400 54.600 13.200 59.800 ;
        RECT 18.800 56.600 19.600 59.800 ;
        RECT 20.400 57.000 21.200 59.800 ;
        RECT 22.000 57.000 22.800 59.800 ;
        RECT 23.600 57.000 24.400 59.800 ;
        RECT 25.200 57.000 26.000 59.800 ;
        RECT 28.400 57.000 29.200 59.800 ;
        RECT 31.600 57.000 32.400 59.800 ;
        RECT 33.200 57.000 34.000 59.800 ;
        RECT 34.800 57.000 35.600 59.800 ;
        RECT 17.200 55.800 19.600 56.600 ;
        RECT 36.400 56.600 37.200 59.800 ;
        RECT 17.200 55.200 18.000 55.800 ;
        RECT 12.000 54.000 13.200 54.600 ;
        RECT 16.200 54.600 18.000 55.200 ;
        RECT 22.000 55.600 23.000 56.400 ;
        RECT 26.000 55.600 27.600 56.400 ;
        RECT 28.400 55.800 33.000 56.400 ;
        RECT 36.400 55.800 39.000 56.600 ;
        RECT 28.400 55.600 29.200 55.800 ;
        RECT 12.000 52.000 12.600 54.000 ;
        RECT 16.200 53.400 17.000 54.600 ;
        RECT 13.200 52.600 17.000 53.400 ;
        RECT 22.000 52.800 22.800 55.600 ;
        RECT 28.400 54.800 29.200 55.000 ;
        RECT 24.800 54.200 29.200 54.800 ;
        RECT 24.800 54.000 25.600 54.200 ;
        RECT 30.000 53.600 30.800 55.200 ;
        RECT 32.200 53.400 33.000 55.800 ;
        RECT 38.200 55.200 39.000 55.800 ;
        RECT 38.200 54.400 41.200 55.200 ;
        RECT 42.800 53.800 43.600 59.800 ;
        RECT 46.000 56.000 46.800 59.800 ;
        RECT 25.200 52.600 28.400 53.400 ;
        RECT 32.200 52.600 34.200 53.400 ;
        RECT 34.800 53.000 43.600 53.800 ;
        RECT 18.800 52.000 19.600 52.600 ;
        RECT 36.400 52.000 37.200 52.400 ;
        RECT 38.000 52.000 38.800 52.400 ;
        RECT 39.600 52.000 40.400 52.400 ;
        RECT 41.400 52.000 42.200 52.200 ;
        RECT 12.000 51.400 12.800 52.000 ;
        RECT 18.800 51.400 42.200 52.000 ;
        RECT 10.600 50.000 11.600 50.800 ;
        RECT 10.800 42.200 11.600 50.000 ;
        RECT 12.200 49.600 12.800 51.400 ;
        RECT 12.200 49.000 21.200 49.600 ;
        RECT 12.200 47.400 12.800 49.000 ;
        RECT 20.400 48.800 21.200 49.000 ;
        RECT 23.600 49.000 32.200 49.600 ;
        RECT 23.600 48.800 24.400 49.000 ;
        RECT 15.400 47.600 18.000 48.400 ;
        RECT 12.200 46.800 14.800 47.400 ;
        RECT 14.000 42.200 14.800 46.800 ;
        RECT 17.200 42.200 18.000 47.600 ;
        RECT 18.600 46.800 22.800 47.600 ;
        RECT 20.400 42.200 21.200 45.000 ;
        RECT 22.000 42.200 22.800 45.000 ;
        RECT 23.600 42.200 24.400 45.000 ;
        RECT 25.200 42.200 26.000 48.400 ;
        RECT 28.400 47.600 31.000 48.400 ;
        RECT 31.600 48.200 32.200 49.000 ;
        RECT 33.200 49.400 34.000 49.600 ;
        RECT 33.200 49.000 38.600 49.400 ;
        RECT 33.200 48.800 39.400 49.000 ;
        RECT 38.000 48.200 39.400 48.800 ;
        RECT 31.600 47.600 37.400 48.200 ;
        RECT 40.400 48.000 42.000 48.800 ;
        RECT 40.400 47.600 41.000 48.000 ;
        RECT 28.400 42.200 29.200 47.000 ;
        RECT 31.600 42.200 32.400 47.000 ;
        RECT 36.800 46.800 41.000 47.600 ;
        RECT 42.800 47.400 43.600 53.000 ;
        RECT 45.800 55.200 46.800 56.000 ;
        RECT 45.800 50.800 46.600 55.200 ;
        RECT 47.600 54.600 48.400 59.800 ;
        RECT 54.000 56.600 54.800 59.800 ;
        RECT 55.600 57.000 56.400 59.800 ;
        RECT 57.200 57.000 58.000 59.800 ;
        RECT 58.800 57.000 59.600 59.800 ;
        RECT 60.400 57.000 61.200 59.800 ;
        RECT 63.600 57.000 64.400 59.800 ;
        RECT 66.800 57.000 67.600 59.800 ;
        RECT 68.400 57.000 69.200 59.800 ;
        RECT 70.000 57.000 70.800 59.800 ;
        RECT 52.400 55.800 54.800 56.600 ;
        RECT 71.600 56.600 72.400 59.800 ;
        RECT 52.400 55.200 53.200 55.800 ;
        RECT 47.200 54.000 48.400 54.600 ;
        RECT 51.400 54.600 53.200 55.200 ;
        RECT 57.200 55.600 58.200 56.400 ;
        RECT 61.200 55.600 62.800 56.400 ;
        RECT 63.600 55.800 68.200 56.400 ;
        RECT 71.600 55.800 74.200 56.600 ;
        RECT 63.600 55.600 64.400 55.800 ;
        RECT 47.200 52.000 47.800 54.000 ;
        RECT 51.400 53.400 52.200 54.600 ;
        RECT 48.400 52.600 52.200 53.400 ;
        RECT 57.200 52.800 58.000 55.600 ;
        RECT 63.600 54.800 64.400 55.000 ;
        RECT 60.000 54.200 64.400 54.800 ;
        RECT 60.000 54.000 60.800 54.200 ;
        RECT 65.200 53.600 66.000 55.200 ;
        RECT 67.400 53.400 68.200 55.800 ;
        RECT 73.400 55.200 74.200 55.800 ;
        RECT 73.400 54.400 76.400 55.200 ;
        RECT 78.000 53.800 78.800 59.800 ;
        RECT 60.400 52.600 63.600 53.400 ;
        RECT 67.400 52.600 69.400 53.400 ;
        RECT 70.000 53.000 78.800 53.800 ;
        RECT 79.600 54.300 80.400 54.400 ;
        RECT 86.000 54.300 86.800 59.800 ;
        RECT 89.200 55.200 90.000 59.800 ;
        RECT 79.600 53.700 86.800 54.300 ;
        RECT 79.600 53.600 80.400 53.700 ;
        RECT 54.000 52.000 54.800 52.600 ;
        RECT 71.600 52.000 72.400 52.400 ;
        RECT 74.800 52.000 75.600 52.400 ;
        RECT 76.600 52.000 77.400 52.200 ;
        RECT 47.200 51.400 48.000 52.000 ;
        RECT 54.000 51.400 77.400 52.000 ;
        RECT 45.800 50.000 46.800 50.800 ;
        RECT 41.600 46.800 43.600 47.400 ;
        RECT 33.200 42.200 34.000 45.000 ;
        RECT 34.800 42.200 35.600 45.000 ;
        RECT 38.000 42.200 38.800 46.800 ;
        RECT 41.600 46.200 42.200 46.800 ;
        RECT 41.200 45.600 42.200 46.200 ;
        RECT 41.200 42.200 42.000 45.600 ;
        RECT 46.000 42.200 46.800 50.000 ;
        RECT 47.400 49.600 48.000 51.400 ;
        RECT 47.400 49.000 56.400 49.600 ;
        RECT 47.400 47.400 48.000 49.000 ;
        RECT 55.600 48.800 56.400 49.000 ;
        RECT 58.800 49.000 67.400 49.600 ;
        RECT 58.800 48.800 59.600 49.000 ;
        RECT 50.600 47.600 53.200 48.400 ;
        RECT 47.400 46.800 50.000 47.400 ;
        RECT 49.200 42.200 50.000 46.800 ;
        RECT 52.400 42.200 53.200 47.600 ;
        RECT 53.800 46.800 58.000 47.600 ;
        RECT 55.600 42.200 56.400 45.000 ;
        RECT 57.200 42.200 58.000 45.000 ;
        RECT 58.800 42.200 59.600 45.000 ;
        RECT 60.400 42.200 61.200 48.400 ;
        RECT 63.600 47.600 66.200 48.400 ;
        RECT 66.800 48.200 67.400 49.000 ;
        RECT 68.400 49.400 69.200 49.600 ;
        RECT 68.400 49.000 73.800 49.400 ;
        RECT 68.400 48.800 74.600 49.000 ;
        RECT 73.200 48.200 74.600 48.800 ;
        RECT 66.800 47.600 72.600 48.200 ;
        RECT 75.600 48.000 77.200 48.800 ;
        RECT 75.600 47.600 76.200 48.000 ;
        RECT 63.600 42.200 64.400 47.000 ;
        RECT 66.800 42.200 67.600 47.000 ;
        RECT 72.000 46.800 76.200 47.600 ;
        RECT 78.000 47.400 78.800 53.000 ;
        RECT 76.800 46.800 78.800 47.400 ;
        RECT 86.000 52.400 86.800 53.700 ;
        RECT 87.800 54.600 90.000 55.200 ;
        RECT 86.000 50.200 86.600 52.400 ;
        RECT 87.800 51.600 88.400 54.600 ;
        RECT 89.200 51.600 90.000 53.200 ;
        RECT 90.800 52.400 91.600 59.800 ;
        RECT 94.000 55.200 94.800 59.800 ;
        RECT 92.600 54.600 94.800 55.200 ;
        RECT 95.600 55.200 96.400 59.800 ;
        RECT 95.600 54.600 97.800 55.200 ;
        RECT 87.200 50.800 88.400 51.600 ;
        RECT 87.800 50.200 88.400 50.800 ;
        RECT 90.800 50.200 91.400 52.400 ;
        RECT 92.600 51.600 93.200 54.600 ;
        RECT 94.000 51.600 94.800 53.200 ;
        RECT 95.600 51.600 96.400 53.200 ;
        RECT 97.200 51.600 97.800 54.600 ;
        RECT 98.800 52.400 99.600 59.800 ;
        RECT 102.000 57.800 102.800 59.800 ;
        RECT 102.000 54.400 102.600 57.800 ;
        RECT 103.600 55.600 104.400 57.200 ;
        RECT 102.000 53.600 102.800 54.400 ;
        RECT 105.200 53.800 106.000 59.800 ;
        RECT 111.600 56.600 112.400 59.800 ;
        RECT 113.200 57.000 114.000 59.800 ;
        RECT 114.800 57.000 115.600 59.800 ;
        RECT 116.400 57.000 117.200 59.800 ;
        RECT 119.600 57.000 120.400 59.800 ;
        RECT 122.800 57.000 123.600 59.800 ;
        RECT 124.400 57.000 125.200 59.800 ;
        RECT 126.000 57.000 126.800 59.800 ;
        RECT 127.600 57.000 128.400 59.800 ;
        RECT 109.800 55.800 112.400 56.600 ;
        RECT 129.200 56.600 130.000 59.800 ;
        RECT 115.800 55.800 120.400 56.400 ;
        RECT 109.800 55.200 110.600 55.800 ;
        RECT 107.600 54.400 110.600 55.200 ;
        RECT 92.000 50.800 93.200 51.600 ;
        RECT 92.600 50.200 93.200 50.800 ;
        RECT 97.200 50.800 98.400 51.600 ;
        RECT 97.200 50.200 97.800 50.800 ;
        RECT 99.000 50.200 99.600 52.400 ;
        RECT 100.400 50.800 101.200 52.400 ;
        RECT 102.000 50.200 102.600 53.600 ;
        RECT 105.200 53.000 114.000 53.800 ;
        RECT 115.800 53.400 116.600 55.800 ;
        RECT 119.600 55.600 120.400 55.800 ;
        RECT 121.200 55.600 122.800 56.400 ;
        RECT 125.800 55.600 126.800 56.400 ;
        RECT 129.200 55.800 131.600 56.600 ;
        RECT 118.000 53.600 118.800 55.200 ;
        RECT 119.600 54.800 120.400 55.000 ;
        RECT 119.600 54.200 124.000 54.800 ;
        RECT 123.200 54.000 124.000 54.200 ;
        RECT 68.400 42.200 69.200 45.000 ;
        RECT 70.000 42.200 70.800 45.000 ;
        RECT 73.200 42.200 74.000 46.800 ;
        RECT 76.800 46.200 77.400 46.800 ;
        RECT 76.400 45.600 77.400 46.200 ;
        RECT 76.400 42.200 77.200 45.600 ;
        RECT 86.000 42.200 86.800 50.200 ;
        RECT 87.800 49.600 90.000 50.200 ;
        RECT 89.200 42.200 90.000 49.600 ;
        RECT 90.800 42.200 91.600 50.200 ;
        RECT 92.600 49.600 94.800 50.200 ;
        RECT 94.000 42.200 94.800 49.600 ;
        RECT 95.600 49.600 97.800 50.200 ;
        RECT 95.600 42.200 96.400 49.600 ;
        RECT 98.800 42.200 99.600 50.200 ;
        RECT 101.000 49.400 102.800 50.200 ;
        RECT 101.000 42.200 101.800 49.400 ;
        RECT 105.200 47.400 106.000 53.000 ;
        RECT 114.600 52.600 116.600 53.400 ;
        RECT 120.400 52.600 123.600 53.400 ;
        RECT 126.000 52.800 126.800 55.600 ;
        RECT 130.800 55.200 131.600 55.800 ;
        RECT 130.800 54.600 132.600 55.200 ;
        RECT 131.800 53.400 132.600 54.600 ;
        RECT 135.600 54.600 136.400 59.800 ;
        RECT 137.200 56.000 138.000 59.800 ;
        RECT 137.200 55.200 138.200 56.000 ;
        RECT 135.600 54.000 136.800 54.600 ;
        RECT 131.800 52.600 135.600 53.400 ;
        RECT 106.600 52.000 107.400 52.200 ;
        RECT 108.400 52.000 109.200 52.400 ;
        RECT 111.600 52.000 112.400 52.400 ;
        RECT 129.200 52.000 130.000 52.600 ;
        RECT 136.200 52.000 136.800 54.000 ;
        RECT 106.600 51.400 130.000 52.000 ;
        RECT 136.000 51.400 136.800 52.000 ;
        RECT 136.000 49.600 136.600 51.400 ;
        RECT 137.400 50.800 138.200 55.200 ;
        RECT 138.800 54.300 139.600 54.400 ;
        RECT 140.400 54.300 141.200 59.800 ;
        RECT 144.200 58.400 145.000 59.800 ;
        RECT 143.600 57.600 145.000 58.400 ;
        RECT 142.000 55.600 142.800 57.200 ;
        RECT 144.200 56.400 145.000 57.600 ;
        RECT 144.200 55.800 146.000 56.400 ;
        RECT 138.800 53.700 141.200 54.300 ;
        RECT 138.800 53.600 139.600 53.700 ;
        RECT 114.800 49.400 115.600 49.600 ;
        RECT 110.200 49.000 115.600 49.400 ;
        RECT 109.400 48.800 115.600 49.000 ;
        RECT 116.600 49.000 125.200 49.600 ;
        RECT 106.800 48.000 108.400 48.800 ;
        RECT 109.400 48.200 110.800 48.800 ;
        RECT 116.600 48.200 117.200 49.000 ;
        RECT 124.400 48.800 125.200 49.000 ;
        RECT 127.600 49.000 136.600 49.600 ;
        RECT 127.600 48.800 128.400 49.000 ;
        RECT 107.800 47.600 108.400 48.000 ;
        RECT 111.400 47.600 117.200 48.200 ;
        RECT 117.800 47.600 120.400 48.400 ;
        RECT 105.200 46.800 107.200 47.400 ;
        RECT 107.800 46.800 112.000 47.600 ;
        RECT 106.600 46.200 107.200 46.800 ;
        RECT 106.600 45.600 107.600 46.200 ;
        RECT 106.800 42.200 107.600 45.600 ;
        RECT 110.000 42.200 110.800 46.800 ;
        RECT 113.200 42.200 114.000 45.000 ;
        RECT 114.800 42.200 115.600 45.000 ;
        RECT 116.400 42.200 117.200 47.000 ;
        RECT 119.600 42.200 120.400 47.000 ;
        RECT 122.800 42.200 123.600 48.400 ;
        RECT 130.800 47.600 133.400 48.400 ;
        RECT 126.000 46.800 130.200 47.600 ;
        RECT 124.400 42.200 125.200 45.000 ;
        RECT 126.000 42.200 126.800 45.000 ;
        RECT 127.600 42.200 128.400 45.000 ;
        RECT 130.800 42.200 131.600 47.600 ;
        RECT 136.000 47.400 136.600 49.000 ;
        RECT 134.000 46.800 136.600 47.400 ;
        RECT 137.200 50.000 138.200 50.800 ;
        RECT 140.400 50.300 141.200 53.700 ;
        RECT 143.600 50.300 144.400 50.400 ;
        RECT 134.000 42.200 134.800 46.800 ;
        RECT 137.200 42.200 138.000 50.000 ;
        RECT 140.400 49.700 144.400 50.300 ;
        RECT 140.400 42.200 141.200 49.700 ;
        RECT 143.600 48.800 144.400 49.700 ;
        RECT 145.200 42.200 146.000 55.800 ;
        RECT 148.400 55.600 149.200 57.200 ;
        RECT 150.000 56.300 150.800 59.800 ;
        RECT 151.600 56.300 152.400 56.400 ;
        RECT 150.000 55.700 152.400 56.300 ;
        RECT 153.200 56.000 154.000 59.800 ;
        RECT 146.800 54.300 147.600 55.200 ;
        RECT 148.400 54.300 149.200 54.400 ;
        RECT 146.800 53.700 149.200 54.300 ;
        RECT 146.800 53.600 147.600 53.700 ;
        RECT 148.400 53.600 149.200 53.700 ;
        RECT 150.000 42.200 150.800 55.700 ;
        RECT 151.600 55.600 152.400 55.700 ;
        RECT 153.000 55.200 154.000 56.000 ;
        RECT 153.000 50.800 153.800 55.200 ;
        RECT 154.800 54.600 155.600 59.800 ;
        RECT 161.200 56.600 162.000 59.800 ;
        RECT 162.800 57.000 163.600 59.800 ;
        RECT 164.400 57.000 165.200 59.800 ;
        RECT 166.000 57.000 166.800 59.800 ;
        RECT 167.600 57.000 168.400 59.800 ;
        RECT 170.800 57.000 171.600 59.800 ;
        RECT 174.000 57.000 174.800 59.800 ;
        RECT 175.600 57.000 176.400 59.800 ;
        RECT 177.200 57.000 178.000 59.800 ;
        RECT 159.600 55.800 162.000 56.600 ;
        RECT 178.800 56.600 179.600 59.800 ;
        RECT 159.600 55.200 160.400 55.800 ;
        RECT 154.400 54.000 155.600 54.600 ;
        RECT 158.600 54.600 160.400 55.200 ;
        RECT 164.400 55.600 165.400 56.400 ;
        RECT 168.400 55.600 170.000 56.400 ;
        RECT 170.800 55.800 175.400 56.400 ;
        RECT 178.800 55.800 181.400 56.600 ;
        RECT 170.800 55.600 171.600 55.800 ;
        RECT 154.400 52.000 155.000 54.000 ;
        RECT 158.600 53.400 159.400 54.600 ;
        RECT 155.600 52.600 159.400 53.400 ;
        RECT 164.400 52.800 165.200 55.600 ;
        RECT 170.800 54.800 171.600 55.000 ;
        RECT 167.200 54.200 171.600 54.800 ;
        RECT 167.200 54.000 168.000 54.200 ;
        RECT 172.400 53.600 173.200 55.200 ;
        RECT 174.600 53.400 175.400 55.800 ;
        RECT 180.600 55.200 181.400 55.800 ;
        RECT 180.600 54.400 183.600 55.200 ;
        RECT 185.200 53.800 186.000 59.800 ;
        RECT 195.800 56.400 196.600 59.800 ;
        RECT 194.800 55.800 196.600 56.400 ;
        RECT 167.600 52.600 170.800 53.400 ;
        RECT 174.600 52.600 176.600 53.400 ;
        RECT 177.200 53.000 186.000 53.800 ;
        RECT 193.200 53.600 194.000 55.200 ;
        RECT 161.200 52.000 162.000 52.600 ;
        RECT 172.400 52.000 173.200 52.400 ;
        RECT 178.800 52.000 179.600 52.400 ;
        RECT 183.800 52.000 184.600 52.200 ;
        RECT 154.400 51.400 155.200 52.000 ;
        RECT 161.200 51.400 184.600 52.000 ;
        RECT 153.000 50.000 154.000 50.800 ;
        RECT 153.200 42.200 154.000 50.000 ;
        RECT 154.600 49.600 155.200 51.400 ;
        RECT 154.600 49.000 163.600 49.600 ;
        RECT 154.600 47.400 155.200 49.000 ;
        RECT 162.800 48.800 163.600 49.000 ;
        RECT 166.000 49.000 174.600 49.600 ;
        RECT 166.000 48.800 166.800 49.000 ;
        RECT 157.800 47.600 160.400 48.400 ;
        RECT 154.600 46.800 157.200 47.400 ;
        RECT 156.400 42.200 157.200 46.800 ;
        RECT 159.600 42.200 160.400 47.600 ;
        RECT 161.000 46.800 165.200 47.600 ;
        RECT 162.800 42.200 163.600 45.000 ;
        RECT 164.400 42.200 165.200 45.000 ;
        RECT 166.000 42.200 166.800 45.000 ;
        RECT 167.600 42.200 168.400 48.400 ;
        RECT 170.800 47.600 173.400 48.400 ;
        RECT 174.000 48.200 174.600 49.000 ;
        RECT 175.600 49.400 176.400 49.600 ;
        RECT 175.600 49.000 181.000 49.400 ;
        RECT 175.600 48.800 181.800 49.000 ;
        RECT 180.400 48.200 181.800 48.800 ;
        RECT 174.000 47.600 179.800 48.200 ;
        RECT 182.800 48.000 184.400 48.800 ;
        RECT 182.800 47.600 183.400 48.000 ;
        RECT 170.800 42.200 171.600 47.000 ;
        RECT 174.000 42.200 174.800 47.000 ;
        RECT 179.200 46.800 183.400 47.600 ;
        RECT 185.200 47.400 186.000 53.000 ;
        RECT 184.000 46.800 186.000 47.400 ;
        RECT 194.800 52.300 195.600 55.800 ;
        RECT 196.400 54.300 197.200 54.400 ;
        RECT 199.200 54.300 200.000 59.800 ;
        RECT 207.000 56.400 207.800 59.800 ;
        RECT 206.000 55.800 207.800 56.400 ;
        RECT 196.400 53.800 200.000 54.300 ;
        RECT 196.400 53.700 199.800 53.800 ;
        RECT 196.400 53.600 197.200 53.700 ;
        RECT 198.200 53.600 199.800 53.700 ;
        RECT 204.400 53.600 205.200 55.200 ;
        RECT 196.400 52.300 197.200 52.400 ;
        RECT 194.800 51.700 197.200 52.300 ;
        RECT 175.600 42.200 176.400 45.000 ;
        RECT 177.200 42.200 178.000 45.000 ;
        RECT 180.400 42.200 181.200 46.800 ;
        RECT 184.000 46.200 184.600 46.800 ;
        RECT 183.600 45.600 184.600 46.200 ;
        RECT 183.600 42.200 184.400 45.600 ;
        RECT 194.800 42.200 195.600 51.700 ;
        RECT 196.400 51.600 197.200 51.700 ;
        RECT 198.200 50.400 198.800 53.600 ;
        RECT 200.400 51.600 202.000 52.400 ;
        RECT 196.400 48.800 197.200 50.400 ;
        RECT 198.000 49.600 198.800 50.400 ;
        RECT 202.800 50.300 203.600 51.200 ;
        RECT 206.000 50.300 206.800 55.800 ;
        RECT 209.200 53.800 210.000 59.800 ;
        RECT 215.600 56.600 216.400 59.800 ;
        RECT 217.200 57.000 218.000 59.800 ;
        RECT 218.800 57.000 219.600 59.800 ;
        RECT 220.400 57.000 221.200 59.800 ;
        RECT 223.600 57.000 224.400 59.800 ;
        RECT 226.800 57.000 227.600 59.800 ;
        RECT 228.400 57.000 229.200 59.800 ;
        RECT 230.000 57.000 230.800 59.800 ;
        RECT 231.600 57.000 232.400 59.800 ;
        RECT 213.800 55.800 216.400 56.600 ;
        RECT 233.200 56.600 234.000 59.800 ;
        RECT 219.800 55.800 224.400 56.400 ;
        RECT 213.800 55.200 214.600 55.800 ;
        RECT 211.600 54.400 214.600 55.200 ;
        RECT 209.200 53.000 218.000 53.800 ;
        RECT 219.800 53.400 220.600 55.800 ;
        RECT 223.600 55.600 224.400 55.800 ;
        RECT 225.200 55.600 226.800 56.400 ;
        RECT 229.800 55.600 230.800 56.400 ;
        RECT 233.200 55.800 235.600 56.600 ;
        RECT 222.000 53.600 222.800 55.200 ;
        RECT 223.600 54.800 224.400 55.000 ;
        RECT 223.600 54.200 228.000 54.800 ;
        RECT 227.200 54.000 228.000 54.200 ;
        RECT 202.800 49.700 206.800 50.300 ;
        RECT 202.800 49.600 203.600 49.700 ;
        RECT 198.200 47.000 198.800 49.600 ;
        RECT 199.600 47.600 200.400 49.200 ;
        RECT 198.200 46.400 201.800 47.000 ;
        RECT 198.200 46.200 198.800 46.400 ;
        RECT 198.000 42.200 198.800 46.200 ;
        RECT 201.200 46.200 201.800 46.400 ;
        RECT 201.200 42.200 202.000 46.200 ;
        RECT 206.000 42.200 206.800 49.700 ;
        RECT 207.600 48.800 208.400 50.400 ;
        RECT 209.200 47.400 210.000 53.000 ;
        RECT 218.600 52.600 220.600 53.400 ;
        RECT 224.400 52.600 227.600 53.400 ;
        RECT 230.000 52.800 230.800 55.600 ;
        RECT 234.800 55.200 235.600 55.800 ;
        RECT 234.800 54.600 236.600 55.200 ;
        RECT 235.800 53.400 236.600 54.600 ;
        RECT 239.600 54.600 240.400 59.800 ;
        RECT 241.200 56.000 242.000 59.800 ;
        RECT 241.200 55.200 242.200 56.000 ;
        RECT 239.600 54.000 240.800 54.600 ;
        RECT 235.800 52.600 239.600 53.400 ;
        RECT 210.600 52.000 211.400 52.200 ;
        RECT 214.000 52.000 214.800 52.400 ;
        RECT 215.600 52.000 216.400 52.400 ;
        RECT 233.200 52.000 234.000 52.600 ;
        RECT 240.200 52.000 240.800 54.000 ;
        RECT 210.600 51.400 234.000 52.000 ;
        RECT 240.000 51.400 240.800 52.000 ;
        RECT 241.400 52.300 242.200 55.200 ;
        RECT 244.400 55.200 245.200 59.800 ;
        RECT 249.800 58.400 250.600 59.800 ;
        RECT 249.800 57.600 251.600 58.400 ;
        RECT 249.800 56.400 250.600 57.600 ;
        RECT 249.800 55.800 251.600 56.400 ;
        RECT 244.400 54.600 246.600 55.200 ;
        RECT 244.400 52.300 245.200 53.200 ;
        RECT 241.400 51.700 245.200 52.300 ;
        RECT 240.000 49.600 240.600 51.400 ;
        RECT 241.400 50.800 242.200 51.700 ;
        RECT 244.400 51.600 245.200 51.700 ;
        RECT 246.000 51.600 246.600 54.600 ;
        RECT 218.800 49.400 219.600 49.600 ;
        RECT 214.200 49.000 219.600 49.400 ;
        RECT 213.400 48.800 219.600 49.000 ;
        RECT 220.600 49.000 229.200 49.600 ;
        RECT 210.800 48.000 212.400 48.800 ;
        RECT 213.400 48.200 214.800 48.800 ;
        RECT 220.600 48.200 221.200 49.000 ;
        RECT 228.400 48.800 229.200 49.000 ;
        RECT 231.600 49.000 240.600 49.600 ;
        RECT 231.600 48.800 232.400 49.000 ;
        RECT 211.800 47.600 212.400 48.000 ;
        RECT 215.400 47.600 221.200 48.200 ;
        RECT 221.800 47.600 224.400 48.400 ;
        RECT 209.200 46.800 211.200 47.400 ;
        RECT 211.800 46.800 216.000 47.600 ;
        RECT 210.600 46.200 211.200 46.800 ;
        RECT 210.600 45.600 211.600 46.200 ;
        RECT 210.800 42.200 211.600 45.600 ;
        RECT 214.000 42.200 214.800 46.800 ;
        RECT 217.200 42.200 218.000 45.000 ;
        RECT 218.800 42.200 219.600 45.000 ;
        RECT 220.400 42.200 221.200 47.000 ;
        RECT 223.600 42.200 224.400 47.000 ;
        RECT 226.800 42.200 227.600 48.400 ;
        RECT 234.800 47.600 237.400 48.400 ;
        RECT 230.000 46.800 234.200 47.600 ;
        RECT 228.400 42.200 229.200 45.000 ;
        RECT 230.000 42.200 230.800 45.000 ;
        RECT 231.600 42.200 232.400 45.000 ;
        RECT 234.800 42.200 235.600 47.600 ;
        RECT 240.000 47.400 240.600 49.000 ;
        RECT 238.000 46.800 240.600 47.400 ;
        RECT 241.200 50.000 242.200 50.800 ;
        RECT 246.000 50.800 247.200 51.600 ;
        RECT 246.000 50.200 246.600 50.800 ;
        RECT 238.000 42.200 238.800 46.800 ;
        RECT 241.200 42.200 242.000 50.000 ;
        RECT 244.400 49.600 246.600 50.200 ;
        RECT 244.400 42.200 245.200 49.600 ;
        RECT 249.200 48.800 250.000 50.400 ;
        RECT 250.800 42.200 251.600 55.800 ;
        RECT 252.400 53.600 253.200 55.200 ;
        RECT 4.400 32.400 5.200 39.800 ;
        RECT 3.000 31.800 5.200 32.400 ;
        RECT 7.600 32.000 8.400 39.800 ;
        RECT 10.800 35.200 11.600 39.800 ;
        RECT 3.000 31.200 3.600 31.800 ;
        RECT 2.400 30.400 3.600 31.200 ;
        RECT 7.400 31.200 8.400 32.000 ;
        RECT 9.000 34.600 11.600 35.200 ;
        RECT 9.000 33.000 9.600 34.600 ;
        RECT 14.000 34.400 14.800 39.800 ;
        RECT 17.200 37.000 18.000 39.800 ;
        RECT 18.800 37.000 19.600 39.800 ;
        RECT 20.400 37.000 21.200 39.800 ;
        RECT 15.400 34.400 19.600 35.200 ;
        RECT 12.200 33.600 14.800 34.400 ;
        RECT 22.000 33.600 22.800 39.800 ;
        RECT 25.200 35.000 26.000 39.800 ;
        RECT 28.400 35.000 29.200 39.800 ;
        RECT 30.000 37.000 30.800 39.800 ;
        RECT 31.600 37.000 32.400 39.800 ;
        RECT 34.800 35.200 35.600 39.800 ;
        RECT 38.000 36.400 38.800 39.800 ;
        RECT 38.000 35.800 39.000 36.400 ;
        RECT 38.400 35.200 39.000 35.800 ;
        RECT 33.600 34.400 37.800 35.200 ;
        RECT 38.400 34.600 40.400 35.200 ;
        RECT 25.200 33.600 27.800 34.400 ;
        RECT 28.400 33.800 34.200 34.400 ;
        RECT 37.200 34.000 37.800 34.400 ;
        RECT 17.200 33.000 18.000 33.200 ;
        RECT 9.000 32.400 18.000 33.000 ;
        RECT 20.400 33.000 21.200 33.200 ;
        RECT 28.400 33.000 29.000 33.800 ;
        RECT 34.800 33.200 36.200 33.800 ;
        RECT 37.200 33.200 38.800 34.000 ;
        RECT 20.400 32.400 29.000 33.000 ;
        RECT 30.000 33.000 36.200 33.200 ;
        RECT 30.000 32.600 35.400 33.000 ;
        RECT 30.000 32.400 30.800 32.600 ;
        RECT 3.000 27.400 3.600 30.400 ;
        RECT 4.400 30.300 5.200 30.400 ;
        RECT 7.400 30.300 8.200 31.200 ;
        RECT 9.000 30.600 9.600 32.400 ;
        RECT 4.400 29.700 8.200 30.300 ;
        RECT 4.400 28.800 5.200 29.700 ;
        RECT 3.000 26.800 5.200 27.400 ;
        RECT 4.400 22.200 5.200 26.800 ;
        RECT 7.400 26.800 8.200 29.700 ;
        RECT 8.800 30.000 9.600 30.600 ;
        RECT 15.600 30.000 39.000 30.600 ;
        RECT 8.800 28.000 9.400 30.000 ;
        RECT 15.600 29.400 16.400 30.000 ;
        RECT 33.200 29.600 34.000 30.000 ;
        RECT 36.400 29.600 37.200 30.000 ;
        RECT 38.200 29.800 39.000 30.000 ;
        RECT 10.000 28.600 13.800 29.400 ;
        RECT 8.800 27.400 10.000 28.000 ;
        RECT 7.400 26.000 8.400 26.800 ;
        RECT 7.600 22.200 8.400 26.000 ;
        RECT 9.200 22.200 10.000 27.400 ;
        RECT 13.000 27.400 13.800 28.600 ;
        RECT 13.000 26.800 14.800 27.400 ;
        RECT 14.000 26.200 14.800 26.800 ;
        RECT 18.800 26.400 19.600 29.200 ;
        RECT 22.000 28.600 25.200 29.400 ;
        RECT 29.000 28.600 31.000 29.400 ;
        RECT 39.600 29.000 40.400 34.600 ;
        RECT 41.200 31.800 42.000 39.800 ;
        RECT 42.800 32.400 43.600 39.800 ;
        RECT 46.000 32.400 46.800 39.800 ;
        RECT 50.200 32.600 51.000 39.800 ;
        RECT 42.800 31.800 46.800 32.400 ;
        RECT 49.200 31.800 51.000 32.600 ;
        RECT 52.400 31.800 53.200 39.800 ;
        RECT 55.600 32.400 56.400 39.800 ;
        RECT 65.200 36.400 66.000 39.800 ;
        RECT 65.000 35.800 66.000 36.400 ;
        RECT 65.000 35.200 65.600 35.800 ;
        RECT 68.400 35.200 69.200 39.800 ;
        RECT 71.600 37.000 72.400 39.800 ;
        RECT 73.200 37.000 74.000 39.800 ;
        RECT 54.200 31.800 56.400 32.400 ;
        RECT 63.600 34.600 65.600 35.200 ;
        RECT 41.400 30.400 42.000 31.800 ;
        RECT 45.200 30.400 46.000 30.800 ;
        RECT 41.200 29.800 43.600 30.400 ;
        RECT 45.200 29.800 46.800 30.400 ;
        RECT 41.200 29.600 42.000 29.800 ;
        RECT 21.600 27.800 22.400 28.000 ;
        RECT 21.600 27.200 26.000 27.800 ;
        RECT 25.200 27.000 26.000 27.200 ;
        RECT 26.800 26.800 27.600 28.400 ;
        RECT 14.000 25.400 16.400 26.200 ;
        RECT 18.800 25.600 19.800 26.400 ;
        RECT 22.800 25.600 24.400 26.400 ;
        RECT 25.200 26.200 26.000 26.400 ;
        RECT 29.000 26.200 29.800 28.600 ;
        RECT 31.600 28.200 40.400 29.000 ;
        RECT 43.000 28.400 43.600 29.800 ;
        RECT 46.000 29.600 46.800 29.800 ;
        RECT 47.600 30.300 48.400 30.400 ;
        RECT 49.400 30.300 50.000 31.800 ;
        RECT 47.600 29.700 50.000 30.300 ;
        RECT 47.600 29.600 48.400 29.700 ;
        RECT 35.000 26.800 38.000 27.600 ;
        RECT 35.000 26.200 35.800 26.800 ;
        RECT 25.200 25.600 29.800 26.200 ;
        RECT 15.600 22.200 16.400 25.400 ;
        RECT 33.200 25.400 35.800 26.200 ;
        RECT 17.200 22.200 18.000 25.000 ;
        RECT 18.800 22.200 19.600 25.000 ;
        RECT 20.400 22.200 21.200 25.000 ;
        RECT 22.000 22.200 22.800 25.000 ;
        RECT 25.200 22.200 26.000 25.000 ;
        RECT 28.400 22.200 29.200 25.000 ;
        RECT 30.000 22.200 30.800 25.000 ;
        RECT 31.600 22.200 32.400 25.000 ;
        RECT 33.200 22.200 34.000 25.400 ;
        RECT 39.600 22.200 40.400 28.200 ;
        RECT 42.800 27.600 43.600 28.400 ;
        RECT 44.400 27.600 45.200 29.200 ;
        RECT 49.400 28.400 50.000 29.700 ;
        RECT 50.800 29.600 51.600 31.200 ;
        RECT 52.400 29.600 53.000 31.800 ;
        RECT 54.200 31.200 54.800 31.800 ;
        RECT 53.600 30.400 54.800 31.200 ;
        RECT 49.200 27.600 50.000 28.400 ;
        RECT 50.900 28.300 51.500 29.600 ;
        RECT 52.400 28.300 53.200 29.600 ;
        RECT 50.900 27.700 53.200 28.300 ;
        RECT 41.200 25.600 42.000 26.400 ;
        RECT 43.000 26.200 43.600 27.600 ;
        RECT 41.400 24.800 42.200 25.600 ;
        RECT 42.800 22.200 43.600 26.200 ;
        RECT 47.600 24.800 48.400 26.400 ;
        RECT 49.400 24.200 50.000 27.600 ;
        RECT 49.200 22.200 50.000 24.200 ;
        RECT 52.400 22.200 53.200 27.700 ;
        RECT 54.200 27.400 54.800 30.400 ;
        RECT 55.600 28.800 56.400 30.400 ;
        RECT 63.600 29.000 64.400 34.600 ;
        RECT 66.200 34.400 70.400 35.200 ;
        RECT 74.800 35.000 75.600 39.800 ;
        RECT 78.000 35.000 78.800 39.800 ;
        RECT 66.200 34.000 66.800 34.400 ;
        RECT 65.200 33.200 66.800 34.000 ;
        RECT 69.800 33.800 75.600 34.400 ;
        RECT 67.800 33.200 69.200 33.800 ;
        RECT 67.800 33.000 74.000 33.200 ;
        RECT 68.600 32.600 74.000 33.000 ;
        RECT 73.200 32.400 74.000 32.600 ;
        RECT 75.000 33.000 75.600 33.800 ;
        RECT 76.200 33.600 78.800 34.400 ;
        RECT 81.200 33.600 82.000 39.800 ;
        RECT 82.800 37.000 83.600 39.800 ;
        RECT 84.400 37.000 85.200 39.800 ;
        RECT 86.000 37.000 86.800 39.800 ;
        RECT 84.400 34.400 88.600 35.200 ;
        RECT 89.200 34.400 90.000 39.800 ;
        RECT 92.400 35.200 93.200 39.800 ;
        RECT 92.400 34.600 95.000 35.200 ;
        RECT 89.200 33.600 91.800 34.400 ;
        RECT 82.800 33.000 83.600 33.200 ;
        RECT 75.000 32.400 83.600 33.000 ;
        RECT 86.000 33.000 86.800 33.200 ;
        RECT 94.400 33.000 95.000 34.600 ;
        RECT 86.000 32.400 95.000 33.000 ;
        RECT 94.400 30.600 95.000 32.400 ;
        RECT 95.600 32.000 96.400 39.800 ;
        RECT 101.400 32.600 102.200 39.800 ;
        RECT 95.600 31.200 96.600 32.000 ;
        RECT 100.400 31.800 102.200 32.600 ;
        RECT 103.600 31.800 104.400 39.800 ;
        RECT 105.200 32.400 106.000 39.800 ;
        RECT 108.400 32.400 109.200 39.800 ;
        RECT 105.200 31.800 109.200 32.400 ;
        RECT 65.000 30.000 88.400 30.600 ;
        RECT 94.400 30.000 95.200 30.600 ;
        RECT 65.000 29.800 66.000 30.000 ;
        RECT 65.200 29.600 66.000 29.800 ;
        RECT 70.000 29.600 70.800 30.000 ;
        RECT 76.400 29.600 77.200 30.000 ;
        RECT 87.600 29.400 88.400 30.000 ;
        RECT 63.600 28.200 72.400 29.000 ;
        RECT 73.000 28.600 75.000 29.400 ;
        RECT 78.800 28.600 82.000 29.400 ;
        RECT 54.200 26.800 56.400 27.400 ;
        RECT 55.600 22.200 56.400 26.800 ;
        RECT 63.600 22.200 64.400 28.200 ;
        RECT 66.000 26.800 69.000 27.600 ;
        RECT 68.200 26.200 69.000 26.800 ;
        RECT 74.200 26.200 75.000 28.600 ;
        RECT 76.400 26.800 77.200 28.400 ;
        RECT 81.600 27.800 82.400 28.000 ;
        RECT 78.000 27.200 82.400 27.800 ;
        RECT 78.000 27.000 78.800 27.200 ;
        RECT 84.400 26.400 85.200 29.200 ;
        RECT 90.200 28.600 94.000 29.400 ;
        RECT 90.200 27.400 91.000 28.600 ;
        RECT 94.600 28.000 95.200 30.000 ;
        RECT 78.000 26.200 78.800 26.400 ;
        RECT 68.200 25.400 70.800 26.200 ;
        RECT 74.200 25.600 78.800 26.200 ;
        RECT 79.600 25.600 81.200 26.400 ;
        RECT 84.200 25.600 85.200 26.400 ;
        RECT 89.200 26.800 91.000 27.400 ;
        RECT 94.000 27.400 95.200 28.000 ;
        RECT 89.200 26.200 90.000 26.800 ;
        RECT 70.000 22.200 70.800 25.400 ;
        RECT 87.600 25.400 90.000 26.200 ;
        RECT 71.600 22.200 72.400 25.000 ;
        RECT 73.200 22.200 74.000 25.000 ;
        RECT 74.800 22.200 75.600 25.000 ;
        RECT 78.000 22.200 78.800 25.000 ;
        RECT 81.200 22.200 82.000 25.000 ;
        RECT 82.800 22.200 83.600 25.000 ;
        RECT 84.400 22.200 85.200 25.000 ;
        RECT 86.000 22.200 86.800 25.000 ;
        RECT 87.600 22.200 88.400 25.400 ;
        RECT 94.000 22.200 94.800 27.400 ;
        RECT 95.800 26.800 96.600 31.200 ;
        RECT 100.600 28.400 101.200 31.800 ;
        RECT 102.000 29.600 102.800 31.200 ;
        RECT 103.800 30.400 104.400 31.800 ;
        RECT 111.600 31.200 112.400 39.800 ;
        RECT 114.800 31.200 115.600 39.800 ;
        RECT 118.000 31.200 118.800 39.800 ;
        RECT 121.200 31.200 122.000 39.800 ;
        RECT 124.400 31.600 125.200 33.200 ;
        RECT 107.600 30.400 108.400 30.800 ;
        RECT 111.600 30.400 113.400 31.200 ;
        RECT 114.800 30.400 117.000 31.200 ;
        RECT 118.000 30.400 120.200 31.200 ;
        RECT 121.200 30.400 123.600 31.200 ;
        RECT 103.600 29.800 106.000 30.400 ;
        RECT 107.600 29.800 109.200 30.400 ;
        RECT 103.600 29.600 104.400 29.800 ;
        RECT 100.400 27.600 101.200 28.400 ;
        RECT 102.000 28.300 102.800 28.400 ;
        RECT 105.400 28.300 106.000 29.800 ;
        RECT 108.400 29.600 109.200 29.800 ;
        RECT 102.000 27.700 106.000 28.300 ;
        RECT 102.000 27.600 102.800 27.700 ;
        RECT 95.600 26.300 96.600 26.800 ;
        RECT 98.800 26.300 99.600 26.400 ;
        RECT 100.600 26.300 101.200 27.600 ;
        RECT 103.600 26.300 104.400 26.400 ;
        RECT 95.600 25.700 99.600 26.300 ;
        RECT 100.500 25.700 104.400 26.300 ;
        RECT 105.400 26.200 106.000 27.700 ;
        RECT 106.800 27.600 107.600 29.200 ;
        RECT 112.600 29.000 113.400 30.400 ;
        RECT 116.200 29.000 117.000 30.400 ;
        RECT 119.400 29.000 120.200 30.400 ;
        RECT 112.600 28.200 115.200 29.000 ;
        RECT 116.200 28.200 118.600 29.000 ;
        RECT 119.400 28.200 122.000 29.000 ;
        RECT 112.600 27.600 113.400 28.200 ;
        RECT 116.200 27.600 117.000 28.200 ;
        RECT 119.400 27.600 120.200 28.200 ;
        RECT 122.800 27.600 123.600 30.400 ;
        RECT 95.600 22.200 96.400 25.700 ;
        RECT 98.800 24.800 99.600 25.700 ;
        RECT 100.600 24.200 101.200 25.700 ;
        RECT 103.600 25.600 104.400 25.700 ;
        RECT 103.800 24.800 104.600 25.600 ;
        RECT 100.400 22.200 101.200 24.200 ;
        RECT 105.200 22.200 106.000 26.200 ;
        RECT 111.600 26.800 113.400 27.600 ;
        RECT 114.800 26.800 117.000 27.600 ;
        RECT 118.000 26.800 120.200 27.600 ;
        RECT 121.200 26.800 123.600 27.600 ;
        RECT 111.600 22.200 112.400 26.800 ;
        RECT 114.800 22.200 115.600 26.800 ;
        RECT 118.000 22.200 118.800 26.800 ;
        RECT 121.200 22.200 122.000 26.800 ;
        RECT 126.000 26.200 126.800 39.800 ;
        RECT 130.800 31.200 131.600 39.800 ;
        RECT 134.000 31.200 134.800 39.800 ;
        RECT 137.200 31.200 138.000 39.800 ;
        RECT 140.400 31.200 141.200 39.800 ;
        RECT 143.600 32.400 144.400 39.800 ;
        RECT 143.600 31.800 145.800 32.400 ;
        RECT 146.800 31.800 147.600 39.800 ;
        RECT 150.000 36.400 150.800 39.800 ;
        RECT 149.800 35.800 150.800 36.400 ;
        RECT 149.800 35.200 150.400 35.800 ;
        RECT 153.200 35.200 154.000 39.800 ;
        RECT 156.400 37.000 157.200 39.800 ;
        RECT 158.000 37.000 158.800 39.800 ;
        RECT 145.200 31.200 145.800 31.800 ;
        RECT 130.800 30.400 132.600 31.200 ;
        RECT 134.000 30.400 136.200 31.200 ;
        RECT 137.200 30.400 139.400 31.200 ;
        RECT 140.400 30.400 142.800 31.200 ;
        RECT 145.200 30.400 146.400 31.200 ;
        RECT 131.800 29.000 132.600 30.400 ;
        RECT 135.400 29.000 136.200 30.400 ;
        RECT 138.600 29.000 139.400 30.400 ;
        RECT 131.800 28.200 134.400 29.000 ;
        RECT 135.400 28.200 137.800 29.000 ;
        RECT 138.600 28.200 141.200 29.000 ;
        RECT 131.800 27.600 132.600 28.200 ;
        RECT 135.400 27.600 136.200 28.200 ;
        RECT 138.600 27.600 139.400 28.200 ;
        RECT 142.000 27.600 142.800 30.400 ;
        RECT 143.600 28.800 144.400 30.400 ;
        RECT 125.000 25.600 126.800 26.200 ;
        RECT 130.800 26.800 132.600 27.600 ;
        RECT 134.000 26.800 136.200 27.600 ;
        RECT 137.200 26.800 139.400 27.600 ;
        RECT 140.400 26.800 142.800 27.600 ;
        RECT 145.200 27.400 145.800 30.400 ;
        RECT 147.000 29.600 147.600 31.800 ;
        RECT 143.600 26.800 145.800 27.400 ;
        RECT 125.000 24.400 125.800 25.600 ;
        RECT 124.400 23.600 125.800 24.400 ;
        RECT 125.000 22.200 125.800 23.600 ;
        RECT 130.800 22.200 131.600 26.800 ;
        RECT 134.000 22.200 134.800 26.800 ;
        RECT 137.200 22.200 138.000 26.800 ;
        RECT 140.400 22.200 141.200 26.800 ;
        RECT 143.600 22.200 144.400 26.800 ;
        RECT 146.800 22.200 147.600 29.600 ;
        RECT 148.400 34.600 150.400 35.200 ;
        RECT 148.400 29.000 149.200 34.600 ;
        RECT 151.000 34.400 155.200 35.200 ;
        RECT 159.600 35.000 160.400 39.800 ;
        RECT 162.800 35.000 163.600 39.800 ;
        RECT 151.000 34.000 151.600 34.400 ;
        RECT 150.000 33.200 151.600 34.000 ;
        RECT 154.600 33.800 160.400 34.400 ;
        RECT 152.600 33.200 154.000 33.800 ;
        RECT 152.600 33.000 158.800 33.200 ;
        RECT 153.400 32.600 158.800 33.000 ;
        RECT 158.000 32.400 158.800 32.600 ;
        RECT 159.800 33.000 160.400 33.800 ;
        RECT 161.000 33.600 163.600 34.400 ;
        RECT 166.000 33.600 166.800 39.800 ;
        RECT 167.600 37.000 168.400 39.800 ;
        RECT 169.200 37.000 170.000 39.800 ;
        RECT 170.800 37.000 171.600 39.800 ;
        RECT 169.200 34.400 173.400 35.200 ;
        RECT 174.000 34.400 174.800 39.800 ;
        RECT 177.200 35.200 178.000 39.800 ;
        RECT 177.200 34.600 179.800 35.200 ;
        RECT 174.000 33.600 176.600 34.400 ;
        RECT 167.600 33.000 168.400 33.200 ;
        RECT 159.800 32.400 168.400 33.000 ;
        RECT 170.800 33.000 171.600 33.200 ;
        RECT 179.200 33.000 179.800 34.600 ;
        RECT 170.800 32.400 179.800 33.000 ;
        RECT 179.200 30.600 179.800 32.400 ;
        RECT 180.400 32.000 181.200 39.800 ;
        RECT 193.200 32.400 194.000 39.800 ;
        RECT 180.400 31.200 181.400 32.000 ;
        RECT 191.800 31.800 194.000 32.400 ;
        RECT 196.400 32.300 197.200 39.800 ;
        RECT 198.800 33.600 199.600 34.400 ;
        RECT 198.800 32.400 199.400 33.600 ;
        RECT 200.200 32.400 201.000 39.800 ;
        RECT 198.000 32.300 199.400 32.400 ;
        RECT 196.400 31.800 199.400 32.300 ;
        RECT 200.000 31.800 201.000 32.400 ;
        RECT 191.800 31.200 192.400 31.800 ;
        RECT 149.800 30.000 173.200 30.600 ;
        RECT 179.200 30.000 180.000 30.600 ;
        RECT 149.800 29.800 150.600 30.000 ;
        RECT 151.600 29.600 152.400 30.000 ;
        RECT 154.800 29.600 155.600 30.000 ;
        RECT 172.400 29.400 173.200 30.000 ;
        RECT 148.400 28.200 157.200 29.000 ;
        RECT 157.800 28.600 159.800 29.400 ;
        RECT 163.600 28.600 166.800 29.400 ;
        RECT 148.400 22.200 149.200 28.200 ;
        RECT 150.800 26.800 153.800 27.600 ;
        RECT 153.000 26.200 153.800 26.800 ;
        RECT 159.000 26.200 159.800 28.600 ;
        RECT 161.200 26.800 162.000 28.400 ;
        RECT 166.400 27.800 167.200 28.000 ;
        RECT 162.800 27.200 167.200 27.800 ;
        RECT 162.800 27.000 163.600 27.200 ;
        RECT 169.200 26.400 170.000 29.200 ;
        RECT 175.000 28.600 178.800 29.400 ;
        RECT 175.000 27.400 175.800 28.600 ;
        RECT 179.400 28.000 180.000 30.000 ;
        RECT 162.800 26.200 163.600 26.400 ;
        RECT 153.000 25.400 155.600 26.200 ;
        RECT 159.000 25.600 163.600 26.200 ;
        RECT 164.400 25.600 166.000 26.400 ;
        RECT 169.000 25.600 170.000 26.400 ;
        RECT 174.000 26.800 175.800 27.400 ;
        RECT 178.800 27.400 180.000 28.000 ;
        RECT 174.000 26.200 174.800 26.800 ;
        RECT 154.800 22.200 155.600 25.400 ;
        RECT 172.400 25.400 174.800 26.200 ;
        RECT 156.400 22.200 157.200 25.000 ;
        RECT 158.000 22.200 158.800 25.000 ;
        RECT 159.600 22.200 160.400 25.000 ;
        RECT 162.800 22.200 163.600 25.000 ;
        RECT 166.000 22.200 166.800 25.000 ;
        RECT 167.600 22.200 168.400 25.000 ;
        RECT 169.200 22.200 170.000 25.000 ;
        RECT 170.800 22.200 171.600 25.000 ;
        RECT 172.400 22.200 173.200 25.400 ;
        RECT 178.800 22.200 179.600 27.400 ;
        RECT 180.600 26.800 181.400 31.200 ;
        RECT 191.200 30.400 192.400 31.200 ;
        RECT 196.400 31.700 198.800 31.800 ;
        RECT 191.800 27.400 192.400 30.400 ;
        RECT 193.200 28.800 194.000 30.400 ;
        RECT 191.800 26.800 194.000 27.400 ;
        RECT 180.400 26.000 181.400 26.800 ;
        RECT 180.400 22.200 181.200 26.000 ;
        RECT 193.200 22.200 194.000 26.800 ;
        RECT 194.800 24.800 195.600 26.400 ;
        RECT 196.400 22.200 197.200 31.700 ;
        RECT 198.000 31.600 198.800 31.700 ;
        RECT 200.000 28.400 200.600 31.800 ;
        RECT 201.200 30.300 202.000 30.400 ;
        RECT 202.800 30.300 203.600 30.400 ;
        RECT 201.200 29.700 203.600 30.300 ;
        RECT 201.200 28.800 202.000 29.700 ;
        RECT 202.800 29.600 203.600 29.700 ;
        RECT 198.000 27.600 200.600 28.400 ;
        RECT 202.800 28.300 203.600 28.400 ;
        RECT 204.400 28.300 205.200 39.800 ;
        RECT 209.200 36.400 210.000 39.800 ;
        RECT 209.000 35.800 210.000 36.400 ;
        RECT 209.000 35.200 209.600 35.800 ;
        RECT 212.400 35.200 213.200 39.800 ;
        RECT 215.600 37.000 216.400 39.800 ;
        RECT 217.200 37.000 218.000 39.800 ;
        RECT 202.800 28.200 205.200 28.300 ;
        RECT 202.000 27.700 205.200 28.200 ;
        RECT 202.000 27.600 203.600 27.700 ;
        RECT 198.200 26.200 198.800 27.600 ;
        RECT 202.000 27.200 202.800 27.600 ;
        RECT 199.800 26.200 203.400 26.600 ;
        RECT 198.000 22.200 198.800 26.200 ;
        RECT 199.600 26.000 203.600 26.200 ;
        RECT 199.600 22.200 200.400 26.000 ;
        RECT 202.800 22.200 203.600 26.000 ;
        RECT 204.400 22.200 205.200 27.700 ;
        RECT 207.600 34.600 209.600 35.200 ;
        RECT 207.600 29.000 208.400 34.600 ;
        RECT 210.200 34.400 214.400 35.200 ;
        RECT 218.800 35.000 219.600 39.800 ;
        RECT 222.000 35.000 222.800 39.800 ;
        RECT 210.200 34.000 210.800 34.400 ;
        RECT 209.200 33.200 210.800 34.000 ;
        RECT 213.800 33.800 219.600 34.400 ;
        RECT 211.800 33.200 213.200 33.800 ;
        RECT 211.800 33.000 218.000 33.200 ;
        RECT 212.600 32.600 218.000 33.000 ;
        RECT 217.200 32.400 218.000 32.600 ;
        RECT 219.000 33.000 219.600 33.800 ;
        RECT 220.200 33.600 222.800 34.400 ;
        RECT 225.200 33.600 226.000 39.800 ;
        RECT 226.800 37.000 227.600 39.800 ;
        RECT 228.400 37.000 229.200 39.800 ;
        RECT 230.000 37.000 230.800 39.800 ;
        RECT 228.400 34.400 232.600 35.200 ;
        RECT 233.200 34.400 234.000 39.800 ;
        RECT 236.400 35.200 237.200 39.800 ;
        RECT 236.400 34.600 239.000 35.200 ;
        RECT 233.200 33.600 235.800 34.400 ;
        RECT 226.800 33.000 227.600 33.200 ;
        RECT 219.000 32.400 227.600 33.000 ;
        RECT 230.000 33.000 230.800 33.200 ;
        RECT 238.400 33.000 239.000 34.600 ;
        RECT 230.000 32.400 239.000 33.000 ;
        RECT 210.800 31.800 211.600 32.400 ;
        RECT 214.000 31.800 215.000 32.000 ;
        RECT 210.800 31.200 237.800 31.800 ;
        RECT 237.000 31.000 237.800 31.200 ;
        RECT 238.400 30.600 239.000 32.400 ;
        RECT 239.600 32.000 240.400 39.800 ;
        RECT 239.600 31.200 240.600 32.000 ;
        RECT 238.400 30.000 239.200 30.600 ;
        RECT 207.600 28.200 216.400 29.000 ;
        RECT 217.000 28.600 219.000 29.400 ;
        RECT 222.800 28.600 226.000 29.400 ;
        RECT 206.000 24.800 206.800 26.400 ;
        RECT 207.600 22.200 208.400 28.200 ;
        RECT 210.000 26.800 213.000 27.600 ;
        RECT 212.200 26.200 213.000 26.800 ;
        RECT 218.200 26.200 219.000 28.600 ;
        RECT 220.400 26.800 221.200 28.400 ;
        RECT 225.600 27.800 226.400 28.000 ;
        RECT 222.000 27.200 226.400 27.800 ;
        RECT 222.000 27.000 222.800 27.200 ;
        RECT 228.400 26.400 229.200 29.200 ;
        RECT 234.200 28.600 238.000 29.400 ;
        RECT 234.200 27.400 235.000 28.600 ;
        RECT 238.600 28.000 239.200 30.000 ;
        RECT 222.000 26.200 222.800 26.400 ;
        RECT 212.200 25.400 214.800 26.200 ;
        RECT 218.200 25.600 222.800 26.200 ;
        RECT 223.600 25.600 225.200 26.400 ;
        RECT 228.200 25.600 229.200 26.400 ;
        RECT 233.200 26.800 235.000 27.400 ;
        RECT 238.000 27.400 239.200 28.000 ;
        RECT 233.200 26.200 234.000 26.800 ;
        RECT 214.000 22.200 214.800 25.400 ;
        RECT 231.600 25.400 234.000 26.200 ;
        RECT 215.600 22.200 216.400 25.000 ;
        RECT 217.200 22.200 218.000 25.000 ;
        RECT 218.800 22.200 219.600 25.000 ;
        RECT 222.000 22.200 222.800 25.000 ;
        RECT 225.200 22.200 226.000 25.000 ;
        RECT 226.800 22.200 227.600 25.000 ;
        RECT 228.400 22.200 229.200 25.000 ;
        RECT 230.000 22.200 230.800 25.000 ;
        RECT 231.600 22.200 232.400 25.400 ;
        RECT 238.000 22.200 238.800 27.400 ;
        RECT 239.800 26.800 240.600 31.200 ;
        RECT 239.600 26.000 240.600 26.800 ;
        RECT 239.600 22.200 240.400 26.000 ;
        RECT 242.800 22.200 243.600 39.800 ;
        RECT 246.000 32.400 246.800 39.800 ;
        RECT 246.000 31.800 248.200 32.400 ;
        RECT 247.600 31.200 248.200 31.800 ;
        RECT 247.600 30.400 248.800 31.200 ;
        RECT 246.000 28.800 246.800 30.400 ;
        RECT 247.600 27.400 248.200 30.400 ;
        RECT 246.000 26.800 248.200 27.400 ;
        RECT 246.000 22.200 246.800 26.800 ;
        RECT 4.400 15.200 5.200 19.800 ;
        RECT 7.600 16.000 8.400 19.800 ;
        RECT 3.000 14.600 5.200 15.200 ;
        RECT 7.400 15.200 8.400 16.000 ;
        RECT 3.000 11.600 3.600 14.600 ;
        RECT 4.400 12.300 5.200 13.200 ;
        RECT 7.400 12.300 8.200 15.200 ;
        RECT 9.200 14.600 10.000 19.800 ;
        RECT 15.600 16.600 16.400 19.800 ;
        RECT 17.200 17.000 18.000 19.800 ;
        RECT 18.800 17.000 19.600 19.800 ;
        RECT 20.400 17.000 21.200 19.800 ;
        RECT 22.000 17.000 22.800 19.800 ;
        RECT 25.200 17.000 26.000 19.800 ;
        RECT 28.400 17.000 29.200 19.800 ;
        RECT 30.000 17.000 30.800 19.800 ;
        RECT 31.600 17.000 32.400 19.800 ;
        RECT 14.000 15.800 16.400 16.600 ;
        RECT 33.200 16.600 34.000 19.800 ;
        RECT 14.000 15.200 14.800 15.800 ;
        RECT 4.400 11.700 8.200 12.300 ;
        RECT 4.400 11.600 5.200 11.700 ;
        RECT 2.400 10.800 3.600 11.600 ;
        RECT 3.000 10.200 3.600 10.800 ;
        RECT 7.400 10.800 8.200 11.700 ;
        RECT 8.800 14.000 10.000 14.600 ;
        RECT 13.000 14.600 14.800 15.200 ;
        RECT 18.800 15.600 19.800 16.400 ;
        RECT 22.800 15.600 24.400 16.400 ;
        RECT 25.200 15.800 29.800 16.400 ;
        RECT 33.200 15.800 35.800 16.600 ;
        RECT 25.200 15.600 26.000 15.800 ;
        RECT 8.800 12.000 9.400 14.000 ;
        RECT 13.000 13.400 13.800 14.600 ;
        RECT 10.000 12.600 13.800 13.400 ;
        RECT 18.800 12.800 19.600 15.600 ;
        RECT 25.200 14.800 26.000 15.000 ;
        RECT 21.600 14.200 26.000 14.800 ;
        RECT 21.600 14.000 22.400 14.200 ;
        RECT 26.800 13.600 27.600 15.200 ;
        RECT 29.000 13.400 29.800 15.800 ;
        RECT 35.000 15.200 35.800 15.800 ;
        RECT 35.000 14.400 38.000 15.200 ;
        RECT 39.600 13.800 40.400 19.800 ;
        RECT 42.800 17.800 43.600 19.800 ;
        RECT 41.200 15.600 42.000 17.200 ;
        RECT 43.000 16.300 43.600 17.800 ;
        RECT 46.200 16.400 47.000 17.200 ;
        RECT 46.000 16.300 46.800 16.400 ;
        RECT 42.900 15.700 46.800 16.300 ;
        RECT 43.000 14.400 43.600 15.700 ;
        RECT 46.000 15.600 46.800 15.700 ;
        RECT 47.600 15.600 48.400 19.800 ;
        RECT 22.000 12.600 25.200 13.400 ;
        RECT 29.000 12.600 31.000 13.400 ;
        RECT 31.600 13.000 40.400 13.800 ;
        RECT 42.800 13.600 43.600 14.400 ;
        RECT 15.600 12.000 16.400 12.600 ;
        RECT 33.200 12.000 34.000 12.400 ;
        RECT 36.400 12.000 37.200 12.400 ;
        RECT 38.200 12.000 39.000 12.200 ;
        RECT 8.800 11.400 9.600 12.000 ;
        RECT 15.600 11.400 39.000 12.000 ;
        RECT 3.000 9.600 5.200 10.200 ;
        RECT 7.400 10.000 8.400 10.800 ;
        RECT 4.400 2.200 5.200 9.600 ;
        RECT 7.600 2.200 8.400 10.000 ;
        RECT 9.000 9.600 9.600 11.400 ;
        RECT 9.000 9.000 18.000 9.600 ;
        RECT 9.000 7.400 9.600 9.000 ;
        RECT 17.200 8.800 18.000 9.000 ;
        RECT 20.400 9.000 29.000 9.600 ;
        RECT 20.400 8.800 21.200 9.000 ;
        RECT 12.200 7.600 14.800 8.400 ;
        RECT 9.000 6.800 11.600 7.400 ;
        RECT 10.800 2.200 11.600 6.800 ;
        RECT 14.000 2.200 14.800 7.600 ;
        RECT 15.400 6.800 19.600 7.600 ;
        RECT 17.200 2.200 18.000 5.000 ;
        RECT 18.800 2.200 19.600 5.000 ;
        RECT 20.400 2.200 21.200 5.000 ;
        RECT 22.000 2.200 22.800 8.400 ;
        RECT 25.200 7.600 27.800 8.400 ;
        RECT 28.400 8.200 29.000 9.000 ;
        RECT 30.000 9.400 30.800 9.600 ;
        RECT 30.000 9.000 35.400 9.400 ;
        RECT 30.000 8.800 36.200 9.000 ;
        RECT 34.800 8.200 36.200 8.800 ;
        RECT 28.400 7.600 34.200 8.200 ;
        RECT 37.200 8.000 38.800 8.800 ;
        RECT 37.200 7.600 37.800 8.000 ;
        RECT 25.200 2.200 26.000 7.000 ;
        RECT 28.400 2.200 29.200 7.000 ;
        RECT 33.600 6.800 37.800 7.600 ;
        RECT 39.600 7.400 40.400 13.000 ;
        RECT 43.000 10.200 43.600 13.600 ;
        RECT 44.400 10.800 45.200 12.400 ;
        RECT 46.000 12.200 46.800 12.400 ;
        RECT 47.800 12.200 48.400 15.600 ;
        RECT 49.200 14.300 50.000 14.400 ;
        RECT 52.400 14.300 53.200 14.400 ;
        RECT 49.200 13.700 53.200 14.300 ;
        RECT 49.200 12.800 50.000 13.700 ;
        RECT 52.400 13.600 53.200 13.700 ;
        RECT 58.800 13.800 59.600 19.800 ;
        RECT 65.200 16.600 66.000 19.800 ;
        RECT 66.800 17.000 67.600 19.800 ;
        RECT 68.400 17.000 69.200 19.800 ;
        RECT 70.000 17.000 70.800 19.800 ;
        RECT 73.200 17.000 74.000 19.800 ;
        RECT 76.400 17.000 77.200 19.800 ;
        RECT 78.000 17.000 78.800 19.800 ;
        RECT 79.600 17.000 80.400 19.800 ;
        RECT 81.200 17.000 82.000 19.800 ;
        RECT 63.400 15.800 66.000 16.600 ;
        RECT 82.800 16.600 83.600 19.800 ;
        RECT 69.400 15.800 74.000 16.400 ;
        RECT 63.400 15.200 64.200 15.800 ;
        RECT 61.200 14.400 64.200 15.200 ;
        RECT 58.800 13.000 67.600 13.800 ;
        RECT 69.400 13.400 70.200 15.800 ;
        RECT 73.200 15.600 74.000 15.800 ;
        RECT 74.800 15.600 76.400 16.400 ;
        RECT 79.400 15.600 80.400 16.400 ;
        RECT 82.800 15.800 85.200 16.600 ;
        RECT 73.200 14.800 74.000 15.000 ;
        RECT 73.200 14.200 77.600 14.800 ;
        RECT 76.800 14.000 77.600 14.200 ;
        RECT 50.800 12.200 51.600 12.400 ;
        RECT 46.000 11.600 48.400 12.200 ;
        RECT 50.000 11.600 51.600 12.200 ;
        RECT 46.200 10.200 46.800 11.600 ;
        RECT 50.000 11.200 50.800 11.600 ;
        RECT 42.800 9.400 44.600 10.200 ;
        RECT 38.400 6.800 40.400 7.400 ;
        RECT 30.000 2.200 30.800 5.000 ;
        RECT 31.600 2.200 32.400 5.000 ;
        RECT 34.800 2.200 35.600 6.800 ;
        RECT 38.400 6.200 39.000 6.800 ;
        RECT 38.000 5.600 39.000 6.200 ;
        RECT 38.000 2.200 38.800 5.600 ;
        RECT 43.800 2.200 44.600 9.400 ;
        RECT 46.000 2.200 46.800 10.200 ;
        RECT 47.600 9.600 51.600 10.200 ;
        RECT 47.600 2.200 48.400 9.600 ;
        RECT 50.800 2.200 51.600 9.600 ;
        RECT 58.800 7.400 59.600 13.000 ;
        RECT 68.200 12.600 70.200 13.400 ;
        RECT 74.000 12.600 77.200 13.400 ;
        RECT 79.600 12.800 80.400 15.600 ;
        RECT 84.400 15.200 85.200 15.800 ;
        RECT 84.400 14.600 86.200 15.200 ;
        RECT 85.400 13.400 86.200 14.600 ;
        RECT 89.200 14.600 90.000 19.800 ;
        RECT 90.800 16.000 91.600 19.800 ;
        RECT 90.800 15.200 91.800 16.000 ;
        RECT 89.200 14.000 90.400 14.600 ;
        RECT 85.400 12.600 89.200 13.400 ;
        RECT 60.200 12.000 61.000 12.200 ;
        RECT 63.600 12.000 64.400 12.400 ;
        RECT 65.200 12.000 66.000 12.400 ;
        RECT 82.800 12.000 83.600 12.600 ;
        RECT 89.800 12.000 90.400 14.000 ;
        RECT 60.200 11.400 83.600 12.000 ;
        RECT 89.600 11.400 90.400 12.000 ;
        RECT 89.600 9.600 90.200 11.400 ;
        RECT 91.000 10.800 91.800 15.200 ;
        RECT 94.000 15.200 94.800 19.800 ;
        RECT 100.400 15.200 101.200 19.800 ;
        RECT 103.600 15.200 104.400 19.800 ;
        RECT 110.000 15.200 110.800 19.800 ;
        RECT 111.600 15.600 112.400 17.200 ;
        RECT 94.000 14.600 96.200 15.200 ;
        RECT 94.000 11.600 94.800 13.200 ;
        RECT 95.600 11.600 96.200 14.600 ;
        RECT 100.400 14.400 104.400 15.200 ;
        RECT 108.600 14.600 110.800 15.200 ;
        RECT 100.400 11.600 101.200 14.400 ;
        RECT 108.600 11.600 109.200 14.600 ;
        RECT 113.200 14.300 114.000 19.800 ;
        RECT 114.800 16.000 115.600 19.800 ;
        RECT 118.000 16.000 118.800 19.800 ;
        RECT 114.800 15.800 118.800 16.000 ;
        RECT 119.600 16.300 120.400 19.800 ;
        RECT 121.200 16.300 122.000 16.400 ;
        RECT 115.000 15.400 118.600 15.800 ;
        RECT 119.600 15.700 122.000 16.300 ;
        RECT 122.800 16.000 123.600 19.800 ;
        RECT 115.600 14.400 116.400 14.800 ;
        RECT 119.600 14.400 120.200 15.700 ;
        RECT 121.200 15.600 122.000 15.700 ;
        RECT 122.600 15.200 123.600 16.000 ;
        RECT 114.800 14.300 116.400 14.400 ;
        RECT 113.200 13.800 116.400 14.300 ;
        RECT 113.200 13.700 115.600 13.800 ;
        RECT 110.000 12.300 110.800 13.200 ;
        RECT 111.600 12.300 112.400 12.400 ;
        RECT 110.000 11.700 112.400 12.300 ;
        RECT 110.000 11.600 110.800 11.700 ;
        RECT 111.600 11.600 112.400 11.700 ;
        RECT 68.400 9.400 69.200 9.600 ;
        RECT 63.800 9.000 69.200 9.400 ;
        RECT 63.000 8.800 69.200 9.000 ;
        RECT 70.200 9.000 78.800 9.600 ;
        RECT 60.400 8.000 62.000 8.800 ;
        RECT 63.000 8.200 64.400 8.800 ;
        RECT 70.200 8.200 70.800 9.000 ;
        RECT 78.000 8.800 78.800 9.000 ;
        RECT 81.200 9.000 90.200 9.600 ;
        RECT 81.200 8.800 82.000 9.000 ;
        RECT 61.400 7.600 62.000 8.000 ;
        RECT 65.000 7.600 70.800 8.200 ;
        RECT 71.400 7.600 74.000 8.400 ;
        RECT 58.800 6.800 60.800 7.400 ;
        RECT 61.400 6.800 65.600 7.600 ;
        RECT 60.200 6.200 60.800 6.800 ;
        RECT 60.200 5.600 61.200 6.200 ;
        RECT 60.400 2.200 61.200 5.600 ;
        RECT 63.600 2.200 64.400 6.800 ;
        RECT 66.800 2.200 67.600 5.000 ;
        RECT 68.400 2.200 69.200 5.000 ;
        RECT 70.000 2.200 70.800 7.000 ;
        RECT 73.200 2.200 74.000 7.000 ;
        RECT 76.400 2.200 77.200 8.400 ;
        RECT 84.400 7.600 87.000 8.400 ;
        RECT 79.600 6.800 83.800 7.600 ;
        RECT 78.000 2.200 78.800 5.000 ;
        RECT 79.600 2.200 80.400 5.000 ;
        RECT 81.200 2.200 82.000 5.000 ;
        RECT 84.400 2.200 85.200 7.600 ;
        RECT 89.600 7.400 90.200 9.000 ;
        RECT 87.600 6.800 90.200 7.400 ;
        RECT 90.800 10.000 91.800 10.800 ;
        RECT 95.600 10.800 96.800 11.600 ;
        RECT 100.400 10.800 104.400 11.600 ;
        RECT 108.000 10.800 109.200 11.600 ;
        RECT 95.600 10.200 96.200 10.800 ;
        RECT 87.600 2.200 88.400 6.800 ;
        RECT 90.800 2.200 91.600 10.000 ;
        RECT 94.000 9.600 96.200 10.200 ;
        RECT 94.000 2.200 94.800 9.600 ;
        RECT 100.400 2.200 101.200 10.800 ;
        RECT 103.600 2.200 104.400 10.800 ;
        RECT 108.600 10.200 109.200 10.800 ;
        RECT 108.600 9.600 110.800 10.200 ;
        RECT 110.000 2.200 110.800 9.600 ;
        RECT 113.200 2.200 114.000 13.700 ;
        RECT 114.800 13.600 115.600 13.700 ;
        RECT 117.800 13.600 120.400 14.400 ;
        RECT 116.400 11.600 117.200 13.200 ;
        RECT 117.800 10.200 118.400 13.600 ;
        RECT 122.600 10.800 123.400 15.200 ;
        RECT 124.400 14.600 125.200 19.800 ;
        RECT 130.800 16.600 131.600 19.800 ;
        RECT 132.400 17.000 133.200 19.800 ;
        RECT 134.000 17.000 134.800 19.800 ;
        RECT 135.600 17.000 136.400 19.800 ;
        RECT 137.200 17.000 138.000 19.800 ;
        RECT 140.400 17.000 141.200 19.800 ;
        RECT 143.600 17.000 144.400 19.800 ;
        RECT 145.200 17.000 146.000 19.800 ;
        RECT 146.800 17.000 147.600 19.800 ;
        RECT 129.200 15.800 131.600 16.600 ;
        RECT 148.400 16.600 149.200 19.800 ;
        RECT 129.200 15.200 130.000 15.800 ;
        RECT 124.000 14.000 125.200 14.600 ;
        RECT 128.200 14.600 130.000 15.200 ;
        RECT 134.000 15.600 135.000 16.400 ;
        RECT 138.000 15.600 139.600 16.400 ;
        RECT 140.400 15.800 145.000 16.400 ;
        RECT 148.400 15.800 151.000 16.600 ;
        RECT 140.400 15.600 141.200 15.800 ;
        RECT 124.000 12.000 124.600 14.000 ;
        RECT 128.200 13.400 129.000 14.600 ;
        RECT 125.200 12.600 129.000 13.400 ;
        RECT 134.000 12.800 134.800 15.600 ;
        RECT 140.400 14.800 141.200 15.000 ;
        RECT 136.800 14.200 141.200 14.800 ;
        RECT 136.800 14.000 137.600 14.200 ;
        RECT 142.000 13.600 142.800 15.200 ;
        RECT 144.200 13.400 145.000 15.800 ;
        RECT 150.200 15.200 151.000 15.800 ;
        RECT 150.200 14.400 153.200 15.200 ;
        RECT 154.800 13.800 155.600 19.800 ;
        RECT 137.200 12.600 140.400 13.400 ;
        RECT 144.200 12.600 146.200 13.400 ;
        RECT 146.800 13.000 155.600 13.800 ;
        RECT 130.800 12.000 131.600 12.600 ;
        RECT 148.400 12.000 149.200 12.400 ;
        RECT 151.600 12.000 152.400 12.400 ;
        RECT 153.400 12.000 154.200 12.200 ;
        RECT 124.000 11.400 124.800 12.000 ;
        RECT 130.800 11.400 154.200 12.000 ;
        RECT 119.600 10.200 120.400 10.400 ;
        RECT 117.400 9.600 118.400 10.200 ;
        RECT 119.000 9.600 120.400 10.200 ;
        RECT 122.600 10.000 123.600 10.800 ;
        RECT 117.400 2.200 118.200 9.600 ;
        RECT 119.000 8.400 119.600 9.600 ;
        RECT 118.800 7.600 119.600 8.400 ;
        RECT 122.800 2.200 123.600 10.000 ;
        RECT 124.200 9.600 124.800 11.400 ;
        RECT 124.200 9.000 133.200 9.600 ;
        RECT 124.200 7.400 124.800 9.000 ;
        RECT 132.400 8.800 133.200 9.000 ;
        RECT 135.600 9.000 144.200 9.600 ;
        RECT 135.600 8.800 136.400 9.000 ;
        RECT 127.400 7.600 130.000 8.400 ;
        RECT 124.200 6.800 126.800 7.400 ;
        RECT 126.000 2.200 126.800 6.800 ;
        RECT 129.200 2.200 130.000 7.600 ;
        RECT 130.600 6.800 134.800 7.600 ;
        RECT 132.400 2.200 133.200 5.000 ;
        RECT 134.000 2.200 134.800 5.000 ;
        RECT 135.600 2.200 136.400 5.000 ;
        RECT 137.200 2.200 138.000 8.400 ;
        RECT 140.400 7.600 143.000 8.400 ;
        RECT 143.600 8.200 144.200 9.000 ;
        RECT 145.200 9.400 146.000 9.600 ;
        RECT 145.200 9.000 150.600 9.400 ;
        RECT 145.200 8.800 151.400 9.000 ;
        RECT 150.000 8.200 151.400 8.800 ;
        RECT 143.600 7.600 149.400 8.200 ;
        RECT 152.400 8.000 154.000 8.800 ;
        RECT 152.400 7.600 153.000 8.000 ;
        RECT 140.400 2.200 141.200 7.000 ;
        RECT 143.600 2.200 144.400 7.000 ;
        RECT 148.800 6.800 153.000 7.600 ;
        RECT 154.800 7.400 155.600 13.000 ;
        RECT 153.600 6.800 155.600 7.400 ;
        RECT 156.400 13.800 157.200 19.800 ;
        RECT 162.800 16.600 163.600 19.800 ;
        RECT 164.400 17.000 165.200 19.800 ;
        RECT 166.000 17.000 166.800 19.800 ;
        RECT 167.600 17.000 168.400 19.800 ;
        RECT 170.800 17.000 171.600 19.800 ;
        RECT 174.000 17.000 174.800 19.800 ;
        RECT 175.600 17.000 176.400 19.800 ;
        RECT 177.200 17.000 178.000 19.800 ;
        RECT 178.800 17.000 179.600 19.800 ;
        RECT 161.000 15.800 163.600 16.600 ;
        RECT 180.400 16.600 181.200 19.800 ;
        RECT 167.000 15.800 171.600 16.400 ;
        RECT 161.000 15.200 161.800 15.800 ;
        RECT 158.800 14.400 161.800 15.200 ;
        RECT 156.400 13.000 165.200 13.800 ;
        RECT 167.000 13.400 167.800 15.800 ;
        RECT 170.800 15.600 171.600 15.800 ;
        RECT 172.400 15.600 174.000 16.400 ;
        RECT 177.000 15.600 178.000 16.400 ;
        RECT 180.400 15.800 182.800 16.600 ;
        RECT 169.200 13.600 170.000 15.200 ;
        RECT 170.800 14.800 171.600 15.000 ;
        RECT 170.800 14.200 175.200 14.800 ;
        RECT 174.400 14.000 175.200 14.200 ;
        RECT 156.400 7.400 157.200 13.000 ;
        RECT 165.800 12.600 167.800 13.400 ;
        RECT 171.600 12.600 174.800 13.400 ;
        RECT 177.200 12.800 178.000 15.600 ;
        RECT 182.000 15.200 182.800 15.800 ;
        RECT 182.000 14.600 183.800 15.200 ;
        RECT 183.000 13.400 183.800 14.600 ;
        RECT 186.800 14.600 187.600 19.800 ;
        RECT 188.400 16.000 189.200 19.800 ;
        RECT 190.000 16.300 190.800 16.400 ;
        RECT 198.000 16.300 198.800 17.200 ;
        RECT 188.400 15.200 189.400 16.000 ;
        RECT 190.000 15.700 198.800 16.300 ;
        RECT 190.000 15.600 190.800 15.700 ;
        RECT 198.000 15.600 198.800 15.700 ;
        RECT 186.800 14.000 188.000 14.600 ;
        RECT 183.000 12.600 186.800 13.400 ;
        RECT 157.800 12.000 158.600 12.200 ;
        RECT 159.600 12.000 160.400 12.400 ;
        RECT 162.800 12.000 163.600 12.400 ;
        RECT 180.400 12.000 181.200 12.600 ;
        RECT 187.400 12.000 188.000 14.000 ;
        RECT 157.800 11.400 181.200 12.000 ;
        RECT 187.200 11.400 188.000 12.000 ;
        RECT 187.200 9.600 187.800 11.400 ;
        RECT 188.600 10.800 189.400 15.200 ;
        RECT 166.000 9.400 166.800 9.600 ;
        RECT 161.400 9.000 166.800 9.400 ;
        RECT 160.600 8.800 166.800 9.000 ;
        RECT 167.800 9.000 176.400 9.600 ;
        RECT 158.000 8.000 159.600 8.800 ;
        RECT 160.600 8.200 162.000 8.800 ;
        RECT 167.800 8.200 168.400 9.000 ;
        RECT 175.600 8.800 176.400 9.000 ;
        RECT 178.800 9.000 187.800 9.600 ;
        RECT 178.800 8.800 179.600 9.000 ;
        RECT 159.000 7.600 159.600 8.000 ;
        RECT 162.600 7.600 168.400 8.200 ;
        RECT 169.000 7.600 171.600 8.400 ;
        RECT 156.400 6.800 158.400 7.400 ;
        RECT 159.000 6.800 163.200 7.600 ;
        RECT 145.200 2.200 146.000 5.000 ;
        RECT 146.800 2.200 147.600 5.000 ;
        RECT 150.000 2.200 150.800 6.800 ;
        RECT 153.600 6.200 154.200 6.800 ;
        RECT 153.200 5.600 154.200 6.200 ;
        RECT 157.800 6.200 158.400 6.800 ;
        RECT 157.800 5.600 158.800 6.200 ;
        RECT 153.200 2.200 154.000 5.600 ;
        RECT 158.000 2.200 158.800 5.600 ;
        RECT 161.200 2.200 162.000 6.800 ;
        RECT 164.400 2.200 165.200 5.000 ;
        RECT 166.000 2.200 166.800 5.000 ;
        RECT 167.600 2.200 168.400 7.000 ;
        RECT 170.800 2.200 171.600 7.000 ;
        RECT 174.000 2.200 174.800 8.400 ;
        RECT 182.000 7.600 184.600 8.400 ;
        RECT 177.200 6.800 181.400 7.600 ;
        RECT 175.600 2.200 176.400 5.000 ;
        RECT 177.200 2.200 178.000 5.000 ;
        RECT 178.800 2.200 179.600 5.000 ;
        RECT 182.000 2.200 182.800 7.600 ;
        RECT 187.200 7.400 187.800 9.000 ;
        RECT 185.200 6.800 187.800 7.400 ;
        RECT 188.400 10.000 189.400 10.800 ;
        RECT 199.600 12.300 200.400 19.800 ;
        RECT 202.800 17.600 203.600 19.800 ;
        RECT 201.200 15.600 202.000 17.200 ;
        RECT 203.000 14.400 203.600 17.600 ;
        RECT 206.000 15.800 206.800 19.800 ;
        RECT 210.200 18.400 211.000 19.800 ;
        RECT 210.200 17.600 211.600 18.400 ;
        RECT 210.200 16.800 211.000 17.600 ;
        RECT 210.200 15.800 211.600 16.800 ;
        RECT 206.200 15.600 206.800 15.800 ;
        RECT 206.200 15.200 208.000 15.600 ;
        RECT 206.200 15.000 210.400 15.200 ;
        RECT 207.400 14.600 210.400 15.000 ;
        RECT 209.600 14.400 210.400 14.600 ;
        RECT 202.800 14.300 203.600 14.400 ;
        RECT 206.000 14.300 206.800 14.400 ;
        RECT 202.800 13.700 206.800 14.300 ;
        RECT 208.000 13.800 208.800 14.000 ;
        RECT 202.800 13.600 203.600 13.700 ;
        RECT 201.200 12.300 202.000 12.400 ;
        RECT 199.600 11.700 202.000 12.300 ;
        RECT 185.200 2.200 186.000 6.800 ;
        RECT 188.400 2.200 189.200 10.000 ;
        RECT 199.600 2.200 200.400 11.700 ;
        RECT 201.200 11.600 202.000 11.700 ;
        RECT 203.000 10.200 203.600 13.600 ;
        RECT 206.000 12.800 206.800 13.700 ;
        RECT 207.800 13.200 208.800 13.800 ;
        RECT 207.800 12.400 208.400 13.200 ;
        RECT 204.400 10.800 205.200 12.400 ;
        RECT 207.600 11.600 208.400 12.400 ;
        RECT 209.600 11.000 210.200 14.400 ;
        RECT 211.000 12.400 211.600 15.800 ;
        RECT 210.800 11.600 211.600 12.400 ;
        RECT 207.800 10.400 210.200 11.000 ;
        RECT 202.800 9.400 204.600 10.200 ;
        RECT 203.800 2.200 204.600 9.400 ;
        RECT 207.800 6.200 208.400 10.400 ;
        RECT 211.000 10.200 211.600 11.600 ;
        RECT 207.600 2.200 208.400 6.200 ;
        RECT 210.800 2.200 211.600 10.200 ;
        RECT 212.400 13.800 213.200 19.800 ;
        RECT 218.800 16.600 219.600 19.800 ;
        RECT 220.400 17.000 221.200 19.800 ;
        RECT 222.000 17.000 222.800 19.800 ;
        RECT 223.600 17.000 224.400 19.800 ;
        RECT 226.800 17.000 227.600 19.800 ;
        RECT 230.000 17.000 230.800 19.800 ;
        RECT 231.600 17.000 232.400 19.800 ;
        RECT 233.200 17.000 234.000 19.800 ;
        RECT 234.800 17.000 235.600 19.800 ;
        RECT 217.000 15.800 219.600 16.600 ;
        RECT 236.400 16.600 237.200 19.800 ;
        RECT 223.000 15.800 227.600 16.400 ;
        RECT 217.000 15.200 217.800 15.800 ;
        RECT 214.800 14.400 217.800 15.200 ;
        RECT 212.400 13.000 221.200 13.800 ;
        RECT 223.000 13.400 223.800 15.800 ;
        RECT 226.800 15.600 227.600 15.800 ;
        RECT 228.400 15.600 230.000 16.400 ;
        RECT 233.000 15.600 234.000 16.400 ;
        RECT 236.400 15.800 238.800 16.600 ;
        RECT 225.200 13.600 226.000 15.200 ;
        RECT 226.800 14.800 227.600 15.000 ;
        RECT 226.800 14.200 231.200 14.800 ;
        RECT 230.400 14.000 231.200 14.200 ;
        RECT 212.400 7.400 213.200 13.000 ;
        RECT 221.800 12.600 223.800 13.400 ;
        RECT 227.600 12.600 230.800 13.400 ;
        RECT 233.200 12.800 234.000 15.600 ;
        RECT 238.000 15.200 238.800 15.800 ;
        RECT 238.000 14.600 239.800 15.200 ;
        RECT 239.000 13.400 239.800 14.600 ;
        RECT 242.800 14.600 243.600 19.800 ;
        RECT 244.400 16.000 245.200 19.800 ;
        RECT 247.600 16.000 248.400 19.800 ;
        RECT 250.800 16.000 251.600 19.800 ;
        RECT 244.400 15.200 245.400 16.000 ;
        RECT 247.600 15.800 251.600 16.000 ;
        RECT 252.400 15.800 253.200 19.800 ;
        RECT 247.800 15.400 251.400 15.800 ;
        RECT 242.800 14.000 244.000 14.600 ;
        RECT 239.000 12.600 242.800 13.400 ;
        RECT 213.800 12.000 214.600 12.200 ;
        RECT 215.600 12.000 216.400 12.400 ;
        RECT 218.800 12.000 219.600 12.400 ;
        RECT 236.400 12.000 237.200 12.600 ;
        RECT 243.400 12.000 244.000 14.000 ;
        RECT 213.800 11.400 237.200 12.000 ;
        RECT 243.200 11.400 244.000 12.000 ;
        RECT 243.200 9.600 243.800 11.400 ;
        RECT 244.600 10.800 245.400 15.200 ;
        RECT 252.400 14.400 253.000 15.800 ;
        RECT 250.600 13.600 253.200 14.400 ;
        RECT 249.200 11.600 250.000 13.200 ;
        RECT 222.000 9.400 222.800 9.600 ;
        RECT 217.400 9.000 222.800 9.400 ;
        RECT 216.600 8.800 222.800 9.000 ;
        RECT 223.800 9.000 232.400 9.600 ;
        RECT 214.000 8.000 215.600 8.800 ;
        RECT 216.600 8.200 218.000 8.800 ;
        RECT 223.800 8.200 224.400 9.000 ;
        RECT 231.600 8.800 232.400 9.000 ;
        RECT 234.800 9.000 243.800 9.600 ;
        RECT 234.800 8.800 235.600 9.000 ;
        RECT 215.000 7.600 215.600 8.000 ;
        RECT 218.600 7.600 224.400 8.200 ;
        RECT 225.000 7.600 227.600 8.400 ;
        RECT 212.400 6.800 214.400 7.400 ;
        RECT 215.000 6.800 219.200 7.600 ;
        RECT 213.800 6.200 214.400 6.800 ;
        RECT 213.800 5.600 214.800 6.200 ;
        RECT 214.000 2.200 214.800 5.600 ;
        RECT 217.200 2.200 218.000 6.800 ;
        RECT 220.400 2.200 221.200 5.000 ;
        RECT 222.000 2.200 222.800 5.000 ;
        RECT 223.600 2.200 224.400 7.000 ;
        RECT 226.800 2.200 227.600 7.000 ;
        RECT 230.000 2.200 230.800 8.400 ;
        RECT 238.000 7.600 240.600 8.400 ;
        RECT 233.200 6.800 237.400 7.600 ;
        RECT 231.600 2.200 232.400 5.000 ;
        RECT 233.200 2.200 234.000 5.000 ;
        RECT 234.800 2.200 235.600 5.000 ;
        RECT 238.000 2.200 238.800 7.600 ;
        RECT 243.200 7.400 243.800 9.000 ;
        RECT 241.200 6.800 243.800 7.400 ;
        RECT 244.400 10.000 245.400 10.800 ;
        RECT 250.600 10.200 251.200 13.600 ;
        RECT 241.200 2.200 242.000 6.800 ;
        RECT 244.400 2.200 245.200 10.000 ;
        RECT 250.200 9.600 251.200 10.200 ;
        RECT 250.200 2.200 251.000 9.600 ;
      LAYER via1 ;
        RECT 7.600 175.600 8.400 176.400 ;
        RECT 23.600 175.600 24.400 176.400 ;
        RECT 25.200 174.200 26.000 175.000 ;
        RECT 47.600 177.600 48.400 178.400 ;
        RECT 34.800 171.600 35.600 172.400 ;
        RECT 18.800 166.800 19.600 167.600 ;
        RECT 22.000 166.200 22.800 167.000 ;
        RECT 17.200 164.200 18.000 165.000 ;
        RECT 18.800 164.200 19.600 165.000 ;
        RECT 20.400 164.200 21.200 165.000 ;
        RECT 25.200 166.200 26.000 167.000 ;
        RECT 28.400 166.200 29.200 167.000 ;
        RECT 44.400 171.600 45.200 172.400 ;
        RECT 49.200 173.600 50.000 174.400 ;
        RECT 50.800 171.600 51.600 172.400 ;
        RECT 71.600 173.000 72.400 173.800 ;
        RECT 30.000 164.200 30.800 165.000 ;
        RECT 31.600 164.200 32.400 165.000 ;
        RECT 81.200 172.600 82.000 173.400 ;
        RECT 66.800 171.600 67.600 172.400 ;
        RECT 73.200 168.800 74.000 169.600 ;
        RECT 78.000 167.600 78.800 168.400 ;
        RECT 74.800 166.200 75.600 167.000 ;
        RECT 71.600 164.200 72.400 165.000 ;
        RECT 73.200 164.200 74.000 165.000 ;
        RECT 78.000 166.200 78.800 167.000 ;
        RECT 81.200 166.200 82.000 167.000 ;
        RECT 82.800 164.200 83.600 165.000 ;
        RECT 84.400 164.200 85.200 165.000 ;
        RECT 86.000 164.200 86.800 165.000 ;
        RECT 95.600 163.600 96.400 164.400 ;
        RECT 126.000 175.600 126.800 176.400 ;
        RECT 127.600 174.200 128.400 175.000 ;
        RECT 138.800 171.600 139.600 172.400 ;
        RECT 110.000 163.600 110.800 164.400 ;
        RECT 121.200 166.800 122.000 167.600 ;
        RECT 124.400 166.200 125.200 167.000 ;
        RECT 119.600 164.200 120.400 165.000 ;
        RECT 121.200 164.200 122.000 165.000 ;
        RECT 122.800 164.200 123.600 165.000 ;
        RECT 127.600 166.200 128.400 167.000 ;
        RECT 130.800 166.200 131.600 167.000 ;
        RECT 161.200 173.000 162.000 173.800 ;
        RECT 132.400 164.200 133.200 165.000 ;
        RECT 134.000 164.200 134.800 165.000 ;
        RECT 170.800 172.600 171.600 173.400 ;
        RECT 166.000 171.600 166.800 172.400 ;
        RECT 207.600 173.000 208.400 173.800 ;
        RECT 162.800 168.800 163.600 169.600 ;
        RECT 167.600 167.600 168.400 168.400 ;
        RECT 164.400 166.200 165.200 167.000 ;
        RECT 161.200 164.200 162.000 165.000 ;
        RECT 162.800 164.200 163.600 165.000 ;
        RECT 167.600 166.200 168.400 167.000 ;
        RECT 170.800 166.200 171.600 167.000 ;
        RECT 172.400 164.200 173.200 165.000 ;
        RECT 174.000 164.200 174.800 165.000 ;
        RECT 175.600 164.200 176.400 165.000 ;
        RECT 217.200 172.600 218.000 173.400 ;
        RECT 202.800 171.600 203.600 172.400 ;
        RECT 209.200 168.800 210.000 169.600 ;
        RECT 214.000 167.600 214.800 168.400 ;
        RECT 210.800 166.200 211.600 167.000 ;
        RECT 207.600 164.200 208.400 165.000 ;
        RECT 209.200 164.200 210.000 165.000 ;
        RECT 214.000 166.200 214.800 167.000 ;
        RECT 217.200 166.200 218.000 167.000 ;
        RECT 218.800 164.200 219.600 165.000 ;
        RECT 220.400 164.200 221.200 165.000 ;
        RECT 222.000 164.200 222.800 165.000 ;
        RECT 231.600 163.600 232.400 164.400 ;
        RECT 18.800 154.400 19.600 155.200 ;
        RECT 22.000 155.000 22.800 155.800 ;
        RECT 17.200 152.400 18.000 153.200 ;
        RECT 7.400 147.600 8.200 148.400 ;
        RECT 26.800 147.600 27.600 148.400 ;
        RECT 23.600 145.600 24.400 146.400 ;
        RECT 17.200 144.200 18.000 145.000 ;
        RECT 18.800 144.200 19.600 145.000 ;
        RECT 20.400 144.200 21.200 145.000 ;
        RECT 22.000 144.200 22.800 145.000 ;
        RECT 25.200 144.200 26.000 145.000 ;
        RECT 28.400 144.200 29.200 145.000 ;
        RECT 30.000 144.200 30.800 145.000 ;
        RECT 31.600 144.200 32.400 145.000 ;
        RECT 41.200 145.600 42.000 146.400 ;
        RECT 42.800 143.600 43.600 144.400 ;
        RECT 62.000 155.000 62.800 155.800 ;
        RECT 58.800 153.600 59.600 154.400 ;
        RECT 63.600 152.400 64.400 153.200 ;
        RECT 90.800 157.600 91.600 158.400 ;
        RECT 122.800 157.600 123.600 158.400 ;
        RECT 52.400 148.200 53.200 149.000 ;
        RECT 62.000 148.600 62.800 149.400 ;
        RECT 57.200 147.600 58.000 148.400 ;
        RECT 52.400 144.200 53.200 145.000 ;
        RECT 54.000 144.200 54.800 145.000 ;
        RECT 55.600 144.200 56.400 145.000 ;
        RECT 58.800 144.200 59.600 145.000 ;
        RECT 62.000 144.200 62.800 145.000 ;
        RECT 63.600 144.200 64.400 145.000 ;
        RECT 65.200 144.200 66.000 145.000 ;
        RECT 66.800 144.200 67.600 145.000 ;
        RECT 76.400 143.600 77.200 144.400 ;
        RECT 92.400 145.600 93.200 146.400 ;
        RECT 103.600 149.600 104.400 150.400 ;
        RECT 106.800 147.600 107.600 148.400 ;
        RECT 100.400 143.600 101.200 144.400 ;
        RECT 111.600 145.600 112.400 146.400 ;
        RECT 118.000 145.600 118.800 146.400 ;
        RECT 132.400 149.600 133.200 150.400 ;
        RECT 137.200 147.600 138.000 148.400 ;
        RECT 130.800 145.600 131.600 146.400 ;
        RECT 159.600 155.000 160.400 155.800 ;
        RECT 156.400 153.600 157.200 154.400 ;
        RECT 161.200 152.400 162.000 153.200 ;
        RECT 166.000 149.600 166.800 150.400 ;
        RECT 150.000 148.200 150.800 149.000 ;
        RECT 159.600 148.600 160.400 149.400 ;
        RECT 154.800 147.600 155.600 148.400 ;
        RECT 150.000 144.200 150.800 145.000 ;
        RECT 151.600 144.200 152.400 145.000 ;
        RECT 153.200 144.200 154.000 145.000 ;
        RECT 156.400 144.200 157.200 145.000 ;
        RECT 159.600 144.200 160.400 145.000 ;
        RECT 161.200 144.200 162.000 145.000 ;
        RECT 162.800 144.200 163.600 145.000 ;
        RECT 164.400 144.200 165.200 145.000 ;
        RECT 180.400 149.600 181.200 150.400 ;
        RECT 183.600 149.600 184.400 150.400 ;
        RECT 174.000 143.600 174.800 144.400 ;
        RECT 198.000 147.600 198.800 148.400 ;
        RECT 210.800 149.600 211.600 150.400 ;
        RECT 212.400 149.600 213.200 150.400 ;
        RECT 221.800 151.800 222.600 152.600 ;
        RECT 244.400 153.600 245.200 154.400 ;
        RECT 207.600 147.600 208.400 148.400 ;
        RECT 233.200 149.600 234.000 150.400 ;
        RECT 218.800 147.600 219.600 148.400 ;
        RECT 206.000 143.600 206.800 144.400 ;
        RECT 221.800 146.200 222.600 147.000 ;
        RECT 234.800 147.600 235.600 148.400 ;
        RECT 249.200 143.600 250.000 144.400 ;
        RECT 7.600 135.600 8.400 136.400 ;
        RECT 23.600 135.600 24.400 136.400 ;
        RECT 25.200 134.200 26.000 135.000 ;
        RECT 34.800 131.600 35.600 132.400 ;
        RECT 18.800 126.800 19.600 127.600 ;
        RECT 22.000 126.200 22.800 127.000 ;
        RECT 17.200 124.200 18.000 125.000 ;
        RECT 18.800 124.200 19.600 125.000 ;
        RECT 20.400 124.200 21.200 125.000 ;
        RECT 25.200 126.200 26.000 127.000 ;
        RECT 28.400 126.200 29.200 127.000 ;
        RECT 30.000 124.200 30.800 125.000 ;
        RECT 31.600 124.200 32.400 125.000 ;
        RECT 50.800 133.600 51.600 134.400 ;
        RECT 58.800 133.600 59.600 134.400 ;
        RECT 74.800 137.600 75.600 138.400 ;
        RECT 78.000 137.600 78.800 138.400 ;
        RECT 42.800 123.600 43.600 124.400 ;
        RECT 76.400 133.600 77.200 134.400 ;
        RECT 90.800 133.000 91.600 133.800 ;
        RECT 78.000 123.600 78.800 124.400 ;
        RECT 100.400 132.600 101.200 133.400 ;
        RECT 114.800 137.600 115.600 138.400 ;
        RECT 119.600 137.600 120.400 138.400 ;
        RECT 106.800 131.600 107.600 132.400 ;
        RECT 92.400 128.800 93.200 129.600 ;
        RECT 97.200 127.600 98.000 128.400 ;
        RECT 94.000 126.200 94.800 127.000 ;
        RECT 90.800 124.200 91.600 125.000 ;
        RECT 92.400 124.200 93.200 125.000 ;
        RECT 97.200 126.200 98.000 127.000 ;
        RECT 100.400 126.200 101.200 127.000 ;
        RECT 102.000 124.200 102.800 125.000 ;
        RECT 103.600 124.200 104.400 125.000 ;
        RECT 105.200 124.200 106.000 125.000 ;
        RECT 135.600 135.600 136.400 136.400 ;
        RECT 137.200 134.200 138.000 135.000 ;
        RECT 146.800 131.600 147.600 132.400 ;
        RECT 130.800 126.800 131.600 127.600 ;
        RECT 134.000 126.200 134.800 127.000 ;
        RECT 129.200 124.200 130.000 125.000 ;
        RECT 130.800 124.200 131.600 125.000 ;
        RECT 132.400 124.200 133.200 125.000 ;
        RECT 137.200 126.200 138.000 127.000 ;
        RECT 140.400 126.200 141.200 127.000 ;
        RECT 154.800 137.600 155.600 138.400 ;
        RECT 142.000 124.200 142.800 125.000 ;
        RECT 143.600 124.200 144.400 125.000 ;
        RECT 161.200 137.600 162.000 138.400 ;
        RECT 159.600 133.600 160.400 134.400 ;
        RECT 164.400 133.600 165.200 134.400 ;
        RECT 193.200 137.600 194.000 138.400 ;
        RECT 180.400 133.600 181.200 134.400 ;
        RECT 191.600 133.600 192.400 134.400 ;
        RECT 207.600 137.600 208.400 138.400 ;
        RECT 174.000 123.600 174.800 124.400 ;
        RECT 199.600 131.600 200.400 132.400 ;
        RECT 199.600 127.600 200.400 128.400 ;
        RECT 206.000 129.600 206.800 130.400 ;
        RECT 218.800 137.600 219.600 138.400 ;
        RECT 220.400 133.600 221.200 134.400 ;
        RECT 236.400 137.600 237.200 138.400 ;
        RECT 222.000 131.600 222.800 132.400 ;
        RECT 214.000 123.600 214.800 124.400 ;
        RECT 236.400 129.600 237.200 130.400 ;
        RECT 242.800 123.600 243.600 124.400 ;
        RECT 249.200 123.600 250.000 124.400 ;
        RECT 18.800 114.400 19.600 115.200 ;
        RECT 22.000 115.000 22.800 115.800 ;
        RECT 17.200 112.400 18.000 113.200 ;
        RECT 7.600 105.600 8.400 106.400 ;
        RECT 26.800 107.600 27.600 108.400 ;
        RECT 23.600 105.600 24.400 106.400 ;
        RECT 17.200 104.200 18.000 105.000 ;
        RECT 18.800 104.200 19.600 105.000 ;
        RECT 20.400 104.200 21.200 105.000 ;
        RECT 22.000 104.200 22.800 105.000 ;
        RECT 25.200 104.200 26.000 105.000 ;
        RECT 28.400 104.200 29.200 105.000 ;
        RECT 30.000 104.200 30.800 105.000 ;
        RECT 31.600 104.200 32.400 105.000 ;
        RECT 63.600 117.600 64.400 118.400 ;
        RECT 54.000 109.600 54.800 110.400 ;
        RECT 55.600 109.600 56.400 110.400 ;
        RECT 47.600 105.600 48.400 106.400 ;
        RECT 44.400 103.600 45.200 104.400 ;
        RECT 78.000 111.800 78.800 112.600 ;
        RECT 78.000 106.200 78.800 107.000 ;
        RECT 89.200 109.600 90.000 110.400 ;
        RECT 92.400 109.600 93.200 110.400 ;
        RECT 113.200 115.000 114.000 115.800 ;
        RECT 110.000 113.600 110.800 114.400 ;
        RECT 127.600 117.600 128.400 118.400 ;
        RECT 114.800 112.400 115.600 113.200 ;
        RECT 119.600 109.600 120.400 110.400 ;
        RECT 86.000 107.600 86.800 108.400 ;
        RECT 90.800 107.600 91.600 108.400 ;
        RECT 82.800 106.400 83.600 107.200 ;
        RECT 94.000 107.600 94.800 108.400 ;
        RECT 103.600 108.200 104.400 109.000 ;
        RECT 113.200 108.600 114.000 109.400 ;
        RECT 108.400 107.600 109.200 108.400 ;
        RECT 103.600 104.200 104.400 105.000 ;
        RECT 105.200 104.200 106.000 105.000 ;
        RECT 106.800 104.200 107.600 105.000 ;
        RECT 110.000 104.200 110.800 105.000 ;
        RECT 113.200 104.200 114.000 105.000 ;
        RECT 114.800 104.200 115.600 105.000 ;
        RECT 116.400 104.200 117.200 105.000 ;
        RECT 118.000 104.200 118.800 105.000 ;
        RECT 140.400 109.600 141.200 110.400 ;
        RECT 145.200 109.600 146.000 110.400 ;
        RECT 151.600 109.600 152.400 110.400 ;
        RECT 154.800 109.600 155.600 110.400 ;
        RECT 142.000 107.600 142.800 108.400 ;
        RECT 153.200 107.600 154.000 108.400 ;
        RECT 156.400 107.600 157.200 108.400 ;
        RECT 167.600 109.600 168.400 110.400 ;
        RECT 169.200 107.600 170.000 108.400 ;
        RECT 159.600 103.600 160.400 104.400 ;
        RECT 170.800 105.600 171.600 106.400 ;
        RECT 175.600 105.600 176.400 106.400 ;
        RECT 182.000 105.600 182.800 106.400 ;
        RECT 206.000 109.600 206.800 110.400 ;
        RECT 226.800 115.000 227.600 115.800 ;
        RECT 223.600 113.600 224.400 114.400 ;
        RECT 228.400 112.400 229.200 113.200 ;
        RECT 204.400 107.600 205.200 108.400 ;
        RECT 198.000 105.600 198.800 106.400 ;
        RECT 194.800 103.600 195.600 104.400 ;
        RECT 207.600 107.600 208.400 108.400 ;
        RECT 217.200 108.200 218.000 109.000 ;
        RECT 226.800 108.600 227.600 109.400 ;
        RECT 222.000 107.600 222.800 108.400 ;
        RECT 217.200 104.200 218.000 105.000 ;
        RECT 218.800 104.200 219.600 105.000 ;
        RECT 220.400 104.200 221.200 105.000 ;
        RECT 223.600 104.200 224.400 105.000 ;
        RECT 226.800 104.200 227.600 105.000 ;
        RECT 228.400 104.200 229.200 105.000 ;
        RECT 230.000 104.200 230.800 105.000 ;
        RECT 231.600 104.200 232.400 105.000 ;
        RECT 247.600 109.600 248.400 110.400 ;
        RECT 241.200 103.600 242.000 104.400 ;
        RECT 23.600 95.600 24.400 96.400 ;
        RECT 25.200 94.200 26.000 95.000 ;
        RECT 54.000 97.600 54.800 98.400 ;
        RECT 36.400 91.600 37.200 92.400 ;
        RECT 7.600 89.600 8.400 90.400 ;
        RECT 18.800 86.800 19.600 87.600 ;
        RECT 22.000 86.200 22.800 87.000 ;
        RECT 17.200 84.200 18.000 85.000 ;
        RECT 18.800 84.200 19.600 85.000 ;
        RECT 20.400 84.200 21.200 85.000 ;
        RECT 25.200 86.200 26.000 87.000 ;
        RECT 28.400 86.200 29.200 87.000 ;
        RECT 41.200 93.600 42.000 94.400 ;
        RECT 55.600 94.800 56.400 95.600 ;
        RECT 58.800 93.600 59.600 94.400 ;
        RECT 78.000 97.600 78.800 98.400 ;
        RECT 62.000 93.600 62.800 94.400 ;
        RECT 30.000 84.200 30.800 85.000 ;
        RECT 31.600 84.200 32.400 85.000 ;
        RECT 98.800 95.600 99.600 96.400 ;
        RECT 100.400 94.200 101.200 95.000 ;
        RECT 90.800 91.600 91.600 92.400 ;
        RECT 113.200 91.600 114.000 92.400 ;
        RECT 78.000 83.600 78.800 84.400 ;
        RECT 94.000 86.800 94.800 87.600 ;
        RECT 97.200 86.200 98.000 87.000 ;
        RECT 92.400 84.200 93.200 85.000 ;
        RECT 94.000 84.200 94.800 85.000 ;
        RECT 95.600 84.200 96.400 85.000 ;
        RECT 100.400 86.200 101.200 87.000 ;
        RECT 103.600 86.200 104.400 87.000 ;
        RECT 124.400 93.000 125.200 93.800 ;
        RECT 134.000 92.600 134.800 93.400 ;
        RECT 148.400 97.600 149.200 98.400 ;
        RECT 119.600 91.600 120.400 92.400 ;
        RECT 126.000 88.800 126.800 89.600 ;
        RECT 130.800 87.600 131.600 88.400 ;
        RECT 105.200 84.200 106.000 85.000 ;
        RECT 106.800 84.200 107.600 85.000 ;
        RECT 127.600 86.200 128.400 87.000 ;
        RECT 124.400 84.200 125.200 85.000 ;
        RECT 126.000 84.200 126.800 85.000 ;
        RECT 130.800 86.200 131.600 87.000 ;
        RECT 134.000 86.200 134.800 87.000 ;
        RECT 135.600 84.200 136.400 85.000 ;
        RECT 137.200 84.200 138.000 85.000 ;
        RECT 138.800 84.200 139.600 85.000 ;
        RECT 182.000 97.600 182.800 98.400 ;
        RECT 148.400 83.600 149.200 84.400 ;
        RECT 169.200 91.600 170.000 92.400 ;
        RECT 169.200 87.600 170.000 88.400 ;
        RECT 175.600 89.600 176.400 90.400 ;
        RECT 196.400 89.600 197.200 90.400 ;
        RECT 191.600 83.600 192.400 84.400 ;
        RECT 206.000 89.600 206.800 90.400 ;
        RECT 214.000 89.600 214.800 90.400 ;
        RECT 210.800 87.600 211.600 88.400 ;
        RECT 226.800 97.600 227.600 98.400 ;
        RECT 225.200 93.600 226.000 94.400 ;
        RECT 218.800 91.600 219.600 92.400 ;
        RECT 234.800 93.600 235.600 94.400 ;
        RECT 247.600 97.600 248.400 98.400 ;
        RECT 241.200 93.600 242.000 94.400 ;
        RECT 249.200 93.600 250.000 94.400 ;
        RECT 17.200 77.600 18.000 78.400 ;
        RECT 36.400 73.600 37.200 74.400 ;
        RECT 4.400 69.600 5.200 70.400 ;
        RECT 34.800 65.600 35.600 66.400 ;
        RECT 31.600 63.600 32.400 64.400 ;
        RECT 39.600 69.600 40.400 70.400 ;
        RECT 42.800 69.600 43.600 70.400 ;
        RECT 46.000 69.600 46.800 70.400 ;
        RECT 47.600 69.600 48.400 70.400 ;
        RECT 76.400 77.600 77.200 78.400 ;
        RECT 79.600 77.600 80.400 78.400 ;
        RECT 52.400 67.600 53.200 68.400 ;
        RECT 55.600 67.600 56.400 68.400 ;
        RECT 42.800 63.600 43.600 64.400 ;
        RECT 47.600 63.600 48.400 64.400 ;
        RECT 57.200 67.600 58.000 68.400 ;
        RECT 82.800 69.600 83.600 70.400 ;
        RECT 102.000 75.000 102.800 75.800 ;
        RECT 98.800 73.600 99.600 74.400 ;
        RECT 116.400 77.600 117.200 78.400 ;
        RECT 103.600 72.400 104.400 73.200 ;
        RECT 108.400 69.600 109.200 70.400 ;
        RECT 92.400 68.200 93.200 69.000 ;
        RECT 102.000 68.600 102.800 69.400 ;
        RECT 97.200 67.600 98.000 68.400 ;
        RECT 92.400 64.200 93.200 65.000 ;
        RECT 94.000 64.200 94.800 65.000 ;
        RECT 95.600 64.200 96.400 65.000 ;
        RECT 98.800 64.200 99.600 65.000 ;
        RECT 102.000 64.200 102.800 65.000 ;
        RECT 103.600 64.200 104.400 65.000 ;
        RECT 105.200 64.200 106.000 65.000 ;
        RECT 106.800 64.200 107.600 65.000 ;
        RECT 129.200 77.600 130.000 78.400 ;
        RECT 126.000 69.600 126.800 70.400 ;
        RECT 145.200 69.600 146.000 70.400 ;
        RECT 151.600 69.600 152.400 70.400 ;
        RECT 135.600 67.600 136.400 68.400 ;
        RECT 138.800 67.600 139.600 68.400 ;
        RECT 148.400 63.600 149.200 64.400 ;
        RECT 154.800 63.600 155.600 64.400 ;
        RECT 161.200 65.600 162.000 66.400 ;
        RECT 166.000 67.600 166.800 68.400 ;
        RECT 169.200 65.600 170.000 66.400 ;
        RECT 174.000 65.600 174.800 66.400 ;
        RECT 202.800 75.000 203.600 75.800 ;
        RECT 199.600 73.600 200.400 74.400 ;
        RECT 217.200 77.600 218.000 78.400 ;
        RECT 204.400 72.400 205.200 73.200 ;
        RECT 209.200 69.600 210.000 70.400 ;
        RECT 193.200 68.200 194.000 69.000 ;
        RECT 202.800 68.600 203.600 69.400 ;
        RECT 198.000 67.600 198.800 68.400 ;
        RECT 193.200 64.200 194.000 65.000 ;
        RECT 194.800 64.200 195.600 65.000 ;
        RECT 196.400 64.200 197.200 65.000 ;
        RECT 199.600 64.200 200.400 65.000 ;
        RECT 202.800 64.200 203.600 65.000 ;
        RECT 204.400 64.200 205.200 65.000 ;
        RECT 206.000 64.200 206.800 65.000 ;
        RECT 207.600 64.200 208.400 65.000 ;
        RECT 233.400 71.800 234.200 72.600 ;
        RECT 246.000 73.600 246.800 74.400 ;
        RECT 228.400 69.600 229.200 70.400 ;
        RECT 234.600 69.800 235.400 70.600 ;
        RECT 242.800 71.600 243.600 72.400 ;
        RECT 217.200 63.600 218.000 64.400 ;
        RECT 223.600 63.600 224.400 64.400 ;
        RECT 230.000 65.600 230.800 66.400 ;
        RECT 233.400 66.200 234.200 67.000 ;
        RECT 7.600 57.600 8.400 58.400 ;
        RECT 26.800 55.600 27.600 56.400 ;
        RECT 28.400 54.200 29.200 55.000 ;
        RECT 46.000 57.600 46.800 58.400 ;
        RECT 38.000 51.600 38.800 52.400 ;
        RECT 39.600 51.600 40.400 52.400 ;
        RECT 22.000 46.800 22.800 47.600 ;
        RECT 25.200 46.200 26.000 47.000 ;
        RECT 20.400 44.200 21.200 45.000 ;
        RECT 22.000 44.200 22.800 45.000 ;
        RECT 23.600 44.200 24.400 45.000 ;
        RECT 28.400 46.200 29.200 47.000 ;
        RECT 31.600 46.200 32.400 47.000 ;
        RECT 62.000 55.600 62.800 56.400 ;
        RECT 63.600 54.200 64.400 55.000 ;
        RECT 54.000 51.600 54.800 52.400 ;
        RECT 74.800 51.600 75.600 52.400 ;
        RECT 33.200 44.200 34.000 45.000 ;
        RECT 34.800 44.200 35.600 45.000 ;
        RECT 57.200 46.800 58.000 47.600 ;
        RECT 60.400 46.200 61.200 47.000 ;
        RECT 55.600 44.200 56.400 45.000 ;
        RECT 57.200 44.200 58.000 45.000 ;
        RECT 58.800 44.200 59.600 45.000 ;
        RECT 63.600 46.200 64.400 47.000 ;
        RECT 66.800 46.200 67.600 47.000 ;
        RECT 90.800 57.600 91.600 58.400 ;
        RECT 100.400 51.600 101.200 52.400 ;
        RECT 113.200 53.000 114.000 53.800 ;
        RECT 68.400 44.200 69.200 45.000 ;
        RECT 70.000 44.200 70.800 45.000 ;
        RECT 98.800 43.600 99.600 44.400 ;
        RECT 122.800 52.600 123.600 53.400 ;
        RECT 137.200 55.600 138.000 56.400 ;
        RECT 108.400 51.600 109.200 52.400 ;
        RECT 114.800 48.800 115.600 49.600 ;
        RECT 119.600 47.600 120.400 48.400 ;
        RECT 116.400 46.200 117.200 47.000 ;
        RECT 113.200 44.200 114.000 45.000 ;
        RECT 114.800 44.200 115.600 45.000 ;
        RECT 119.600 46.200 120.400 47.000 ;
        RECT 122.800 46.200 123.600 47.000 ;
        RECT 124.400 44.200 125.200 45.000 ;
        RECT 126.000 44.200 126.800 45.000 ;
        RECT 127.600 44.200 128.400 45.000 ;
        RECT 153.200 57.600 154.000 58.400 ;
        RECT 169.200 55.600 170.000 56.400 ;
        RECT 170.800 54.200 171.600 55.000 ;
        RECT 172.400 51.600 173.200 52.400 ;
        RECT 164.400 46.800 165.200 47.600 ;
        RECT 167.600 46.200 168.400 47.000 ;
        RECT 162.800 44.200 163.600 45.000 ;
        RECT 164.400 44.200 165.200 45.000 ;
        RECT 166.000 44.200 166.800 45.000 ;
        RECT 170.800 46.200 171.600 47.000 ;
        RECT 174.000 46.200 174.800 47.000 ;
        RECT 175.600 44.200 176.400 45.000 ;
        RECT 177.200 44.200 178.000 45.000 ;
        RECT 201.200 51.600 202.000 52.400 ;
        RECT 196.400 49.600 197.200 50.400 ;
        RECT 217.200 53.000 218.000 53.800 ;
        RECT 207.600 49.600 208.400 50.400 ;
        RECT 226.800 52.600 227.600 53.400 ;
        RECT 241.200 57.600 242.000 58.400 ;
        RECT 214.000 51.600 214.800 52.400 ;
        RECT 250.800 57.600 251.600 58.400 ;
        RECT 218.800 48.800 219.600 49.600 ;
        RECT 223.600 47.600 224.400 48.400 ;
        RECT 220.400 46.200 221.200 47.000 ;
        RECT 217.200 44.200 218.000 45.000 ;
        RECT 218.800 44.200 219.600 45.000 ;
        RECT 223.600 46.200 224.400 47.000 ;
        RECT 226.800 46.200 227.600 47.000 ;
        RECT 228.400 44.200 229.200 45.000 ;
        RECT 230.000 44.200 230.800 45.000 ;
        RECT 231.600 44.200 232.400 45.000 ;
        RECT 249.200 49.600 250.000 50.400 ;
        RECT 18.800 34.400 19.600 35.200 ;
        RECT 22.000 35.000 22.800 35.800 ;
        RECT 17.200 32.400 18.000 33.200 ;
        RECT 7.600 25.600 8.400 26.400 ;
        RECT 26.800 27.600 27.600 28.400 ;
        RECT 23.600 25.600 24.400 26.400 ;
        RECT 17.200 24.200 18.000 25.000 ;
        RECT 18.800 24.200 19.600 25.000 ;
        RECT 20.400 24.200 21.200 25.000 ;
        RECT 22.000 24.200 22.800 25.000 ;
        RECT 25.200 24.200 26.000 25.000 ;
        RECT 28.400 24.200 29.200 25.000 ;
        RECT 30.000 24.200 30.800 25.000 ;
        RECT 31.600 24.200 32.400 25.000 ;
        RECT 47.600 25.600 48.400 26.400 ;
        RECT 55.600 29.600 56.400 30.400 ;
        RECT 81.200 35.000 82.000 35.800 ;
        RECT 78.000 33.600 78.800 34.400 ;
        RECT 82.800 32.400 83.600 33.200 ;
        RECT 71.600 28.200 72.400 29.000 ;
        RECT 81.200 28.600 82.000 29.400 ;
        RECT 52.400 23.600 53.200 24.400 ;
        RECT 76.400 27.600 77.200 28.400 ;
        RECT 71.600 24.200 72.400 25.000 ;
        RECT 73.200 24.200 74.000 25.000 ;
        RECT 74.800 24.200 75.600 25.000 ;
        RECT 78.000 24.200 78.800 25.000 ;
        RECT 81.200 24.200 82.000 25.000 ;
        RECT 82.800 24.200 83.600 25.000 ;
        RECT 84.400 24.200 85.200 25.000 ;
        RECT 86.000 24.200 86.800 25.000 ;
        RECT 121.200 37.600 122.000 38.400 ;
        RECT 95.600 23.600 96.400 24.400 ;
        RECT 143.600 29.600 144.400 30.400 ;
        RECT 146.800 27.600 147.600 28.400 ;
        RECT 140.400 23.600 141.200 24.400 ;
        RECT 166.000 35.000 166.800 35.800 ;
        RECT 162.800 33.600 163.600 34.400 ;
        RECT 167.600 32.400 168.400 33.200 ;
        RECT 172.400 29.600 173.200 30.400 ;
        RECT 156.400 28.200 157.200 29.000 ;
        RECT 166.000 28.600 166.800 29.400 ;
        RECT 161.200 27.600 162.000 28.400 ;
        RECT 180.600 27.600 181.400 28.400 ;
        RECT 156.400 24.200 157.200 25.000 ;
        RECT 158.000 24.200 158.800 25.000 ;
        RECT 159.600 24.200 160.400 25.000 ;
        RECT 162.800 24.200 163.600 25.000 ;
        RECT 166.000 24.200 166.800 25.000 ;
        RECT 167.600 24.200 168.400 25.000 ;
        RECT 169.200 24.200 170.000 25.000 ;
        RECT 170.800 24.200 171.600 25.000 ;
        RECT 193.200 29.600 194.000 30.400 ;
        RECT 194.800 25.600 195.600 26.400 ;
        RECT 198.000 23.600 198.800 24.400 ;
        RECT 225.200 35.000 226.000 35.800 ;
        RECT 222.000 33.600 222.800 34.400 ;
        RECT 239.600 37.600 240.400 38.400 ;
        RECT 226.800 32.400 227.600 33.200 ;
        RECT 210.800 31.600 211.600 32.400 ;
        RECT 214.000 31.200 214.800 32.000 ;
        RECT 242.800 37.600 243.600 38.400 ;
        RECT 215.600 28.200 216.400 29.000 ;
        RECT 225.200 28.600 226.000 29.400 ;
        RECT 206.000 25.600 206.800 26.400 ;
        RECT 220.400 27.600 221.200 28.400 ;
        RECT 215.600 24.200 216.400 25.000 ;
        RECT 217.200 24.200 218.000 25.000 ;
        RECT 218.800 24.200 219.600 25.000 ;
        RECT 222.000 24.200 222.800 25.000 ;
        RECT 225.200 24.200 226.000 25.000 ;
        RECT 226.800 24.200 227.600 25.000 ;
        RECT 228.400 24.200 229.200 25.000 ;
        RECT 230.000 24.200 230.800 25.000 ;
        RECT 246.000 29.600 246.800 30.400 ;
        RECT 7.400 13.600 8.200 14.400 ;
        RECT 23.600 15.600 24.400 16.400 ;
        RECT 25.200 14.200 26.000 15.000 ;
        RECT 36.400 11.600 37.200 12.400 ;
        RECT 18.800 6.800 19.600 7.600 ;
        RECT 22.000 6.200 22.800 7.000 ;
        RECT 17.200 4.200 18.000 5.000 ;
        RECT 18.800 4.200 19.600 5.000 ;
        RECT 20.400 4.200 21.200 5.000 ;
        RECT 25.200 6.200 26.000 7.000 ;
        RECT 28.400 6.200 29.200 7.000 ;
        RECT 44.400 11.600 45.200 12.400 ;
        RECT 66.800 13.000 67.600 13.800 ;
        RECT 50.800 11.600 51.600 12.400 ;
        RECT 30.000 4.200 30.800 5.000 ;
        RECT 31.600 4.200 32.400 5.000 ;
        RECT 76.400 12.600 77.200 13.400 ;
        RECT 63.600 11.600 64.400 12.400 ;
        RECT 100.400 17.600 101.200 18.400 ;
        RECT 91.000 13.600 91.800 14.400 ;
        RECT 68.400 8.800 69.200 9.600 ;
        RECT 73.200 7.600 74.000 8.400 ;
        RECT 70.000 6.200 70.800 7.000 ;
        RECT 66.800 4.200 67.600 5.000 ;
        RECT 68.400 4.200 69.200 5.000 ;
        RECT 73.200 6.200 74.000 7.000 ;
        RECT 76.400 6.200 77.200 7.000 ;
        RECT 78.000 4.200 78.800 5.000 ;
        RECT 79.600 4.200 80.400 5.000 ;
        RECT 81.200 4.200 82.000 5.000 ;
        RECT 122.600 11.600 123.400 12.400 ;
        RECT 138.800 15.600 139.600 16.400 ;
        RECT 140.400 14.200 141.200 15.000 ;
        RECT 151.600 11.600 152.400 12.400 ;
        RECT 119.600 9.600 120.400 10.400 ;
        RECT 134.000 6.800 134.800 7.600 ;
        RECT 137.200 6.200 138.000 7.000 ;
        RECT 132.400 4.200 133.200 5.000 ;
        RECT 134.000 4.200 134.800 5.000 ;
        RECT 135.600 4.200 136.400 5.000 ;
        RECT 140.400 6.200 141.200 7.000 ;
        RECT 143.600 6.200 144.400 7.000 ;
        RECT 164.400 13.000 165.200 13.800 ;
        RECT 174.000 12.600 174.800 13.400 ;
        RECT 188.400 15.600 189.200 16.400 ;
        RECT 159.600 11.600 160.400 12.400 ;
        RECT 166.000 8.800 166.800 9.600 ;
        RECT 170.800 7.600 171.600 8.400 ;
        RECT 145.200 4.200 146.000 5.000 ;
        RECT 146.800 4.200 147.600 5.000 ;
        RECT 167.600 6.200 168.400 7.000 ;
        RECT 164.400 4.200 165.200 5.000 ;
        RECT 166.000 4.200 166.800 5.000 ;
        RECT 170.800 6.200 171.600 7.000 ;
        RECT 174.000 6.200 174.800 7.000 ;
        RECT 175.600 4.200 176.400 5.000 ;
        RECT 177.200 4.200 178.000 5.000 ;
        RECT 178.800 4.200 179.600 5.000 ;
        RECT 210.800 17.600 211.600 18.400 ;
        RECT 204.400 11.600 205.200 12.400 ;
        RECT 220.400 13.000 221.200 13.800 ;
        RECT 230.000 12.600 230.800 13.400 ;
        RECT 252.400 17.600 253.200 18.400 ;
        RECT 215.600 11.600 216.400 12.400 ;
        RECT 222.000 8.800 222.800 9.600 ;
        RECT 226.800 7.600 227.600 8.400 ;
        RECT 223.600 6.200 224.400 7.000 ;
        RECT 220.400 4.200 221.200 5.000 ;
        RECT 222.000 4.200 222.800 5.000 ;
        RECT 226.800 6.200 227.600 7.000 ;
        RECT 230.000 6.200 230.800 7.000 ;
        RECT 231.600 4.200 232.400 5.000 ;
        RECT 233.200 4.200 234.000 5.000 ;
        RECT 234.800 4.200 235.600 5.000 ;
        RECT 244.400 9.600 245.200 10.400 ;
      LAYER metal2 ;
        RECT 7.600 175.600 8.400 176.400 ;
        RECT 17.200 164.200 18.000 177.800 ;
        RECT 18.800 164.200 19.600 177.800 ;
        RECT 20.400 164.200 21.200 177.800 ;
        RECT 22.000 166.200 22.800 177.800 ;
        RECT 23.600 175.600 24.400 176.400 ;
        RECT 7.400 147.600 8.400 148.400 ;
        RECT 17.200 144.200 18.000 157.800 ;
        RECT 18.800 144.200 19.600 157.800 ;
        RECT 20.400 144.200 21.200 157.800 ;
        RECT 22.000 144.200 22.800 155.800 ;
        RECT 23.700 146.400 24.300 175.600 ;
        RECT 25.200 166.200 26.000 177.800 ;
        RECT 26.800 177.600 27.600 178.400 ;
        RECT 26.900 174.400 27.500 177.600 ;
        RECT 26.800 173.600 27.600 174.400 ;
        RECT 28.400 166.200 29.200 177.800 ;
        RECT 30.000 164.200 30.800 177.800 ;
        RECT 31.600 164.200 32.400 177.800 ;
        RECT 47.600 177.600 48.400 178.400 ;
        RECT 41.200 175.600 42.000 176.400 ;
        RECT 44.400 173.600 45.200 174.400 ;
        RECT 49.200 173.600 50.000 174.400 ;
        RECT 44.500 172.400 45.100 173.600 ;
        RECT 34.800 171.600 35.600 172.400 ;
        RECT 44.400 171.600 45.200 172.400 ;
        RECT 50.800 171.600 51.600 172.400 ;
        RECT 55.600 171.600 56.400 172.400 ;
        RECT 66.800 171.600 67.600 172.400 ;
        RECT 23.600 145.600 24.400 146.400 ;
        RECT 7.600 135.600 8.400 136.400 ;
        RECT 17.200 124.200 18.000 137.800 ;
        RECT 18.800 124.200 19.600 137.800 ;
        RECT 20.400 124.200 21.200 137.800 ;
        RECT 22.000 126.200 22.800 137.800 ;
        RECT 23.700 136.400 24.300 145.600 ;
        RECT 25.200 144.200 26.000 155.800 ;
        RECT 26.800 147.600 27.600 148.400 ;
        RECT 26.900 142.400 27.500 147.600 ;
        RECT 28.400 144.200 29.200 155.800 ;
        RECT 30.000 144.200 30.800 157.800 ;
        RECT 31.600 144.200 32.400 157.800 ;
        RECT 34.900 150.400 35.500 171.600 ;
        RECT 34.800 149.600 35.600 150.400 ;
        RECT 26.800 141.600 27.600 142.400 ;
        RECT 23.600 135.600 24.400 136.400 ;
        RECT 7.600 105.600 8.400 106.400 ;
        RECT 17.200 104.200 18.000 117.800 ;
        RECT 18.800 104.200 19.600 117.800 ;
        RECT 20.400 104.200 21.200 117.800 ;
        RECT 22.000 104.200 22.800 115.800 ;
        RECT 23.700 106.400 24.300 135.600 ;
        RECT 25.200 126.200 26.000 137.800 ;
        RECT 26.800 133.600 27.600 134.400 ;
        RECT 28.400 126.200 29.200 137.800 ;
        RECT 30.000 124.200 30.800 137.800 ;
        RECT 31.600 124.200 32.400 137.800 ;
        RECT 34.900 132.400 35.500 149.600 ;
        RECT 41.200 147.600 42.000 148.400 ;
        RECT 41.300 146.400 41.900 147.600 ;
        RECT 41.200 145.600 42.000 146.400 ;
        RECT 42.800 143.600 43.600 144.400 ;
        RECT 42.900 136.400 43.500 143.600 ;
        RECT 41.200 135.600 42.000 136.400 ;
        RECT 42.800 135.600 43.600 136.400 ;
        RECT 34.800 131.600 35.600 132.400 ;
        RECT 23.600 105.600 24.400 106.400 ;
        RECT 7.600 89.600 8.400 90.400 ;
        RECT 17.200 84.200 18.000 97.800 ;
        RECT 18.800 84.200 19.600 97.800 ;
        RECT 20.400 84.200 21.200 97.800 ;
        RECT 22.000 86.200 22.800 97.800 ;
        RECT 23.700 96.400 24.300 105.600 ;
        RECT 25.200 104.200 26.000 115.800 ;
        RECT 26.800 107.600 27.600 108.400 ;
        RECT 26.900 104.400 27.500 107.600 ;
        RECT 26.800 103.600 27.600 104.400 ;
        RECT 28.400 104.200 29.200 115.800 ;
        RECT 30.000 104.200 30.800 117.800 ;
        RECT 31.600 104.200 32.400 117.800 ;
        RECT 34.900 110.400 35.500 131.600 ;
        RECT 44.500 124.400 45.100 171.600 ;
        RECT 50.900 150.400 51.500 171.600 ;
        RECT 55.700 158.400 56.300 171.600 ;
        RECT 71.600 164.200 72.400 177.800 ;
        RECT 73.200 164.200 74.000 177.800 ;
        RECT 74.800 166.200 75.600 177.800 ;
        RECT 76.400 173.600 77.200 174.400 ;
        RECT 78.000 166.200 78.800 177.800 ;
        RECT 79.600 175.600 80.400 176.400 ;
        RECT 47.600 149.600 48.400 150.400 ;
        RECT 50.800 149.600 51.600 150.400 ;
        RECT 50.800 143.600 51.600 144.400 ;
        RECT 52.400 144.200 53.200 157.800 ;
        RECT 54.000 144.200 54.800 157.800 ;
        RECT 55.600 157.600 56.400 158.400 ;
        RECT 55.600 144.200 56.400 155.800 ;
        RECT 57.200 147.600 58.000 148.400 ;
        RECT 50.900 136.400 51.500 143.600 ;
        RECT 57.300 142.400 57.900 147.600 ;
        RECT 58.800 144.200 59.600 155.800 ;
        RECT 60.400 145.600 61.200 146.400 ;
        RECT 62.000 144.200 62.800 155.800 ;
        RECT 63.600 144.200 64.400 157.800 ;
        RECT 65.200 144.200 66.000 157.800 ;
        RECT 66.800 144.200 67.600 157.800 ;
        RECT 68.400 157.600 69.200 158.400 ;
        RECT 55.600 141.600 56.400 142.400 ;
        RECT 57.200 141.600 58.000 142.400 ;
        RECT 50.800 135.600 51.600 136.400 ;
        RECT 50.900 134.400 51.500 135.600 ;
        RECT 55.700 134.400 56.300 141.600 ;
        RECT 68.500 138.400 69.100 157.600 ;
        RECT 70.000 149.600 70.800 150.400 ;
        RECT 68.400 137.600 69.200 138.400 ;
        RECT 68.500 136.400 69.100 137.600 ;
        RECT 68.400 135.600 69.200 136.400 ;
        RECT 70.100 134.400 70.700 149.600 ;
        RECT 78.000 147.600 78.800 148.400 ;
        RECT 76.400 143.600 77.200 144.400 ;
        RECT 74.800 141.600 75.600 142.400 ;
        RECT 74.900 138.400 75.500 141.600 ;
        RECT 76.500 138.400 77.100 143.600 ;
        RECT 78.100 138.400 78.700 147.600 ;
        RECT 74.800 137.600 75.600 138.400 ;
        RECT 76.400 137.600 77.200 138.400 ;
        RECT 78.000 137.600 78.800 138.400 ;
        RECT 79.700 134.400 80.300 175.600 ;
        RECT 81.200 166.200 82.000 177.800 ;
        RECT 82.800 164.200 83.600 177.800 ;
        RECT 84.400 164.200 85.200 177.800 ;
        RECT 86.000 164.200 86.800 177.800 ;
        RECT 90.800 173.600 91.600 174.400 ;
        RECT 90.900 158.400 91.500 173.600 ;
        RECT 95.600 163.600 96.400 164.400 ;
        RECT 110.000 163.600 110.800 164.400 ;
        RECT 118.000 163.600 118.800 164.400 ;
        RECT 119.600 164.200 120.400 177.800 ;
        RECT 121.200 164.200 122.000 177.800 ;
        RECT 122.800 164.200 123.600 177.800 ;
        RECT 124.400 166.200 125.200 177.800 ;
        RECT 126.000 175.600 126.800 176.400 ;
        RECT 127.600 166.200 128.400 177.800 ;
        RECT 129.200 173.600 130.000 174.400 ;
        RECT 90.800 157.600 91.600 158.400 ;
        RECT 86.000 149.600 86.800 150.400 ;
        RECT 84.400 137.600 85.200 138.400 ;
        RECT 47.600 133.600 48.400 134.400 ;
        RECT 50.800 133.600 51.600 134.400 ;
        RECT 55.600 133.600 56.400 134.400 ;
        RECT 58.800 133.600 59.600 134.400 ;
        RECT 70.000 133.600 70.800 134.400 ;
        RECT 76.400 133.600 77.200 134.400 ;
        RECT 79.600 133.600 80.400 134.400 ;
        RECT 46.000 131.600 46.800 132.400 ;
        RECT 49.200 131.600 50.000 132.400 ;
        RECT 54.000 131.600 54.800 132.400 ;
        RECT 57.200 132.300 58.000 132.400 ;
        RECT 55.700 131.700 58.000 132.300 ;
        RECT 42.800 123.600 43.600 124.400 ;
        RECT 44.400 123.600 45.200 124.400 ;
        RECT 42.900 110.400 43.500 123.600 ;
        RECT 34.800 109.600 35.600 110.400 ;
        RECT 36.400 109.600 37.200 110.400 ;
        RECT 41.200 109.600 42.000 110.400 ;
        RECT 42.800 109.600 43.600 110.400 ;
        RECT 23.600 95.600 24.400 96.400 ;
        RECT 23.700 82.400 24.300 95.600 ;
        RECT 25.200 86.200 26.000 97.800 ;
        RECT 26.800 93.600 27.600 94.400 ;
        RECT 28.400 86.200 29.200 97.800 ;
        RECT 30.000 84.200 30.800 97.800 ;
        RECT 31.600 84.200 32.400 97.800 ;
        RECT 36.500 92.400 37.100 109.600 ;
        RECT 41.300 94.400 41.900 109.600 ;
        RECT 42.800 107.600 43.600 108.400 ;
        RECT 44.400 103.600 45.200 104.400 ;
        RECT 42.800 95.600 43.600 96.400 ;
        RECT 44.400 95.600 45.200 96.400 ;
        RECT 42.900 94.400 43.500 95.600 ;
        RECT 41.200 93.600 42.000 94.400 ;
        RECT 42.800 93.600 43.600 94.400 ;
        RECT 36.400 91.600 37.200 92.400 ;
        RECT 17.200 81.600 18.000 82.400 ;
        RECT 23.600 81.600 24.400 82.400 ;
        RECT 17.300 78.400 17.900 81.600 ;
        RECT 17.200 77.600 18.000 78.400 ;
        RECT 41.300 74.400 41.900 93.600 ;
        RECT 42.800 91.600 43.600 92.400 ;
        RECT 36.400 73.600 37.200 74.400 ;
        RECT 41.200 73.600 42.000 74.400 ;
        RECT 7.600 71.600 8.400 72.400 ;
        RECT 38.000 71.600 38.800 72.400 ;
        RECT 4.400 69.600 5.200 70.400 ;
        RECT 4.500 62.400 5.100 69.600 ;
        RECT 4.400 61.600 5.200 62.400 ;
        RECT 7.700 58.400 8.300 71.600 ;
        RECT 38.100 68.400 38.700 71.600 ;
        RECT 42.900 70.400 43.500 91.600 ;
        RECT 39.600 69.600 40.400 70.400 ;
        RECT 42.800 69.600 43.600 70.400 ;
        RECT 42.900 68.400 43.500 69.600 ;
        RECT 44.500 68.400 45.100 95.600 ;
        RECT 46.100 92.400 46.700 131.600 ;
        RECT 49.300 130.400 49.900 131.600 ;
        RECT 49.200 129.600 50.000 130.400 ;
        RECT 50.800 123.600 51.600 124.400 ;
        RECT 50.900 110.400 51.500 123.600 ;
        RECT 52.400 111.600 53.200 112.400 ;
        RECT 50.800 109.600 51.600 110.400 ;
        RECT 50.900 108.400 51.500 109.600 ;
        RECT 52.500 108.400 53.100 111.600 ;
        RECT 55.700 110.400 56.300 131.700 ;
        RECT 57.200 131.600 58.000 131.700 ;
        RECT 58.900 118.400 59.500 133.600 ;
        RECT 62.000 131.600 62.800 132.400 ;
        RECT 74.800 131.600 75.600 132.400 ;
        RECT 74.900 130.400 75.500 131.600 ;
        RECT 74.800 129.600 75.600 130.400 ;
        RECT 62.000 127.600 62.800 128.400 ;
        RECT 58.800 117.600 59.600 118.400 ;
        RECT 57.200 111.600 58.000 112.400 ;
        RECT 60.400 111.600 61.200 112.400 ;
        RECT 54.000 109.600 54.800 110.400 ;
        RECT 55.600 109.600 56.400 110.400 ;
        RECT 54.100 108.400 54.700 109.600 ;
        RECT 50.800 107.600 51.600 108.400 ;
        RECT 52.400 107.600 53.200 108.400 ;
        RECT 54.000 107.600 54.800 108.400 ;
        RECT 47.600 105.600 48.400 106.400 ;
        RECT 54.100 98.400 54.700 107.600 ;
        RECT 57.300 106.400 57.900 111.600 ;
        RECT 60.500 110.400 61.100 111.600 ;
        RECT 60.400 109.600 61.200 110.400 ;
        RECT 58.800 107.600 59.600 108.400 ;
        RECT 57.200 105.600 58.000 106.400 ;
        RECT 60.400 105.600 61.200 106.400 ;
        RECT 54.000 97.600 54.800 98.400 ;
        RECT 50.800 95.000 51.600 95.800 ;
        RECT 57.000 95.600 57.800 95.800 ;
        RECT 52.200 95.000 57.800 95.600 ;
        RECT 47.600 93.600 48.400 94.400 ;
        RECT 49.200 93.600 50.000 94.400 ;
        RECT 50.800 94.200 51.400 95.000 ;
        RECT 52.200 94.800 53.000 95.000 ;
        RECT 55.600 94.800 56.400 95.000 ;
        RECT 50.800 93.600 56.400 94.200 ;
        RECT 46.000 91.600 46.800 92.400 ;
        RECT 46.000 71.600 46.800 72.400 ;
        RECT 46.100 70.400 46.700 71.600 ;
        RECT 46.000 69.600 46.800 70.400 ;
        RECT 47.600 69.600 48.400 70.400 ;
        RECT 47.700 68.400 48.300 69.600 ;
        RECT 38.000 67.600 38.800 68.400 ;
        RECT 42.800 67.600 43.600 68.400 ;
        RECT 44.400 67.600 45.200 68.400 ;
        RECT 47.600 67.600 48.400 68.400 ;
        RECT 34.800 65.600 35.600 66.400 ;
        RECT 31.600 63.600 32.400 64.400 ;
        RECT 31.700 60.400 32.300 63.600 ;
        RECT 34.900 62.400 35.500 65.600 ;
        RECT 34.800 61.600 35.600 62.400 ;
        RECT 26.800 59.600 27.600 60.400 ;
        RECT 31.600 59.600 32.400 60.400 ;
        RECT 7.600 57.600 8.400 58.400 ;
        RECT 6.000 55.600 6.800 56.400 ;
        RECT 9.200 55.600 10.000 56.400 ;
        RECT 6.100 52.400 6.700 55.600 ;
        RECT 6.000 51.600 6.800 52.400 ;
        RECT 20.400 44.200 21.200 57.800 ;
        RECT 22.000 44.200 22.800 57.800 ;
        RECT 23.600 44.200 24.400 57.800 ;
        RECT 25.200 46.200 26.000 57.800 ;
        RECT 26.900 56.400 27.500 59.600 ;
        RECT 26.800 55.600 27.600 56.400 ;
        RECT 7.600 25.600 8.400 26.400 ;
        RECT 17.200 24.200 18.000 37.800 ;
        RECT 18.800 24.200 19.600 37.800 ;
        RECT 20.400 24.200 21.200 37.800 ;
        RECT 22.000 24.200 22.800 35.800 ;
        RECT 23.600 29.600 24.400 30.400 ;
        RECT 23.700 26.400 24.300 29.600 ;
        RECT 23.600 25.600 24.400 26.400 ;
        RECT 7.400 13.600 8.400 14.400 ;
        RECT 17.200 4.200 18.000 17.800 ;
        RECT 18.800 4.200 19.600 17.800 ;
        RECT 20.400 4.200 21.200 17.800 ;
        RECT 22.000 6.200 22.800 17.800 ;
        RECT 23.700 16.400 24.300 25.600 ;
        RECT 25.200 24.200 26.000 35.800 ;
        RECT 26.900 30.400 27.500 55.600 ;
        RECT 28.400 46.200 29.200 57.800 ;
        RECT 30.000 55.600 30.800 56.400 ;
        RECT 30.100 54.400 30.700 55.600 ;
        RECT 30.000 53.600 30.800 54.400 ;
        RECT 31.600 46.200 32.400 57.800 ;
        RECT 33.200 44.200 34.000 57.800 ;
        RECT 34.800 44.200 35.600 57.800 ;
        RECT 38.100 54.400 38.700 67.600 ;
        RECT 42.800 63.600 43.600 64.400 ;
        RECT 42.900 56.400 43.500 63.600 ;
        RECT 42.800 55.600 43.600 56.400 ;
        RECT 38.000 53.600 38.800 54.400 ;
        RECT 38.000 51.600 38.800 52.400 ;
        RECT 39.600 51.600 40.400 52.400 ;
        RECT 26.800 29.600 27.600 30.400 ;
        RECT 26.800 27.600 27.600 28.400 ;
        RECT 28.400 24.200 29.200 35.800 ;
        RECT 30.000 24.200 30.800 37.800 ;
        RECT 31.600 24.200 32.400 37.800 ;
        RECT 36.400 30.300 37.200 30.400 ;
        RECT 38.100 30.300 38.700 51.600 ;
        RECT 44.500 32.400 45.100 67.600 ;
        RECT 47.600 63.600 48.400 64.400 ;
        RECT 46.000 61.600 46.800 62.400 ;
        RECT 46.100 58.400 46.700 61.600 ;
        RECT 46.000 57.600 46.800 58.400 ;
        RECT 47.700 54.400 48.300 63.600 ;
        RECT 49.300 62.400 49.900 93.600 ;
        RECT 50.800 90.200 51.400 93.600 ;
        RECT 52.400 91.600 53.200 92.400 ;
        RECT 55.800 92.200 56.400 93.600 ;
        RECT 50.800 89.400 51.600 90.200 ;
        RECT 52.500 86.400 53.100 91.600 ;
        RECT 55.800 91.400 56.600 92.200 ;
        RECT 57.200 90.200 57.800 95.000 ;
        RECT 58.800 93.600 59.600 94.400 ;
        RECT 58.900 90.400 59.500 93.600 ;
        RECT 57.000 89.400 57.800 90.200 ;
        RECT 58.800 89.600 59.600 90.400 ;
        RECT 52.400 85.600 53.200 86.400 ;
        RECT 50.800 73.600 51.600 74.400 ;
        RECT 50.900 68.300 51.500 73.600 ;
        RECT 52.500 70.400 53.100 85.600 ;
        RECT 60.500 74.400 61.100 105.600 ;
        RECT 62.100 94.400 62.700 127.600 ;
        RECT 63.600 117.600 64.400 118.400 ;
        RECT 74.900 110.400 75.500 129.600 ;
        RECT 76.500 122.400 77.100 133.600 ;
        RECT 81.200 131.600 82.000 132.400 ;
        RECT 78.000 123.600 78.800 124.400 ;
        RECT 76.400 121.600 77.200 122.400 ;
        RECT 84.500 116.300 85.100 137.600 ;
        RECT 86.100 128.400 86.700 149.600 ;
        RECT 95.700 148.400 96.300 163.600 ;
        RECT 97.200 149.600 98.000 150.400 ;
        RECT 103.600 149.600 104.400 150.400 ;
        RECT 111.600 149.600 112.400 150.400 ;
        RECT 92.400 147.600 93.200 148.400 ;
        RECT 95.600 147.600 96.400 148.400 ;
        RECT 92.500 146.400 93.100 147.600 ;
        RECT 92.400 145.600 93.200 146.400 ;
        RECT 97.300 144.400 97.900 149.600 ;
        RECT 98.800 147.600 99.600 148.400 ;
        RECT 106.800 147.600 107.600 148.400 ;
        RECT 111.700 146.400 112.300 149.600 ;
        RECT 118.100 146.400 118.700 163.600 ;
        RECT 129.300 162.400 129.900 173.600 ;
        RECT 130.800 166.200 131.600 177.800 ;
        RECT 130.800 163.600 131.600 164.400 ;
        RECT 132.400 164.200 133.200 177.800 ;
        RECT 134.000 164.200 134.800 177.800 ;
        RECT 158.000 175.600 158.800 176.400 ;
        RECT 138.800 171.600 139.600 172.400 ;
        RECT 143.600 171.600 144.400 172.400 ;
        RECT 148.400 171.600 149.200 172.400 ;
        RECT 122.800 161.600 123.600 162.400 ;
        RECT 129.200 161.600 130.000 162.400 ;
        RECT 122.900 158.400 123.500 161.600 ;
        RECT 122.800 157.600 123.600 158.400 ;
        RECT 119.600 149.600 120.400 150.400 ;
        RECT 121.200 149.600 122.000 150.400 ;
        RECT 127.600 149.600 128.400 150.400 ;
        RECT 102.000 145.600 102.800 146.400 ;
        RECT 108.400 145.600 109.200 146.400 ;
        RECT 111.600 145.600 112.400 146.400 ;
        RECT 118.000 145.600 118.800 146.400 ;
        RECT 97.200 143.600 98.000 144.400 ;
        RECT 100.400 143.600 101.200 144.400 ;
        RECT 100.500 140.400 101.100 143.600 ;
        RECT 95.600 139.600 96.400 140.400 ;
        RECT 100.400 139.600 101.200 140.400 ;
        RECT 86.000 127.600 86.800 128.400 ;
        RECT 90.800 124.200 91.600 137.800 ;
        RECT 92.400 124.200 93.200 137.800 ;
        RECT 94.000 126.200 94.800 137.800 ;
        RECT 95.700 134.400 96.300 139.600 ;
        RECT 111.700 138.400 112.300 145.600 ;
        RECT 119.700 138.400 120.300 149.600 ;
        RECT 121.300 148.400 121.900 149.600 ;
        RECT 121.200 147.600 122.000 148.400 ;
        RECT 126.000 147.600 126.800 148.400 ;
        RECT 95.600 133.600 96.400 134.400 ;
        RECT 97.200 126.200 98.000 137.800 ;
        RECT 98.800 135.600 99.600 136.400 ;
        RECT 98.900 130.400 99.500 135.600 ;
        RECT 98.800 129.600 99.600 130.400 ;
        RECT 100.400 126.200 101.200 137.800 ;
        RECT 102.000 124.200 102.800 137.800 ;
        RECT 103.600 124.200 104.400 137.800 ;
        RECT 105.200 124.200 106.000 137.800 ;
        RECT 111.600 137.600 112.400 138.400 ;
        RECT 114.800 137.600 115.600 138.400 ;
        RECT 119.600 137.600 120.400 138.400 ;
        RECT 111.600 135.600 112.400 136.400 ;
        RECT 106.800 131.600 107.600 132.400 ;
        RECT 106.900 126.300 107.500 131.600 ;
        RECT 111.700 130.400 112.300 135.600 ;
        RECT 111.600 129.600 112.400 130.400 ;
        RECT 106.900 125.700 109.100 126.300 ;
        RECT 94.000 121.600 94.800 122.400 ;
        RECT 84.500 115.700 86.700 116.300 ;
        RECT 78.000 111.800 78.800 112.600 ;
        RECT 71.600 109.600 72.400 110.400 ;
        RECT 74.800 109.600 75.600 110.400 ;
        RECT 62.000 93.600 62.800 94.400 ;
        RECT 71.700 92.400 72.300 109.600 ;
        RECT 78.000 108.400 78.600 111.800 ;
        RECT 79.600 111.600 80.400 112.400 ;
        RECT 84.600 111.800 85.400 112.600 ;
        RECT 82.000 108.400 82.800 108.600 ;
        RECT 76.400 107.600 77.200 108.400 ;
        RECT 78.000 107.800 82.800 108.400 ;
        RECT 74.800 101.600 75.600 102.400 ;
        RECT 73.200 93.600 74.000 94.400 ;
        RECT 74.900 92.400 75.500 101.600 ;
        RECT 76.500 100.400 77.100 107.600 ;
        RECT 78.000 107.000 78.600 107.800 ;
        RECT 79.400 107.000 80.200 107.200 ;
        RECT 82.800 107.000 83.600 107.200 ;
        RECT 84.800 107.000 85.400 111.800 ;
        RECT 86.100 108.400 86.700 115.700 ;
        RECT 89.200 109.600 90.000 110.400 ;
        RECT 92.400 109.600 93.200 110.400 ;
        RECT 86.000 107.600 86.800 108.400 ;
        RECT 87.600 107.600 88.400 108.400 ;
        RECT 90.800 107.600 91.600 108.400 ;
        RECT 78.000 106.200 78.800 107.000 ;
        RECT 79.400 106.400 83.600 107.000 ;
        RECT 84.600 106.200 85.400 107.000 ;
        RECT 87.700 104.400 88.300 107.600 ;
        RECT 78.000 103.600 78.800 104.400 ;
        RECT 87.600 103.600 88.400 104.400 ;
        RECT 76.400 99.600 77.200 100.400 ;
        RECT 78.100 98.400 78.700 103.600 ;
        RECT 92.500 102.400 93.100 109.600 ;
        RECT 94.100 108.400 94.700 121.600 ;
        RECT 94.000 107.600 94.800 108.400 ;
        RECT 103.600 104.200 104.400 117.800 ;
        RECT 105.200 104.200 106.000 117.800 ;
        RECT 106.800 104.200 107.600 115.800 ;
        RECT 108.500 110.400 109.100 125.700 ;
        RECT 108.400 109.600 109.200 110.400 ;
        RECT 108.400 107.600 109.200 108.400 ;
        RECT 110.000 104.200 110.800 115.800 ;
        RECT 111.700 106.400 112.300 129.600 ;
        RECT 127.700 122.400 128.300 149.600 ;
        RECT 130.900 146.400 131.500 163.600 ;
        RECT 138.900 156.400 139.500 171.600 ;
        RECT 143.700 164.400 144.300 171.600 ;
        RECT 148.500 170.400 149.100 171.600 ;
        RECT 148.400 169.600 149.200 170.400 ;
        RECT 143.600 163.600 144.400 164.400 ;
        RECT 138.800 155.600 139.600 156.400 ;
        RECT 146.800 155.600 147.600 156.400 ;
        RECT 140.400 151.600 141.200 152.400 ;
        RECT 132.400 149.600 133.200 150.400 ;
        RECT 137.200 149.600 138.000 150.400 ;
        RECT 137.300 148.400 137.900 149.600 ;
        RECT 137.200 147.600 138.000 148.400 ;
        RECT 130.800 145.600 131.600 146.400 ;
        RECT 130.900 140.400 131.500 145.600 ;
        RECT 138.800 143.600 139.600 144.400 ;
        RECT 130.800 139.600 131.600 140.400 ;
        RECT 129.200 124.200 130.000 137.800 ;
        RECT 130.800 124.200 131.600 137.800 ;
        RECT 132.400 124.200 133.200 137.800 ;
        RECT 134.000 126.200 134.800 137.800 ;
        RECT 135.600 135.600 136.400 136.400 ;
        RECT 135.600 133.600 136.400 134.400 ;
        RECT 127.600 121.600 128.400 122.400 ;
        RECT 111.600 105.600 112.400 106.400 ;
        RECT 92.400 101.600 93.200 102.400 ;
        RECT 79.600 99.600 80.400 100.400 ;
        RECT 76.400 97.600 77.200 98.400 ;
        RECT 78.000 97.600 78.800 98.400 ;
        RECT 71.600 91.600 72.400 92.400 ;
        RECT 74.800 91.600 75.600 92.400 ;
        RECT 57.200 73.600 58.000 74.400 ;
        RECT 60.400 73.600 61.200 74.400 ;
        RECT 52.400 69.600 53.200 70.400 ;
        RECT 57.300 68.400 57.900 73.600 ;
        RECT 71.700 68.400 72.300 91.600 ;
        RECT 74.900 86.400 75.500 91.600 ;
        RECT 74.800 85.600 75.600 86.400 ;
        RECT 76.500 78.400 77.100 97.600 ;
        RECT 79.700 96.400 80.300 99.600 ;
        RECT 111.700 98.400 112.300 105.600 ;
        RECT 113.200 104.200 114.000 115.800 ;
        RECT 114.800 104.200 115.600 117.800 ;
        RECT 116.400 104.200 117.200 117.800 ;
        RECT 118.000 104.200 118.800 117.800 ;
        RECT 127.600 117.600 128.400 118.400 ;
        RECT 135.700 112.400 136.300 133.600 ;
        RECT 137.200 126.200 138.000 137.800 ;
        RECT 138.900 136.400 139.500 143.600 ;
        RECT 140.500 140.400 141.100 151.600 ;
        RECT 146.900 150.400 147.500 155.600 ;
        RECT 146.800 149.600 147.600 150.400 ;
        RECT 140.400 139.600 141.200 140.400 ;
        RECT 138.800 135.600 139.600 136.400 ;
        RECT 138.800 133.600 139.600 134.400 ;
        RECT 135.600 111.600 136.400 112.400 ;
        RECT 138.900 110.400 139.500 133.600 ;
        RECT 140.400 126.200 141.200 137.800 ;
        RECT 142.000 124.200 142.800 137.800 ;
        RECT 143.600 124.200 144.400 137.800 ;
        RECT 146.900 132.400 147.500 149.600 ;
        RECT 150.000 144.200 150.800 157.800 ;
        RECT 151.600 144.200 152.400 157.800 ;
        RECT 153.200 144.200 154.000 155.800 ;
        RECT 154.800 147.600 155.600 148.400 ;
        RECT 154.900 142.400 155.500 147.600 ;
        RECT 156.400 144.200 157.200 155.800 ;
        RECT 158.100 146.400 158.700 175.600 ;
        RECT 161.200 164.200 162.000 177.800 ;
        RECT 162.800 164.200 163.600 177.800 ;
        RECT 164.400 166.200 165.200 177.800 ;
        RECT 166.000 173.600 166.800 174.400 ;
        RECT 166.000 171.600 166.800 172.400 ;
        RECT 158.000 145.600 158.800 146.400 ;
        RECT 159.600 144.200 160.400 155.800 ;
        RECT 161.200 144.200 162.000 157.800 ;
        RECT 162.800 144.200 163.600 157.800 ;
        RECT 164.400 144.200 165.200 157.800 ;
        RECT 166.100 150.400 166.700 171.600 ;
        RECT 167.600 166.200 168.400 177.800 ;
        RECT 169.200 175.600 170.000 176.400 ;
        RECT 170.800 166.200 171.600 177.800 ;
        RECT 172.400 164.200 173.200 177.800 ;
        RECT 174.000 164.200 174.800 177.800 ;
        RECT 175.600 164.200 176.400 177.800 ;
        RECT 183.600 173.600 184.400 174.400 ;
        RECT 183.700 158.400 184.300 173.600 ;
        RECT 194.800 171.600 195.600 172.400 ;
        RECT 202.800 171.600 203.600 172.400 ;
        RECT 194.900 160.400 195.500 171.600 ;
        RECT 207.600 164.200 208.400 177.800 ;
        RECT 209.200 164.200 210.000 177.800 ;
        RECT 210.800 166.200 211.600 177.800 ;
        RECT 212.400 173.600 213.200 174.400 ;
        RECT 194.800 159.600 195.600 160.400 ;
        RECT 198.000 159.600 198.800 160.400 ;
        RECT 183.600 157.600 184.400 158.400 ;
        RECT 194.800 151.600 195.600 152.400 ;
        RECT 166.000 149.600 166.800 150.400 ;
        RECT 174.000 149.600 174.800 150.400 ;
        RECT 180.400 149.600 181.200 150.400 ;
        RECT 183.600 149.600 184.400 150.400 ;
        RECT 193.200 149.600 194.000 150.400 ;
        RECT 174.100 144.400 174.700 149.600 ;
        RECT 180.400 147.600 181.200 148.400 ;
        RECT 182.000 147.600 182.800 148.400 ;
        RECT 175.600 145.600 176.400 146.400 ;
        RECT 170.800 143.600 171.600 144.400 ;
        RECT 174.000 143.600 174.800 144.400 ;
        RECT 154.800 141.600 155.600 142.400 ;
        RECT 161.200 141.600 162.000 142.400 ;
        RECT 154.800 139.600 155.600 140.400 ;
        RECT 154.900 138.400 155.500 139.600 ;
        RECT 161.300 138.400 161.900 141.600 ;
        RECT 154.800 137.600 155.600 138.400 ;
        RECT 158.000 137.600 158.800 138.400 ;
        RECT 161.200 137.600 162.000 138.400 ;
        RECT 158.100 132.400 158.700 137.600 ;
        RECT 162.800 135.600 163.600 136.400 ;
        RECT 166.000 135.600 166.800 136.400 ;
        RECT 170.900 134.400 171.500 143.600 ;
        RECT 175.700 134.400 176.300 145.600 ;
        RECT 180.500 134.400 181.100 147.600 ;
        RECT 182.100 146.400 182.700 147.600 ;
        RECT 182.000 145.600 182.800 146.400 ;
        RECT 182.000 139.600 182.800 140.400 ;
        RECT 159.600 133.600 160.400 134.400 ;
        RECT 164.400 133.600 165.200 134.400 ;
        RECT 170.800 133.600 171.600 134.400 ;
        RECT 175.600 133.600 176.400 134.400 ;
        RECT 177.200 133.600 178.000 134.400 ;
        RECT 180.400 133.600 181.200 134.400 ;
        RECT 146.800 131.600 147.600 132.400 ;
        RECT 158.000 131.600 158.800 132.400 ;
        RECT 119.600 109.600 120.400 110.400 ;
        RECT 130.800 109.600 131.600 110.400 ;
        RECT 134.000 109.600 134.800 110.400 ;
        RECT 135.600 109.600 136.400 110.400 ;
        RECT 138.800 109.600 139.600 110.400 ;
        RECT 140.400 109.600 141.200 110.400 ;
        RECT 145.200 109.600 146.000 110.400 ;
        RECT 116.400 99.600 117.200 100.400 ;
        RECT 79.600 95.600 80.400 96.400 ;
        RECT 79.600 91.600 80.400 92.400 ;
        RECT 90.800 91.600 91.600 92.400 ;
        RECT 78.000 83.600 78.800 84.400 ;
        RECT 76.400 77.600 77.200 78.400 ;
        RECT 52.400 68.300 53.200 68.400 ;
        RECT 50.900 67.700 53.200 68.300 ;
        RECT 52.400 67.600 53.200 67.700 ;
        RECT 55.600 67.600 56.400 68.400 ;
        RECT 57.200 67.600 58.000 68.400 ;
        RECT 71.600 67.600 72.400 68.400 ;
        RECT 49.200 61.600 50.000 62.400 ;
        RECT 62.000 59.600 62.800 60.400 ;
        RECT 46.000 53.600 46.800 54.400 ;
        RECT 47.600 53.600 48.400 54.400 ;
        RECT 44.400 31.600 45.200 32.400 ;
        RECT 46.100 30.400 46.700 53.600 ;
        RECT 54.000 51.600 54.800 52.400 ;
        RECT 55.600 44.200 56.400 57.800 ;
        RECT 57.200 44.200 58.000 57.800 ;
        RECT 58.800 44.200 59.600 57.800 ;
        RECT 60.400 46.200 61.200 57.800 ;
        RECT 62.100 56.400 62.700 59.600 ;
        RECT 62.000 55.600 62.800 56.400 ;
        RECT 50.800 31.600 51.600 32.400 ;
        RECT 36.400 29.700 38.700 30.300 ;
        RECT 36.400 29.600 37.200 29.700 ;
        RECT 41.200 29.600 42.000 30.400 ;
        RECT 46.000 29.600 46.800 30.400 ;
        RECT 47.600 29.600 48.400 30.400 ;
        RECT 23.600 15.600 24.400 16.400 ;
        RECT 25.200 6.200 26.000 17.800 ;
        RECT 26.800 15.600 27.600 16.400 ;
        RECT 26.900 14.400 27.500 15.600 ;
        RECT 26.800 13.600 27.600 14.400 ;
        RECT 28.400 6.200 29.200 17.800 ;
        RECT 30.000 4.200 30.800 17.800 ;
        RECT 31.600 4.200 32.400 17.800 ;
        RECT 36.500 12.400 37.100 29.600 ;
        RECT 41.300 26.400 41.900 29.600 ;
        RECT 42.800 27.600 43.600 28.400 ;
        RECT 44.400 27.600 45.200 28.400 ;
        RECT 41.200 25.600 42.000 26.400 ;
        RECT 41.200 15.600 42.000 16.400 ;
        RECT 41.300 14.400 41.900 15.600 ;
        RECT 41.200 13.600 42.000 14.400 ;
        RECT 44.500 12.400 45.100 27.600 ;
        RECT 47.600 25.600 48.400 26.400 ;
        RECT 47.600 15.600 48.400 16.400 ;
        RECT 50.900 12.400 51.500 31.600 ;
        RECT 55.600 29.600 56.400 30.400 ;
        RECT 62.100 26.400 62.700 55.600 ;
        RECT 63.600 46.200 64.400 57.800 ;
        RECT 65.200 53.600 66.000 54.400 ;
        RECT 66.800 46.200 67.600 57.800 ;
        RECT 68.400 44.200 69.200 57.800 ;
        RECT 70.000 44.200 70.800 57.800 ;
        RECT 74.800 51.600 75.600 52.400 ;
        RECT 76.400 51.600 77.200 52.400 ;
        RECT 65.200 29.600 66.000 30.400 ;
        RECT 62.000 25.600 62.800 26.400 ;
        RECT 52.400 23.600 53.200 24.400 ;
        RECT 52.500 14.400 53.100 23.600 ;
        RECT 52.400 13.600 53.200 14.400 ;
        RECT 65.300 14.300 65.900 29.600 ;
        RECT 71.600 24.200 72.400 37.800 ;
        RECT 73.200 24.200 74.000 37.800 ;
        RECT 74.800 24.200 75.600 35.800 ;
        RECT 76.500 30.400 77.100 51.600 ;
        RECT 78.100 38.400 78.700 83.600 ;
        RECT 79.700 78.400 80.300 91.600 ;
        RECT 79.600 77.600 80.400 78.400 ;
        RECT 90.900 70.400 91.500 91.600 ;
        RECT 92.400 84.200 93.200 97.800 ;
        RECT 94.000 84.200 94.800 97.800 ;
        RECT 95.600 84.200 96.400 97.800 ;
        RECT 97.200 86.200 98.000 97.800 ;
        RECT 98.800 97.600 99.600 98.400 ;
        RECT 98.900 96.400 99.500 97.600 ;
        RECT 98.800 95.600 99.600 96.400 ;
        RECT 98.900 84.300 99.500 95.600 ;
        RECT 100.400 86.200 101.200 97.800 ;
        RECT 102.000 93.600 102.800 94.400 ;
        RECT 103.600 86.200 104.400 97.800 ;
        RECT 98.900 83.700 101.100 84.300 ;
        RECT 105.200 84.200 106.000 97.800 ;
        RECT 106.800 84.200 107.600 97.800 ;
        RECT 111.600 97.600 112.400 98.400 ;
        RECT 113.200 91.600 114.000 92.400 ;
        RECT 82.800 69.600 83.600 70.400 ;
        RECT 90.800 69.600 91.600 70.400 ;
        RECT 79.600 53.600 80.400 54.400 ;
        RECT 79.700 52.400 80.300 53.600 ;
        RECT 82.900 52.400 83.500 69.600 ;
        RECT 90.900 58.400 91.500 69.600 ;
        RECT 92.400 64.200 93.200 77.800 ;
        RECT 94.000 64.200 94.800 77.800 ;
        RECT 95.600 64.200 96.400 75.800 ;
        RECT 97.200 75.600 98.000 76.400 ;
        RECT 97.300 68.400 97.900 75.600 ;
        RECT 97.200 67.600 98.000 68.400 ;
        RECT 98.800 64.200 99.600 75.800 ;
        RECT 100.500 66.400 101.100 83.700 ;
        RECT 116.500 78.400 117.100 99.600 ;
        RECT 119.700 92.400 120.300 109.600 ;
        RECT 130.900 106.400 131.500 109.600 ;
        RECT 134.100 108.400 134.700 109.600 ;
        RECT 135.700 108.400 136.300 109.600 ;
        RECT 134.000 107.600 134.800 108.400 ;
        RECT 135.600 107.600 136.400 108.400 ;
        RECT 130.800 105.600 131.600 106.400 ;
        RECT 129.200 103.600 130.000 104.400 ;
        RECT 119.600 91.600 120.400 92.400 ;
        RECT 124.400 84.200 125.200 97.800 ;
        RECT 126.000 84.200 126.800 97.800 ;
        RECT 127.600 86.200 128.400 97.800 ;
        RECT 129.300 94.400 129.900 103.600 ;
        RECT 140.500 102.400 141.100 109.600 ;
        RECT 142.000 107.600 142.800 108.400 ;
        RECT 143.600 107.600 144.400 108.400 ;
        RECT 142.100 106.300 142.700 107.600 ;
        RECT 142.100 105.700 144.300 106.300 ;
        RECT 140.400 101.600 141.200 102.400 ;
        RECT 129.200 93.600 130.000 94.400 ;
        RECT 129.200 91.600 130.000 92.400 ;
        RECT 129.300 78.400 129.900 91.600 ;
        RECT 130.800 86.200 131.600 97.800 ;
        RECT 132.400 97.600 133.200 98.400 ;
        RECT 132.500 96.400 133.100 97.600 ;
        RECT 132.400 95.600 133.200 96.400 ;
        RECT 134.000 86.200 134.800 97.800 ;
        RECT 135.600 84.200 136.400 97.800 ;
        RECT 137.200 84.200 138.000 97.800 ;
        RECT 138.800 84.200 139.600 97.800 ;
        RECT 142.000 83.600 142.800 84.400 ;
        RECT 100.400 65.600 101.200 66.400 ;
        RECT 102.000 64.200 102.800 75.800 ;
        RECT 103.600 64.200 104.400 77.800 ;
        RECT 105.200 64.200 106.000 77.800 ;
        RECT 106.800 64.200 107.600 77.800 ;
        RECT 116.400 77.600 117.200 78.400 ;
        RECT 124.400 77.600 125.200 78.400 ;
        RECT 129.200 77.600 130.000 78.400 ;
        RECT 116.500 72.400 117.100 77.600 ;
        RECT 116.400 71.600 117.200 72.400 ;
        RECT 122.800 71.600 123.600 72.400 ;
        RECT 122.900 70.400 123.500 71.600 ;
        RECT 108.400 69.600 109.200 70.400 ;
        RECT 118.000 69.600 118.800 70.400 ;
        RECT 122.800 69.600 123.600 70.400 ;
        RECT 90.800 57.600 91.600 58.400 ;
        RECT 103.600 55.600 104.400 56.400 ;
        RECT 103.700 54.400 104.300 55.600 ;
        RECT 95.600 53.600 96.400 54.400 ;
        RECT 102.000 53.600 102.800 54.400 ;
        RECT 103.600 53.600 104.400 54.400 ;
        RECT 95.700 52.400 96.300 53.600 ;
        RECT 108.500 52.400 109.100 69.600 ;
        RECT 79.600 51.600 80.400 52.400 ;
        RECT 82.800 51.600 83.600 52.400 ;
        RECT 89.200 51.600 90.000 52.400 ;
        RECT 94.000 51.600 94.800 52.400 ;
        RECT 95.600 51.600 96.400 52.400 ;
        RECT 100.400 51.600 101.200 52.400 ;
        RECT 108.400 51.600 109.200 52.400 ;
        RECT 78.000 37.600 78.800 38.400 ;
        RECT 76.400 29.600 77.200 30.400 ;
        RECT 76.400 27.600 77.200 28.400 ;
        RECT 78.000 24.200 78.800 35.800 ;
        RECT 79.600 25.600 80.400 26.400 ;
        RECT 79.700 20.400 80.300 25.600 ;
        RECT 81.200 24.200 82.000 35.800 ;
        RECT 82.800 24.200 83.600 37.800 ;
        RECT 84.400 24.200 85.200 37.800 ;
        RECT 86.000 24.200 86.800 37.800 ;
        RECT 74.800 19.600 75.600 20.400 ;
        RECT 79.600 19.600 80.400 20.400 ;
        RECT 63.700 13.700 65.900 14.300 ;
        RECT 52.500 12.400 53.100 13.600 ;
        RECT 63.700 12.400 64.300 13.700 ;
        RECT 36.400 11.600 37.200 12.400 ;
        RECT 44.400 11.600 45.200 12.400 ;
        RECT 50.800 11.600 51.600 12.400 ;
        RECT 52.400 11.600 53.200 12.400 ;
        RECT 63.600 11.600 64.400 12.400 ;
        RECT 66.800 4.200 67.600 17.800 ;
        RECT 68.400 4.200 69.200 17.800 ;
        RECT 70.000 6.200 70.800 17.800 ;
        RECT 73.200 6.200 74.000 17.800 ;
        RECT 74.900 16.400 75.500 19.600 ;
        RECT 94.100 18.400 94.700 51.600 ;
        RECT 95.700 30.400 96.300 51.600 ;
        RECT 98.800 43.600 99.600 44.400 ;
        RECT 113.200 44.200 114.000 57.800 ;
        RECT 114.800 44.200 115.600 57.800 ;
        RECT 116.400 46.200 117.200 57.800 ;
        RECT 118.100 54.400 118.700 69.600 ;
        RECT 124.500 68.400 125.100 77.600 ;
        RECT 138.800 71.600 139.600 72.400 ;
        RECT 126.000 69.600 126.800 70.400 ;
        RECT 138.900 68.400 139.500 71.600 ;
        RECT 142.100 68.400 142.700 83.600 ;
        RECT 124.400 67.600 125.200 68.400 ;
        RECT 135.600 67.600 136.400 68.400 ;
        RECT 138.800 67.600 139.600 68.400 ;
        RECT 142.000 67.600 142.800 68.400 ;
        RECT 121.200 65.600 122.000 66.400 ;
        RECT 118.000 53.600 118.800 54.400 ;
        RECT 119.600 46.200 120.400 57.800 ;
        RECT 121.300 56.400 121.900 65.600 ;
        RECT 138.900 60.400 139.500 67.600 ;
        RECT 138.800 59.600 139.600 60.400 ;
        RECT 143.700 58.400 144.300 105.700 ;
        RECT 145.300 82.400 145.900 109.600 ;
        RECT 146.900 92.400 147.500 131.600 ;
        RECT 154.800 119.600 155.600 120.400 ;
        RECT 148.400 111.600 149.200 112.400 ;
        RECT 154.900 110.400 155.500 119.600 ;
        RECT 148.400 109.600 149.200 110.400 ;
        RECT 151.600 109.600 152.400 110.400 ;
        RECT 154.800 109.600 155.600 110.400 ;
        RECT 148.400 107.600 149.200 108.400 ;
        RECT 150.000 107.600 150.800 108.400 ;
        RECT 153.200 107.600 154.000 108.400 ;
        RECT 148.500 98.400 149.100 107.600 ;
        RECT 150.100 106.400 150.700 107.600 ;
        RECT 153.300 106.400 153.900 107.600 ;
        RECT 150.000 105.600 150.800 106.400 ;
        RECT 153.200 105.600 154.000 106.400 ;
        RECT 154.900 102.400 155.500 109.600 ;
        RECT 156.400 107.600 157.200 108.400 ;
        RECT 159.700 108.300 160.300 133.600 ;
        RECT 164.500 128.300 165.100 133.600 ;
        RECT 166.000 131.600 166.800 132.400 ;
        RECT 166.100 130.400 166.700 131.600 ;
        RECT 166.000 129.600 166.800 130.400 ;
        RECT 164.500 127.700 166.700 128.300 ;
        RECT 162.800 113.600 163.600 114.400 ;
        RECT 162.900 110.400 163.500 113.600 ;
        RECT 164.400 111.600 165.200 112.400 ;
        RECT 161.200 109.600 162.000 110.400 ;
        RECT 162.800 109.600 163.600 110.400 ;
        RECT 161.300 108.400 161.900 109.600 ;
        RECT 161.200 108.300 162.000 108.400 ;
        RECT 164.500 108.300 165.100 111.600 ;
        RECT 166.100 110.400 166.700 127.700 ;
        RECT 166.000 109.600 166.800 110.400 ;
        RECT 167.600 109.600 168.400 110.400 ;
        RECT 159.700 107.700 162.000 108.300 ;
        RECT 161.200 107.600 162.000 107.700 ;
        RECT 162.900 107.700 165.100 108.300 ;
        RECT 158.000 105.600 158.800 106.400 ;
        RECT 159.600 103.600 160.400 104.400 ;
        RECT 154.800 101.600 155.600 102.400 ;
        RECT 159.600 101.600 160.400 102.400 ;
        RECT 158.000 99.600 158.800 100.400 ;
        RECT 148.400 97.600 149.200 98.400 ;
        RECT 158.100 96.400 158.700 99.600 ;
        RECT 158.000 95.600 158.800 96.400 ;
        RECT 150.000 93.600 150.800 94.400 ;
        RECT 146.800 91.600 147.600 92.400 ;
        RECT 150.100 90.400 150.700 93.600 ;
        RECT 151.600 91.600 152.400 92.400 ;
        RECT 154.800 91.600 155.600 92.400 ;
        RECT 150.000 89.600 150.800 90.400 ;
        RECT 148.400 83.600 149.200 84.400 ;
        RECT 145.200 81.600 146.000 82.400 ;
        RECT 145.300 70.400 145.900 81.600 ;
        RECT 151.700 76.400 152.300 91.600 ;
        RECT 154.900 86.400 155.500 91.600 ;
        RECT 159.700 88.400 160.300 101.600 ;
        RECT 161.300 96.400 161.900 107.600 ;
        RECT 162.900 98.400 163.500 107.700 ;
        RECT 166.000 107.600 166.800 108.400 ;
        RECT 162.800 97.600 163.600 98.400 ;
        RECT 166.100 96.400 166.700 107.600 ;
        RECT 167.700 98.400 168.300 109.600 ;
        RECT 169.200 108.300 170.000 108.400 ;
        RECT 170.900 108.300 171.500 133.600 ;
        RECT 174.000 123.600 174.800 124.400 ;
        RECT 174.100 120.400 174.700 123.600 ;
        RECT 174.000 119.600 174.800 120.400 ;
        RECT 175.700 114.400 176.300 133.600 ;
        RECT 182.100 132.400 182.700 139.600 ;
        RECT 193.300 138.400 193.900 149.600 ;
        RECT 194.900 148.400 195.500 151.600 ;
        RECT 198.100 148.400 198.700 159.600 ;
        RECT 204.400 151.600 205.200 152.400 ;
        RECT 202.800 149.600 203.600 150.400 ;
        RECT 194.800 147.600 195.600 148.400 ;
        RECT 198.000 147.600 198.800 148.400 ;
        RECT 199.600 145.600 200.400 146.400 ;
        RECT 202.800 145.600 203.600 146.400 ;
        RECT 194.800 139.600 195.600 140.400 ;
        RECT 186.800 137.600 187.600 138.400 ;
        RECT 193.200 137.600 194.000 138.400 ;
        RECT 177.200 131.600 178.000 132.400 ;
        RECT 182.000 131.600 182.800 132.400 ;
        RECT 175.600 113.600 176.400 114.400 ;
        RECT 177.300 110.400 177.900 131.600 ;
        RECT 186.900 130.400 187.500 137.600 ;
        RECT 194.900 136.400 195.500 139.600 ;
        RECT 191.600 135.600 192.400 136.400 ;
        RECT 194.800 135.600 195.600 136.400 ;
        RECT 196.400 135.600 197.200 136.400 ;
        RECT 191.700 134.400 192.300 135.600 ;
        RECT 190.000 133.600 190.800 134.400 ;
        RECT 191.600 133.600 192.400 134.400 ;
        RECT 190.100 132.400 190.700 133.600 ;
        RECT 196.500 132.400 197.100 135.600 ;
        RECT 199.700 134.400 200.300 145.600 ;
        RECT 202.900 136.400 203.500 145.600 ;
        RECT 202.800 135.600 203.600 136.400 ;
        RECT 199.600 133.600 200.400 134.400 ;
        RECT 202.900 132.400 203.500 135.600 ;
        RECT 204.500 134.400 205.100 151.600 ;
        RECT 212.500 150.400 213.100 173.600 ;
        RECT 214.000 166.200 214.800 177.800 ;
        RECT 215.600 175.600 216.400 176.400 ;
        RECT 217.200 166.200 218.000 177.800 ;
        RECT 218.800 164.200 219.600 177.800 ;
        RECT 220.400 164.200 221.200 177.800 ;
        RECT 222.000 164.200 222.800 177.800 ;
        RECT 242.800 173.600 243.600 174.400 ;
        RECT 231.600 163.600 232.400 164.400 ;
        RECT 241.200 163.600 242.000 164.400 ;
        RECT 215.600 151.600 216.400 152.400 ;
        RECT 221.800 151.800 222.600 152.600 ;
        RECT 228.400 151.800 229.200 152.600 ;
        RECT 207.600 149.600 208.400 150.400 ;
        RECT 210.800 149.600 211.600 150.400 ;
        RECT 212.400 149.600 213.200 150.400 ;
        RECT 207.700 148.400 208.300 149.600 ;
        RECT 207.600 147.600 208.400 148.400 ;
        RECT 209.200 147.600 210.000 148.400 ;
        RECT 207.600 145.600 208.400 146.400 ;
        RECT 206.000 143.600 206.800 144.400 ;
        RECT 206.100 138.400 206.700 143.600 ;
        RECT 207.700 138.400 208.300 145.600 ;
        RECT 206.000 137.600 206.800 138.400 ;
        RECT 207.600 137.600 208.400 138.400 ;
        RECT 204.400 133.600 205.200 134.400 ;
        RECT 206.100 132.400 206.700 137.600 ;
        RECT 190.000 131.600 190.800 132.400 ;
        RECT 196.400 131.600 197.200 132.400 ;
        RECT 199.600 131.600 200.400 132.400 ;
        RECT 201.200 131.600 202.000 132.400 ;
        RECT 202.800 131.600 203.600 132.400 ;
        RECT 206.000 131.600 206.800 132.400 ;
        RECT 178.800 129.600 179.600 130.400 ;
        RECT 186.800 129.600 187.600 130.400 ;
        RECT 178.900 118.400 179.500 129.600 ;
        RECT 178.800 117.600 179.600 118.400 ;
        RECT 190.100 110.400 190.700 131.600 ;
        RECT 201.300 130.300 201.900 131.600 ;
        RECT 199.700 129.700 201.900 130.300 ;
        RECT 199.700 128.400 200.300 129.700 ;
        RECT 199.600 127.600 200.400 128.400 ;
        RECT 202.900 126.400 203.500 131.600 ;
        RECT 206.000 129.600 206.800 130.400 ;
        RECT 199.600 125.600 200.400 126.400 ;
        RECT 202.800 125.600 203.600 126.400 ;
        RECT 174.000 109.600 174.800 110.400 ;
        RECT 177.200 109.600 178.000 110.400 ;
        RECT 190.000 109.600 190.800 110.400 ;
        RECT 196.400 109.600 197.200 110.400 ;
        RECT 169.200 107.700 171.500 108.300 ;
        RECT 169.200 107.600 170.000 107.700 ;
        RECT 167.600 97.600 168.400 98.400 ;
        RECT 169.300 96.400 169.900 107.600 ;
        RECT 170.800 105.600 171.600 106.400 ;
        RECT 175.600 105.600 176.400 106.400 ;
        RECT 170.900 100.400 171.500 105.600 ;
        RECT 170.800 99.600 171.600 100.400 ;
        RECT 175.700 98.400 176.300 105.600 ;
        RECT 177.300 104.400 177.900 109.600 ;
        RECT 178.800 107.600 179.600 108.400 ;
        RECT 183.600 107.600 184.400 108.400 ;
        RECT 190.100 106.400 190.700 109.600 ;
        RECT 182.000 105.600 182.800 106.400 ;
        RECT 190.000 105.600 190.800 106.400 ;
        RECT 198.000 105.600 198.800 106.400 ;
        RECT 177.200 103.600 178.000 104.400 ;
        RECT 182.100 98.400 182.700 105.600 ;
        RECT 194.800 103.600 195.600 104.400 ;
        RECT 194.900 102.400 195.500 103.600 ;
        RECT 194.800 101.600 195.600 102.400 ;
        RECT 170.800 97.600 171.600 98.400 ;
        RECT 175.600 97.600 176.400 98.400 ;
        RECT 182.000 97.600 182.800 98.400 ;
        RECT 196.400 97.600 197.200 98.400 ;
        RECT 170.900 96.400 171.500 97.600 ;
        RECT 161.200 95.600 162.000 96.400 ;
        RECT 164.400 95.600 165.200 96.400 ;
        RECT 166.000 95.600 166.800 96.400 ;
        RECT 169.200 95.600 170.000 96.400 ;
        RECT 170.800 95.600 171.600 96.400 ;
        RECT 180.400 95.600 181.200 96.400 ;
        RECT 169.300 92.400 169.900 95.600 ;
        RECT 198.100 94.400 198.700 105.600 ;
        RECT 199.700 94.400 200.300 125.600 ;
        RECT 202.800 123.600 203.600 124.400 ;
        RECT 202.900 112.400 203.500 123.600 ;
        RECT 201.200 111.600 202.000 112.400 ;
        RECT 202.800 111.600 203.600 112.400 ;
        RECT 201.300 110.400 201.900 111.600 ;
        RECT 201.200 109.600 202.000 110.400 ;
        RECT 206.000 109.600 206.800 110.400 ;
        RECT 204.400 107.600 205.200 108.400 ;
        RECT 206.100 102.400 206.700 109.600 ;
        RECT 207.600 108.300 208.400 108.400 ;
        RECT 209.300 108.300 209.900 147.600 ;
        RECT 210.900 146.400 211.500 149.600 ;
        RECT 215.700 148.400 216.300 151.600 ;
        RECT 218.800 149.600 219.600 150.400 ;
        RECT 218.900 148.400 219.500 149.600 ;
        RECT 215.600 147.600 216.400 148.400 ;
        RECT 218.800 147.600 219.600 148.400 ;
        RECT 220.400 147.600 221.200 148.400 ;
        RECT 210.800 145.600 211.600 146.400 ;
        RECT 218.800 139.600 219.600 140.400 ;
        RECT 218.900 138.400 219.500 139.600 ;
        RECT 218.800 137.600 219.600 138.400 ;
        RECT 220.500 136.400 221.100 147.600 ;
        RECT 221.800 147.000 222.400 151.800 ;
        RECT 224.400 148.400 225.200 148.600 ;
        RECT 228.600 148.400 229.200 151.800 ;
        RECT 231.700 150.400 232.300 163.600 ;
        RECT 233.200 153.600 234.000 154.400 ;
        RECT 233.300 150.400 233.900 153.600 ;
        RECT 236.400 151.600 237.200 152.400 ;
        RECT 239.600 151.600 240.400 152.400 ;
        RECT 231.600 149.600 232.400 150.400 ;
        RECT 233.200 149.600 234.000 150.400 ;
        RECT 236.400 149.600 237.200 150.400 ;
        RECT 236.500 148.400 237.100 149.600 ;
        RECT 224.400 147.800 229.200 148.400 ;
        RECT 223.600 147.000 224.400 147.200 ;
        RECT 227.000 147.000 227.800 147.200 ;
        RECT 228.600 147.000 229.200 147.800 ;
        RECT 231.600 147.600 232.400 148.400 ;
        RECT 234.800 147.600 235.600 148.400 ;
        RECT 236.400 147.600 237.200 148.400 ;
        RECT 221.800 146.200 222.600 147.000 ;
        RECT 223.600 146.400 227.800 147.000 ;
        RECT 228.400 146.200 229.200 147.000 ;
        RECT 223.600 143.600 224.400 144.400 ;
        RECT 215.600 135.600 216.400 136.400 ;
        RECT 217.200 135.600 218.000 136.400 ;
        RECT 220.400 135.600 221.200 136.400 ;
        RECT 226.800 135.600 227.600 136.400 ;
        RECT 231.600 135.600 232.400 136.400 ;
        RECT 217.300 134.400 217.900 135.600 ;
        RECT 226.900 134.400 227.500 135.600 ;
        RECT 231.700 134.400 232.300 135.600 ;
        RECT 212.400 133.600 213.200 134.400 ;
        RECT 217.200 133.600 218.000 134.400 ;
        RECT 220.400 133.600 221.200 134.400 ;
        RECT 226.800 133.600 227.600 134.400 ;
        RECT 231.600 133.600 232.400 134.400 ;
        RECT 222.000 131.600 222.800 132.400 ;
        RECT 226.800 131.600 227.600 132.400 ;
        RECT 233.200 131.600 234.000 132.400 ;
        RECT 214.000 123.600 214.800 124.400 ;
        RECT 214.100 112.400 214.700 123.600 ;
        RECT 214.000 111.600 214.800 112.400 ;
        RECT 212.400 109.600 213.200 110.400 ;
        RECT 207.600 107.700 209.900 108.300 ;
        RECT 207.600 107.600 208.400 107.700 ;
        RECT 202.800 101.600 203.600 102.400 ;
        RECT 206.000 101.600 206.800 102.400 ;
        RECT 201.200 97.600 202.000 98.400 ;
        RECT 201.300 94.400 201.900 97.600 ;
        RECT 174.000 93.600 174.800 94.400 ;
        RECT 178.800 93.600 179.600 94.400 ;
        RECT 198.000 93.600 198.800 94.400 ;
        RECT 199.600 93.600 200.400 94.400 ;
        RECT 201.200 93.600 202.000 94.400 ;
        RECT 169.200 91.600 170.000 92.400 ;
        RECT 169.200 89.600 170.000 90.400 ;
        RECT 169.300 88.400 169.900 89.600 ;
        RECT 159.600 87.600 160.400 88.400 ;
        RECT 169.200 87.600 170.000 88.400 ;
        RECT 154.800 85.600 155.600 86.400 ;
        RECT 154.900 78.400 155.500 85.600 ;
        RECT 154.800 77.600 155.600 78.400 ;
        RECT 151.600 75.600 152.400 76.400 ;
        RECT 154.800 75.600 155.600 76.400 ;
        RECT 154.900 74.400 155.500 75.600 ;
        RECT 154.800 73.600 155.600 74.400 ;
        RECT 159.700 74.300 160.300 87.600 ;
        RECT 172.400 85.600 173.200 86.400 ;
        RECT 172.500 84.400 173.100 85.600 ;
        RECT 161.200 83.600 162.000 84.400 ;
        RECT 172.400 83.600 173.200 84.400 ;
        RECT 161.300 76.400 161.900 83.600 ;
        RECT 161.200 75.600 162.000 76.400 ;
        RECT 159.700 73.700 161.900 74.300 ;
        RECT 154.900 72.400 155.500 73.600 ;
        RECT 161.300 72.400 161.900 73.700 ;
        RECT 148.400 71.600 149.200 72.400 ;
        RECT 154.800 71.600 155.600 72.400 ;
        RECT 161.200 71.600 162.000 72.400 ;
        RECT 162.800 71.600 163.600 72.400 ;
        RECT 145.200 69.600 146.000 70.400 ;
        RECT 151.600 69.600 152.400 70.400 ;
        RECT 154.800 69.600 155.600 70.400 ;
        RECT 150.000 67.600 150.800 68.400 ;
        RECT 148.400 63.600 149.200 64.400 ;
        RECT 121.200 55.600 122.000 56.400 ;
        RECT 98.900 30.400 99.500 43.600 ;
        RECT 121.300 38.400 121.900 55.600 ;
        RECT 122.800 46.200 123.600 57.800 ;
        RECT 124.400 44.200 125.200 57.800 ;
        RECT 126.000 44.200 126.800 57.800 ;
        RECT 127.600 44.200 128.400 57.800 ;
        RECT 143.600 57.600 144.400 58.400 ;
        RECT 148.500 56.400 149.100 63.600 ;
        RECT 151.700 56.400 152.300 69.600 ;
        RECT 154.900 68.400 155.500 69.600 ;
        RECT 172.500 68.400 173.100 83.600 ;
        RECT 174.100 72.400 174.700 93.600 ;
        RECT 175.600 89.600 176.400 90.400 ;
        RECT 178.900 78.400 179.500 93.600 ;
        RECT 199.700 92.400 200.300 93.600 ;
        RECT 188.400 91.600 189.200 92.400 ;
        RECT 191.600 91.600 192.400 92.400 ;
        RECT 199.600 91.600 200.400 92.400 ;
        RECT 178.800 77.600 179.600 78.400 ;
        RECT 174.000 71.600 174.800 72.400 ;
        RECT 174.100 70.400 174.700 71.600 ;
        RECT 188.500 70.400 189.100 91.600 ;
        RECT 193.200 89.600 194.000 90.400 ;
        RECT 196.400 89.600 197.200 90.400 ;
        RECT 193.300 88.400 193.900 89.600 ;
        RECT 193.200 87.600 194.000 88.400 ;
        RECT 191.600 83.600 192.400 84.400 ;
        RECT 191.700 82.400 192.300 83.600 ;
        RECT 191.600 81.600 192.400 82.400 ;
        RECT 174.000 69.600 174.800 70.400 ;
        RECT 177.200 69.600 178.000 70.400 ;
        RECT 188.400 69.600 189.200 70.400 ;
        RECT 177.300 68.400 177.900 69.600 ;
        RECT 154.800 67.600 155.600 68.400 ;
        RECT 156.400 67.600 157.200 68.400 ;
        RECT 162.800 67.600 163.600 68.400 ;
        RECT 166.000 67.600 166.800 68.400 ;
        RECT 172.400 67.600 173.200 68.400 ;
        RECT 177.200 67.600 178.000 68.400 ;
        RECT 161.200 65.600 162.000 66.400 ;
        RECT 167.600 65.600 168.400 66.400 ;
        RECT 169.200 65.600 170.000 66.400 ;
        RECT 174.000 65.600 174.800 66.400 ;
        RECT 174.100 64.400 174.700 65.600 ;
        RECT 154.800 63.600 155.600 64.400 ;
        RECT 174.000 63.600 174.800 64.400 ;
        RECT 191.600 63.600 192.400 64.400 ;
        RECT 193.200 64.200 194.000 77.800 ;
        RECT 194.800 64.200 195.600 77.800 ;
        RECT 198.000 77.600 198.800 78.400 ;
        RECT 196.400 64.200 197.200 75.800 ;
        RECT 198.100 68.400 198.700 77.600 ;
        RECT 201.300 76.400 201.900 93.600 ;
        RECT 202.900 92.400 203.500 101.600 ;
        RECT 207.700 98.400 208.300 107.600 ;
        RECT 212.500 106.400 213.100 109.600 ;
        RECT 209.200 105.600 210.000 106.400 ;
        RECT 212.400 105.600 213.200 106.400 ;
        RECT 207.600 97.600 208.400 98.400 ;
        RECT 206.000 95.600 206.800 96.400 ;
        RECT 202.800 91.600 203.600 92.400 ;
        RECT 206.100 90.400 206.700 95.600 ;
        RECT 206.000 89.600 206.800 90.400 ;
        RECT 207.600 89.600 208.400 90.400 ;
        RECT 207.700 88.400 208.300 89.600 ;
        RECT 207.600 87.600 208.400 88.400 ;
        RECT 202.800 83.600 203.600 84.400 ;
        RECT 202.900 78.400 203.500 83.600 ;
        RECT 202.800 77.600 203.600 78.400 ;
        RECT 198.000 67.600 198.800 68.400 ;
        RECT 199.600 64.200 200.400 75.800 ;
        RECT 201.200 75.600 202.000 76.400 ;
        RECT 201.200 71.600 202.000 72.400 ;
        RECT 201.300 66.400 201.900 71.600 ;
        RECT 201.200 65.600 202.000 66.400 ;
        RECT 202.800 64.200 203.600 75.800 ;
        RECT 204.400 64.200 205.200 77.800 ;
        RECT 206.000 64.200 206.800 77.800 ;
        RECT 207.600 64.200 208.400 77.800 ;
        RECT 209.300 70.400 209.900 105.600 ;
        RECT 212.400 103.600 213.200 104.400 ;
        RECT 217.200 104.200 218.000 117.800 ;
        RECT 218.800 104.200 219.600 117.800 ;
        RECT 220.400 104.200 221.200 115.800 ;
        RECT 222.000 107.600 222.800 108.400 ;
        RECT 223.600 104.200 224.400 115.800 ;
        RECT 225.200 105.600 226.000 106.400 ;
        RECT 226.800 104.200 227.600 115.800 ;
        RECT 228.400 104.200 229.200 117.800 ;
        RECT 230.000 104.200 230.800 117.800 ;
        RECT 231.600 104.200 232.400 117.800 ;
        RECT 234.900 114.400 235.500 147.600 ;
        RECT 236.500 138.400 237.100 147.600 ;
        RECT 241.300 138.400 241.900 163.600 ;
        RECT 242.900 156.400 243.500 173.600 ;
        RECT 249.200 171.600 250.000 172.400 ;
        RECT 249.300 168.400 249.900 171.600 ;
        RECT 249.200 167.600 250.000 168.400 ;
        RECT 242.800 155.600 243.600 156.400 ;
        RECT 244.400 153.600 245.200 154.400 ;
        RECT 249.200 143.600 250.000 144.400 ;
        RECT 236.400 137.600 237.200 138.400 ;
        RECT 241.200 137.600 242.000 138.400 ;
        RECT 246.000 137.600 246.800 138.400 ;
        RECT 236.400 135.600 237.200 136.400 ;
        RECT 241.200 135.600 242.000 136.400 ;
        RECT 244.400 135.600 245.200 136.400 ;
        RECT 236.500 130.400 237.100 135.600 ;
        RECT 238.000 131.600 238.800 132.400 ;
        RECT 244.500 130.400 245.100 135.600 ;
        RECT 246.100 132.400 246.700 137.600 ;
        RECT 246.000 131.600 246.800 132.400 ;
        RECT 236.400 129.600 237.200 130.400 ;
        RECT 238.000 129.600 238.800 130.400 ;
        RECT 244.400 129.600 245.200 130.400 ;
        RECT 234.800 113.600 235.600 114.400 ;
        RECT 210.800 97.600 211.600 98.400 ;
        RECT 210.900 92.400 211.500 97.600 ;
        RECT 212.500 94.400 213.100 103.600 ;
        RECT 238.100 102.400 238.700 129.600 ;
        RECT 247.600 128.300 248.400 128.400 ;
        RECT 249.300 128.300 249.900 143.600 ;
        RECT 247.600 127.700 249.900 128.300 ;
        RECT 247.600 127.600 248.400 127.700 ;
        RECT 242.800 123.600 243.600 124.400 ;
        RECT 249.200 123.600 250.000 124.400 ;
        RECT 242.900 110.400 243.500 123.600 ;
        RECT 242.800 109.600 243.600 110.400 ;
        RECT 247.600 109.600 248.400 110.400 ;
        RECT 239.600 103.600 240.400 104.400 ;
        RECT 241.200 103.600 242.000 104.400 ;
        RECT 226.800 101.600 227.600 102.400 ;
        RECT 238.000 101.600 238.800 102.400 ;
        RECT 226.900 98.400 227.500 101.600 ;
        RECT 225.200 97.600 226.000 98.400 ;
        RECT 226.800 97.600 227.600 98.400 ;
        RECT 228.400 97.600 229.200 98.400 ;
        RECT 214.000 95.600 214.800 96.400 ;
        RECT 217.200 95.600 218.000 96.400 ;
        RECT 222.000 95.600 222.800 96.400 ;
        RECT 217.300 94.400 217.900 95.600 ;
        RECT 212.400 93.600 213.200 94.400 ;
        RECT 217.200 93.600 218.000 94.400 ;
        RECT 210.800 91.600 211.600 92.400 ;
        RECT 218.800 91.600 219.600 92.400 ;
        RECT 218.900 90.400 219.500 91.600 ;
        RECT 214.000 89.600 214.800 90.400 ;
        RECT 217.200 89.600 218.000 90.400 ;
        RECT 218.800 89.600 219.600 90.400 ;
        RECT 214.100 88.400 214.700 89.600 ;
        RECT 217.300 88.400 217.900 89.600 ;
        RECT 210.800 87.600 211.600 88.400 ;
        RECT 214.000 87.600 214.800 88.400 ;
        RECT 217.200 87.600 218.000 88.400 ;
        RECT 222.100 78.400 222.700 95.600 ;
        RECT 225.300 94.400 225.900 97.600 ;
        RECT 228.500 96.400 229.100 97.600 ;
        RECT 238.100 96.400 238.700 101.600 ;
        RECT 228.400 95.600 229.200 96.400 ;
        RECT 238.000 95.600 238.800 96.400 ;
        RECT 223.600 93.600 224.400 94.400 ;
        RECT 225.200 93.600 226.000 94.400 ;
        RECT 230.000 93.600 230.800 94.400 ;
        RECT 234.800 93.600 235.600 94.400 ;
        RECT 223.700 92.400 224.300 93.600 ;
        RECT 230.100 92.400 230.700 93.600 ;
        RECT 234.900 92.400 235.500 93.600 ;
        RECT 223.600 91.600 224.400 92.400 ;
        RECT 230.000 91.600 230.800 92.400 ;
        RECT 233.200 91.600 234.000 92.400 ;
        RECT 234.800 91.600 235.600 92.400 ;
        RECT 233.300 90.300 233.900 91.600 ;
        RECT 238.100 90.400 238.700 95.600 ;
        RECT 239.700 90.400 240.300 103.600 ;
        RECT 241.300 102.400 241.900 103.600 ;
        RECT 241.200 101.600 242.000 102.400 ;
        RECT 241.200 95.600 242.000 96.400 ;
        RECT 241.300 94.400 241.900 95.600 ;
        RECT 242.900 94.400 243.500 109.600 ;
        RECT 247.600 97.600 248.400 98.400 ;
        RECT 246.000 95.600 246.800 96.400 ;
        RECT 249.300 96.300 249.900 123.600 ;
        RECT 247.700 95.700 249.900 96.300 ;
        RECT 241.200 93.600 242.000 94.400 ;
        RECT 242.800 93.600 243.600 94.400 ;
        RECT 242.900 92.400 243.500 93.600 ;
        RECT 242.800 91.600 243.600 92.400 ;
        RECT 234.800 90.300 235.600 90.400 ;
        RECT 233.300 89.700 235.600 90.300 ;
        RECT 234.800 89.600 235.600 89.700 ;
        RECT 238.000 89.600 238.800 90.400 ;
        RECT 239.600 89.600 240.400 90.400 ;
        RECT 217.200 77.600 218.000 78.400 ;
        RECT 222.000 77.600 222.800 78.400 ;
        RECT 222.000 75.600 222.800 76.400 ;
        RECT 209.200 69.600 210.000 70.400 ;
        RECT 220.400 69.600 221.200 70.400 ;
        RECT 222.100 68.400 222.700 75.600 ;
        RECT 239.700 74.400 240.300 89.600 ;
        RECT 244.400 75.600 245.200 76.400 ;
        RECT 239.600 73.600 240.400 74.400 ;
        RECT 242.800 73.600 243.600 74.400 ;
        RECT 226.800 71.600 227.600 72.400 ;
        RECT 233.400 71.800 234.200 72.600 ;
        RECT 239.600 71.800 240.400 72.600 ;
        RECT 242.900 72.400 243.500 73.600 ;
        RECT 244.500 72.400 245.100 75.600 ;
        RECT 246.000 73.600 246.800 74.400 ;
        RECT 226.900 70.400 227.500 71.600 ;
        RECT 226.800 69.600 227.600 70.400 ;
        RECT 228.400 69.600 229.200 70.400 ;
        RECT 231.600 69.600 232.400 70.400 ;
        RECT 231.700 68.400 232.300 69.600 ;
        RECT 222.000 67.600 222.800 68.400 ;
        RECT 225.200 67.600 226.000 68.400 ;
        RECT 230.000 67.600 230.800 68.400 ;
        RECT 231.600 67.600 232.400 68.400 ;
        RECT 225.300 66.400 225.900 67.600 ;
        RECT 230.100 66.400 230.700 67.600 ;
        RECT 233.400 67.000 234.000 71.800 ;
        RECT 234.600 69.800 235.400 70.600 ;
        RECT 234.800 68.400 235.400 69.800 ;
        RECT 239.800 68.400 240.400 71.800 ;
        RECT 242.800 71.600 243.600 72.400 ;
        RECT 244.400 71.600 245.200 72.400 ;
        RECT 247.700 72.300 248.300 95.700 ;
        RECT 249.200 93.600 250.000 94.400 ;
        RECT 250.800 73.600 251.600 74.400 ;
        RECT 247.700 71.700 249.900 72.300 ;
        RECT 234.800 67.800 240.400 68.400 ;
        RECT 234.800 67.000 235.600 67.200 ;
        RECT 238.200 67.000 239.000 67.200 ;
        RECT 239.800 67.000 240.400 67.800 ;
        RECT 233.400 66.400 239.000 67.000 ;
        RECT 225.200 65.600 226.000 66.400 ;
        RECT 230.000 65.600 230.800 66.400 ;
        RECT 233.400 66.200 234.200 66.400 ;
        RECT 239.600 66.200 240.400 67.000 ;
        RECT 217.200 63.600 218.000 64.400 ;
        RECT 223.600 63.600 224.400 64.400 ;
        RECT 153.200 59.600 154.000 60.400 ;
        RECT 153.300 58.400 153.900 59.600 ;
        RECT 153.200 57.600 154.000 58.400 ;
        RECT 137.200 55.600 138.000 56.400 ;
        RECT 142.000 55.600 142.800 56.400 ;
        RECT 148.400 55.600 149.200 56.400 ;
        RECT 151.600 55.600 152.400 56.400 ;
        RECT 138.800 53.600 139.600 54.400 ;
        RECT 148.400 53.600 149.200 54.400 ;
        RECT 108.400 37.600 109.200 38.400 ;
        RECT 121.200 37.600 122.000 38.400 ;
        RECT 108.500 30.400 109.100 37.600 ;
        RECT 124.400 31.600 125.200 32.400 ;
        RECT 124.500 30.400 125.100 31.600 ;
        RECT 95.600 29.600 96.400 30.400 ;
        RECT 98.800 29.600 99.600 30.400 ;
        RECT 102.000 29.600 102.800 30.400 ;
        RECT 106.800 29.600 107.600 30.400 ;
        RECT 108.400 29.600 109.200 30.400 ;
        RECT 116.400 29.600 117.200 30.400 ;
        RECT 124.400 29.600 125.200 30.400 ;
        RECT 143.600 29.600 144.400 30.400 ;
        RECT 146.800 29.600 147.600 30.400 ;
        RECT 106.900 28.400 107.500 29.600 ;
        RECT 102.000 27.600 102.800 28.400 ;
        RECT 106.800 27.600 107.600 28.400 ;
        RECT 95.600 23.600 96.400 24.400 ;
        RECT 100.400 23.600 101.200 24.400 ;
        RECT 74.800 15.600 75.600 16.400 ;
        RECT 76.400 6.200 77.200 17.800 ;
        RECT 78.000 4.200 78.800 17.800 ;
        RECT 79.600 4.200 80.400 17.800 ;
        RECT 81.200 4.200 82.000 17.800 ;
        RECT 94.000 17.600 94.800 18.400 ;
        RECT 90.800 13.600 91.800 14.400 ;
        RECT 94.000 12.300 94.800 12.400 ;
        RECT 95.700 12.300 96.300 23.600 ;
        RECT 100.500 18.400 101.100 23.600 ;
        RECT 100.400 17.600 101.200 18.400 ;
        RECT 111.600 15.600 112.400 16.400 ;
        RECT 111.700 12.400 112.300 15.600 ;
        RECT 116.500 12.400 117.100 29.600 ;
        RECT 140.400 25.600 141.200 26.400 ;
        RECT 140.500 24.400 141.100 25.600 ;
        RECT 143.700 24.400 144.300 29.600 ;
        RECT 146.900 28.400 147.500 29.600 ;
        RECT 148.500 28.400 149.100 53.600 ;
        RECT 154.900 48.400 155.500 63.600 ;
        RECT 174.100 60.400 174.700 63.600 ;
        RECT 174.000 59.600 174.800 60.400 ;
        RECT 161.200 55.600 162.000 56.400 ;
        RECT 154.800 47.600 155.600 48.400 ;
        RECT 151.600 29.600 152.400 30.400 ;
        RECT 146.800 27.600 147.600 28.400 ;
        RECT 148.400 27.600 149.200 28.400 ;
        RECT 124.400 23.600 125.200 24.400 ;
        RECT 140.400 23.600 141.200 24.400 ;
        RECT 143.600 23.600 144.400 24.400 ;
        RECT 121.200 15.600 122.000 16.400 ;
        RECT 94.000 11.700 96.300 12.300 ;
        RECT 94.000 11.600 94.800 11.700 ;
        RECT 111.600 11.600 112.400 12.400 ;
        RECT 116.400 11.600 117.200 12.400 ;
        RECT 122.600 11.600 123.600 12.400 ;
        RECT 124.500 10.400 125.100 23.600 ;
        RECT 140.500 20.300 141.100 23.600 ;
        RECT 138.900 19.700 141.100 20.300 ;
        RECT 119.600 9.600 120.400 10.400 ;
        RECT 124.400 9.600 125.200 10.400 ;
        RECT 132.400 4.200 133.200 17.800 ;
        RECT 134.000 4.200 134.800 17.800 ;
        RECT 135.600 4.200 136.400 17.800 ;
        RECT 137.200 6.200 138.000 17.800 ;
        RECT 138.900 16.400 139.500 19.700 ;
        RECT 138.800 15.600 139.600 16.400 ;
        RECT 140.400 6.200 141.200 17.800 ;
        RECT 142.000 15.600 142.800 16.400 ;
        RECT 142.100 14.400 142.700 15.600 ;
        RECT 142.000 13.600 142.800 14.400 ;
        RECT 143.600 6.200 144.400 17.800 ;
        RECT 145.200 4.200 146.000 17.800 ;
        RECT 146.800 4.200 147.600 17.800 ;
        RECT 151.700 12.400 152.300 29.600 ;
        RECT 156.400 24.200 157.200 37.800 ;
        RECT 158.000 24.200 158.800 37.800 ;
        RECT 159.600 24.200 160.400 35.800 ;
        RECT 161.300 28.400 161.900 55.600 ;
        RECT 162.800 44.200 163.600 57.800 ;
        RECT 164.400 44.200 165.200 57.800 ;
        RECT 166.000 44.200 166.800 57.800 ;
        RECT 167.600 46.200 168.400 57.800 ;
        RECT 169.200 55.600 170.000 56.400 ;
        RECT 169.300 42.400 169.900 55.600 ;
        RECT 170.800 46.200 171.600 57.800 ;
        RECT 172.400 53.600 173.200 54.400 ;
        RECT 172.400 51.600 173.200 52.400 ;
        RECT 164.400 41.600 165.200 42.400 ;
        RECT 169.200 41.600 170.000 42.400 ;
        RECT 161.200 27.600 162.000 28.400 ;
        RECT 162.800 24.200 163.600 35.800 ;
        RECT 164.500 26.400 165.100 41.600 ;
        RECT 164.400 25.600 165.200 26.400 ;
        RECT 166.000 24.200 166.800 35.800 ;
        RECT 167.600 24.200 168.400 37.800 ;
        RECT 169.200 24.200 170.000 37.800 ;
        RECT 170.800 24.200 171.600 37.800 ;
        RECT 172.500 32.400 173.100 51.600 ;
        RECT 174.000 46.200 174.800 57.800 ;
        RECT 175.600 44.200 176.400 57.800 ;
        RECT 177.200 44.200 178.000 57.800 ;
        RECT 191.700 54.300 192.300 63.600 ;
        RECT 204.400 59.600 205.200 60.400 ;
        RECT 223.700 60.300 224.300 63.600 ;
        RECT 230.100 62.400 230.700 65.600 ;
        RECT 234.800 63.600 235.600 64.400 ;
        RECT 230.000 61.600 230.800 62.400 ;
        RECT 222.100 59.700 224.300 60.300 ;
        RECT 204.500 54.400 205.100 59.600 ;
        RECT 193.200 54.300 194.000 54.400 ;
        RECT 191.700 53.700 194.000 54.300 ;
        RECT 193.200 53.600 194.000 53.700 ;
        RECT 196.400 53.600 197.200 54.400 ;
        RECT 204.400 53.600 205.200 54.400 ;
        RECT 172.400 31.600 173.200 32.400 ;
        RECT 172.500 30.400 173.100 31.600 ;
        RECT 193.300 30.400 193.900 53.600 ;
        RECT 196.400 51.600 197.200 52.400 ;
        RECT 201.200 51.600 202.000 52.400 ;
        RECT 214.000 51.600 214.800 52.400 ;
        RECT 196.400 49.600 197.200 50.400 ;
        RECT 207.600 49.600 208.400 50.400 ;
        RECT 199.600 47.600 200.400 48.400 ;
        RECT 210.800 31.600 211.600 32.400 ;
        RECT 214.100 32.000 214.700 51.600 ;
        RECT 217.200 44.200 218.000 57.800 ;
        RECT 218.800 44.200 219.600 57.800 ;
        RECT 220.400 46.200 221.200 57.800 ;
        RECT 222.100 54.400 222.700 59.700 ;
        RECT 222.000 53.600 222.800 54.400 ;
        RECT 223.600 46.200 224.400 57.800 ;
        RECT 225.200 55.600 226.000 56.400 ;
        RECT 225.300 44.300 225.900 55.600 ;
        RECT 226.800 46.200 227.600 57.800 ;
        RECT 223.700 43.700 225.900 44.300 ;
        RECT 228.400 44.200 229.200 57.800 ;
        RECT 230.000 44.200 230.800 57.800 ;
        RECT 231.600 44.200 232.400 57.800 ;
        RECT 234.900 50.400 235.500 63.600 ;
        RECT 241.200 61.600 242.000 62.400 ;
        RECT 239.600 59.600 240.400 60.400 ;
        RECT 234.800 49.600 235.600 50.400 ;
        RECT 214.000 31.200 214.800 32.000 ;
        RECT 172.400 29.600 173.200 30.400 ;
        RECT 193.200 29.600 194.000 30.400 ;
        RECT 202.800 29.600 203.600 30.400 ;
        RECT 180.400 27.600 181.400 28.400 ;
        RECT 194.800 27.600 195.600 28.400 ;
        RECT 194.900 26.400 195.500 27.600 ;
        RECT 172.400 25.600 173.200 26.400 ;
        RECT 194.800 25.600 195.600 26.400 ;
        RECT 151.600 11.600 152.400 12.400 ;
        RECT 159.600 11.600 160.400 12.400 ;
        RECT 164.400 4.200 165.200 17.800 ;
        RECT 166.000 4.200 166.800 17.800 ;
        RECT 167.600 6.200 168.400 17.800 ;
        RECT 169.200 13.600 170.000 14.400 ;
        RECT 170.800 6.200 171.600 17.800 ;
        RECT 172.500 16.400 173.100 25.600 ;
        RECT 198.000 23.600 198.800 24.400 ;
        RECT 172.400 15.600 173.200 16.400 ;
        RECT 174.000 6.200 174.800 17.800 ;
        RECT 175.600 4.200 176.400 17.800 ;
        RECT 177.200 4.200 178.000 17.800 ;
        RECT 178.800 4.200 179.600 17.800 ;
        RECT 188.400 15.600 189.200 16.400 ;
        RECT 190.000 15.600 190.800 16.400 ;
        RECT 190.100 14.400 190.700 15.600 ;
        RECT 198.100 14.400 198.700 23.600 ;
        RECT 202.900 18.400 203.500 29.600 ;
        RECT 210.800 27.600 211.600 28.400 ;
        RECT 206.000 25.600 206.800 26.400 ;
        RECT 202.800 17.600 203.600 18.400 ;
        RECT 201.200 15.600 202.000 16.400 ;
        RECT 190.000 13.600 190.800 14.400 ;
        RECT 198.000 13.600 198.800 14.400 ;
        RECT 201.200 11.600 202.000 12.400 ;
        RECT 204.400 11.600 205.200 12.400 ;
        RECT 206.100 12.300 206.700 25.600 ;
        RECT 210.900 18.400 211.500 27.600 ;
        RECT 215.600 24.200 216.400 37.800 ;
        RECT 217.200 24.200 218.000 37.800 ;
        RECT 218.800 24.200 219.600 35.800 ;
        RECT 220.400 27.600 221.200 28.400 ;
        RECT 222.000 24.200 222.800 35.800 ;
        RECT 223.700 26.400 224.300 43.700 ;
        RECT 239.700 38.400 240.300 59.600 ;
        RECT 241.300 58.400 241.900 61.600 ;
        RECT 242.900 60.400 243.500 71.600 ;
        RECT 247.700 70.400 248.300 71.700 ;
        RECT 249.300 70.400 249.900 71.700 ;
        RECT 244.400 69.600 245.200 70.400 ;
        RECT 247.600 69.600 248.400 70.400 ;
        RECT 249.200 69.600 250.000 70.400 ;
        RECT 242.800 59.600 243.600 60.400 ;
        RECT 241.200 57.600 242.000 58.400 ;
        RECT 242.800 53.600 243.600 54.400 ;
        RECT 242.900 38.400 243.500 53.600 ;
        RECT 244.500 52.400 245.100 69.600 ;
        RECT 249.200 65.600 250.000 66.400 ;
        RECT 246.000 63.600 246.800 64.400 ;
        RECT 244.400 51.600 245.200 52.400 ;
        RECT 223.600 25.600 224.400 26.400 ;
        RECT 223.700 20.400 224.300 25.600 ;
        RECT 225.200 24.200 226.000 35.800 ;
        RECT 226.800 24.200 227.600 37.800 ;
        RECT 228.400 24.200 229.200 37.800 ;
        RECT 230.000 24.200 230.800 37.800 ;
        RECT 239.600 37.600 240.400 38.400 ;
        RECT 242.800 37.600 243.600 38.400 ;
        RECT 246.100 30.400 246.700 63.600 ;
        RECT 249.300 50.400 249.900 65.600 ;
        RECT 250.900 58.400 251.500 73.600 ;
        RECT 250.800 57.600 251.600 58.400 ;
        RECT 252.400 53.600 253.200 54.400 ;
        RECT 252.400 51.600 253.200 52.400 ;
        RECT 249.200 49.600 250.000 50.400 ;
        RECT 246.000 29.600 246.800 30.400 ;
        RECT 223.600 19.600 224.400 20.400 ;
        RECT 228.400 19.600 229.200 20.400 ;
        RECT 210.800 17.600 211.600 18.400 ;
        RECT 207.600 12.300 208.400 12.400 ;
        RECT 206.100 11.700 208.400 12.300 ;
        RECT 207.600 11.600 208.400 11.700 ;
        RECT 215.600 11.600 216.400 12.400 ;
        RECT 207.700 10.400 208.300 11.600 ;
        RECT 207.600 9.600 208.400 10.400 ;
        RECT 220.400 4.200 221.200 17.800 ;
        RECT 222.000 4.200 222.800 17.800 ;
        RECT 223.600 6.200 224.400 17.800 ;
        RECT 225.200 13.600 226.000 14.400 ;
        RECT 226.800 6.200 227.600 17.800 ;
        RECT 228.500 16.400 229.100 19.600 ;
        RECT 252.500 18.400 253.100 51.600 ;
        RECT 228.400 15.600 229.200 16.400 ;
        RECT 230.000 6.200 230.800 17.800 ;
        RECT 231.600 4.200 232.400 17.800 ;
        RECT 233.200 4.200 234.000 17.800 ;
        RECT 234.800 4.200 235.600 17.800 ;
        RECT 252.400 17.600 253.200 18.400 ;
        RECT 249.200 11.600 250.000 12.400 ;
        RECT 244.400 9.600 245.200 10.400 ;
      LAYER via2 ;
        RECT 7.600 147.600 8.400 148.400 ;
        RECT 7.600 13.600 8.400 14.400 ;
        RECT 90.800 13.600 91.600 14.400 ;
        RECT 122.800 11.600 123.600 12.400 ;
        RECT 180.400 27.600 181.200 28.400 ;
      LAYER metal3 ;
        RECT 26.800 178.300 27.600 178.400 ;
        RECT 47.600 178.300 48.400 178.400 ;
        RECT 26.800 177.700 48.400 178.300 ;
        RECT 26.800 177.600 27.600 177.700 ;
        RECT 47.600 177.600 48.400 177.700 ;
        RECT 7.600 176.300 8.400 176.400 ;
        RECT 41.200 176.300 42.000 176.400 ;
        RECT 7.600 175.700 42.000 176.300 ;
        RECT 7.600 175.600 8.400 175.700 ;
        RECT 41.200 175.600 42.000 175.700 ;
        RECT 79.600 176.300 80.400 176.400 ;
        RECT 126.000 176.300 126.800 176.400 ;
        RECT 158.000 176.300 158.800 176.400 ;
        RECT 169.200 176.300 170.000 176.400 ;
        RECT 215.600 176.300 216.400 176.400 ;
        RECT 218.800 176.300 219.600 176.400 ;
        RECT 79.600 175.700 219.600 176.300 ;
        RECT 79.600 175.600 80.400 175.700 ;
        RECT 126.000 175.600 126.800 175.700 ;
        RECT 158.000 175.600 158.800 175.700 ;
        RECT 169.200 175.600 170.000 175.700 ;
        RECT 215.600 175.600 216.400 175.700 ;
        RECT 218.800 175.600 219.600 175.700 ;
        RECT 44.400 174.300 45.200 174.400 ;
        RECT 49.200 174.300 50.000 174.400 ;
        RECT 44.400 173.700 50.000 174.300 ;
        RECT 44.400 173.600 45.200 173.700 ;
        RECT 49.200 173.600 50.000 173.700 ;
        RECT 76.400 174.300 77.200 174.400 ;
        RECT 90.800 174.300 91.600 174.400 ;
        RECT 76.400 173.700 91.600 174.300 ;
        RECT 76.400 173.600 77.200 173.700 ;
        RECT 90.800 173.600 91.600 173.700 ;
        RECT 166.000 174.300 166.800 174.400 ;
        RECT 183.600 174.300 184.400 174.400 ;
        RECT 166.000 173.700 184.400 174.300 ;
        RECT 166.000 173.600 166.800 173.700 ;
        RECT 183.600 173.600 184.400 173.700 ;
        RECT 34.800 172.300 35.600 172.400 ;
        RECT 66.800 172.300 67.600 172.400 ;
        RECT 34.800 171.700 67.600 172.300 ;
        RECT 34.800 171.600 35.600 171.700 ;
        RECT 66.800 171.600 67.600 171.700 ;
        RECT 166.000 172.300 166.800 172.400 ;
        RECT 202.800 172.300 203.600 172.400 ;
        RECT 166.000 171.700 203.600 172.300 ;
        RECT 166.000 171.600 166.800 171.700 ;
        RECT 202.800 171.600 203.600 171.700 ;
        RECT 148.400 169.600 149.200 170.400 ;
        RECT 234.800 168.300 235.600 168.400 ;
        RECT 249.200 168.300 250.000 168.400 ;
        RECT 234.800 167.700 250.000 168.300 ;
        RECT 234.800 167.600 235.600 167.700 ;
        RECT 249.200 167.600 250.000 167.700 ;
        RECT 110.000 164.300 110.800 164.400 ;
        RECT 118.000 164.300 118.800 164.400 ;
        RECT 110.000 163.700 118.800 164.300 ;
        RECT 110.000 163.600 110.800 163.700 ;
        RECT 118.000 163.600 118.800 163.700 ;
        RECT 130.800 164.300 131.600 164.400 ;
        RECT 143.600 164.300 144.400 164.400 ;
        RECT 130.800 163.700 144.400 164.300 ;
        RECT 130.800 163.600 131.600 163.700 ;
        RECT 143.600 163.600 144.400 163.700 ;
        RECT 122.800 162.300 123.600 162.400 ;
        RECT 129.200 162.300 130.000 162.400 ;
        RECT 122.800 161.700 130.000 162.300 ;
        RECT 122.800 161.600 123.600 161.700 ;
        RECT 129.200 161.600 130.000 161.700 ;
        RECT 194.800 160.300 195.600 160.400 ;
        RECT 198.000 160.300 198.800 160.400 ;
        RECT 194.800 159.700 198.800 160.300 ;
        RECT 194.800 159.600 195.600 159.700 ;
        RECT 198.000 159.600 198.800 159.700 ;
        RECT 55.600 158.300 56.400 158.400 ;
        RECT 68.400 158.300 69.200 158.400 ;
        RECT 55.600 157.700 69.200 158.300 ;
        RECT 55.600 157.600 56.400 157.700 ;
        RECT 68.400 157.600 69.200 157.700 ;
        RECT 138.800 156.300 139.600 156.400 ;
        RECT 146.800 156.300 147.600 156.400 ;
        RECT 138.800 155.700 147.600 156.300 ;
        RECT 138.800 155.600 139.600 155.700 ;
        RECT 146.800 155.600 147.600 155.700 ;
        RECT 238.000 156.300 238.800 156.400 ;
        RECT 242.800 156.300 243.600 156.400 ;
        RECT 238.000 155.700 243.600 156.300 ;
        RECT 238.000 155.600 238.800 155.700 ;
        RECT 242.800 155.600 243.600 155.700 ;
        RECT 233.200 154.300 234.000 154.400 ;
        RECT 244.400 154.300 245.200 154.400 ;
        RECT 233.200 153.700 245.200 154.300 ;
        RECT 233.200 153.600 234.000 153.700 ;
        RECT 244.400 153.600 245.200 153.700 ;
        RECT 236.400 152.300 237.200 152.400 ;
        RECT 239.600 152.300 240.400 152.400 ;
        RECT 236.400 151.700 240.400 152.300 ;
        RECT 236.400 151.600 237.200 151.700 ;
        RECT 239.600 151.600 240.400 151.700 ;
        RECT 34.800 150.300 35.600 150.400 ;
        RECT 47.600 150.300 48.400 150.400 ;
        RECT 34.800 149.700 48.400 150.300 ;
        RECT 34.800 149.600 35.600 149.700 ;
        RECT 47.600 149.600 48.400 149.700 ;
        RECT 50.800 150.300 51.600 150.400 ;
        RECT 70.000 150.300 70.800 150.400 ;
        RECT 50.800 149.700 70.800 150.300 ;
        RECT 50.800 149.600 51.600 149.700 ;
        RECT 70.000 149.600 70.800 149.700 ;
        RECT 87.600 150.300 88.400 150.400 ;
        RECT 103.600 150.300 104.400 150.400 ;
        RECT 87.600 149.700 104.400 150.300 ;
        RECT 87.600 149.600 88.400 149.700 ;
        RECT 103.600 149.600 104.400 149.700 ;
        RECT 119.600 150.300 120.400 150.400 ;
        RECT 132.400 150.300 133.200 150.400 ;
        RECT 137.200 150.300 138.000 150.400 ;
        RECT 119.600 149.700 138.000 150.300 ;
        RECT 119.600 149.600 120.400 149.700 ;
        RECT 132.400 149.600 133.200 149.700 ;
        RECT 137.200 149.600 138.000 149.700 ;
        RECT 174.000 150.300 174.800 150.400 ;
        RECT 180.400 150.300 181.200 150.400 ;
        RECT 174.000 149.700 181.200 150.300 ;
        RECT 174.000 149.600 174.800 149.700 ;
        RECT 180.400 149.600 181.200 149.700 ;
        RECT 183.600 150.300 184.400 150.400 ;
        RECT 193.200 150.300 194.000 150.400 ;
        RECT 183.600 149.700 194.000 150.300 ;
        RECT 183.600 149.600 184.400 149.700 ;
        RECT 193.200 149.600 194.000 149.700 ;
        RECT 202.800 150.300 203.600 150.400 ;
        RECT 207.600 150.300 208.400 150.400 ;
        RECT 218.800 150.300 219.600 150.400 ;
        RECT 231.600 150.300 232.400 150.400 ;
        RECT 202.800 149.700 232.400 150.300 ;
        RECT 202.800 149.600 203.600 149.700 ;
        RECT 207.600 149.600 208.400 149.700 ;
        RECT 218.800 149.600 219.600 149.700 ;
        RECT 231.600 149.600 232.400 149.700 ;
        RECT 7.600 148.300 8.400 148.400 ;
        RECT 41.200 148.300 42.000 148.400 ;
        RECT 7.600 147.700 42.000 148.300 ;
        RECT 7.600 147.600 8.400 147.700 ;
        RECT 41.200 147.600 42.000 147.700 ;
        RECT 92.400 148.300 93.200 148.400 ;
        RECT 95.600 148.300 96.400 148.400 ;
        RECT 92.400 147.700 96.400 148.300 ;
        RECT 92.400 147.600 93.200 147.700 ;
        RECT 95.600 147.600 96.400 147.700 ;
        RECT 98.800 148.300 99.600 148.400 ;
        RECT 106.800 148.300 107.600 148.400 ;
        RECT 121.200 148.300 122.000 148.400 ;
        RECT 126.000 148.300 126.800 148.400 ;
        RECT 98.800 147.700 126.800 148.300 ;
        RECT 98.800 147.600 99.600 147.700 ;
        RECT 106.800 147.600 107.600 147.700 ;
        RECT 121.200 147.600 122.000 147.700 ;
        RECT 126.000 147.600 126.800 147.700 ;
        RECT 180.400 148.300 181.200 148.400 ;
        RECT 194.800 148.300 195.600 148.400 ;
        RECT 209.200 148.300 210.000 148.400 ;
        RECT 215.600 148.300 216.400 148.400 ;
        RECT 180.400 147.700 195.600 148.300 ;
        RECT 180.400 147.600 181.200 147.700 ;
        RECT 194.800 147.600 195.600 147.700 ;
        RECT 199.700 147.700 216.400 148.300 ;
        RECT 199.700 146.400 200.300 147.700 ;
        RECT 209.200 147.600 210.000 147.700 ;
        RECT 215.600 147.600 216.400 147.700 ;
        RECT 220.400 148.300 221.200 148.400 ;
        RECT 231.600 148.300 232.400 148.400 ;
        RECT 236.400 148.300 237.200 148.400 ;
        RECT 220.400 147.700 237.200 148.300 ;
        RECT 220.400 147.600 221.200 147.700 ;
        RECT 231.600 147.600 232.400 147.700 ;
        RECT 236.400 147.600 237.200 147.700 ;
        RECT 23.600 146.300 24.400 146.400 ;
        RECT 60.400 146.300 61.200 146.400 ;
        RECT 23.600 145.700 61.200 146.300 ;
        RECT 23.600 145.600 24.400 145.700 ;
        RECT 60.400 145.600 61.200 145.700 ;
        RECT 102.000 146.300 102.800 146.400 ;
        RECT 108.400 146.300 109.200 146.400 ;
        RECT 102.000 145.700 109.200 146.300 ;
        RECT 102.000 145.600 102.800 145.700 ;
        RECT 108.400 145.600 109.200 145.700 ;
        RECT 175.600 146.300 176.400 146.400 ;
        RECT 182.000 146.300 182.800 146.400 ;
        RECT 199.600 146.300 200.400 146.400 ;
        RECT 175.600 145.700 200.400 146.300 ;
        RECT 175.600 145.600 176.400 145.700 ;
        RECT 182.000 145.600 182.800 145.700 ;
        RECT 199.600 145.600 200.400 145.700 ;
        RECT 207.600 146.300 208.400 146.400 ;
        RECT 210.800 146.300 211.600 146.400 ;
        RECT 207.600 145.700 211.600 146.300 ;
        RECT 207.600 145.600 208.400 145.700 ;
        RECT 210.800 145.600 211.600 145.700 ;
        RECT 50.800 144.300 51.600 144.400 ;
        RECT 97.200 144.300 98.000 144.400 ;
        RECT 50.800 143.700 98.000 144.300 ;
        RECT 50.800 143.600 51.600 143.700 ;
        RECT 97.200 143.600 98.000 143.700 ;
        RECT 170.800 144.300 171.600 144.400 ;
        RECT 174.000 144.300 174.800 144.400 ;
        RECT 170.800 143.700 174.800 144.300 ;
        RECT 170.800 143.600 171.600 143.700 ;
        RECT 174.000 143.600 174.800 143.700 ;
        RECT 177.200 144.300 178.000 144.400 ;
        RECT 223.600 144.300 224.400 144.400 ;
        RECT 177.200 143.700 224.400 144.300 ;
        RECT 177.200 143.600 178.000 143.700 ;
        RECT 223.600 143.600 224.400 143.700 ;
        RECT 26.800 142.300 27.600 142.400 ;
        RECT 55.600 142.300 56.400 142.400 ;
        RECT 26.800 141.700 56.400 142.300 ;
        RECT 26.800 141.600 27.600 141.700 ;
        RECT 55.600 141.600 56.400 141.700 ;
        RECT 57.200 142.300 58.000 142.400 ;
        RECT 74.800 142.300 75.600 142.400 ;
        RECT 57.200 141.700 75.600 142.300 ;
        RECT 57.200 141.600 58.000 141.700 ;
        RECT 74.800 141.600 75.600 141.700 ;
        RECT 154.800 142.300 155.600 142.400 ;
        RECT 161.200 142.300 162.000 142.400 ;
        RECT 154.800 141.700 162.000 142.300 ;
        RECT 154.800 141.600 155.600 141.700 ;
        RECT 161.200 141.600 162.000 141.700 ;
        RECT 95.600 140.300 96.400 140.400 ;
        RECT 100.400 140.300 101.200 140.400 ;
        RECT 95.600 139.700 101.200 140.300 ;
        RECT 95.600 139.600 96.400 139.700 ;
        RECT 100.400 139.600 101.200 139.700 ;
        RECT 130.800 140.300 131.600 140.400 ;
        RECT 132.400 140.300 133.200 140.400 ;
        RECT 130.800 139.700 133.200 140.300 ;
        RECT 130.800 139.600 131.600 139.700 ;
        RECT 132.400 139.600 133.200 139.700 ;
        RECT 140.400 140.300 141.200 140.400 ;
        RECT 154.800 140.300 155.600 140.400 ;
        RECT 182.000 140.300 182.800 140.400 ;
        RECT 140.400 139.700 182.800 140.300 ;
        RECT 140.400 139.600 141.200 139.700 ;
        RECT 154.800 139.600 155.600 139.700 ;
        RECT 182.000 139.600 182.800 139.700 ;
        RECT 194.800 140.300 195.600 140.400 ;
        RECT 218.800 140.300 219.600 140.400 ;
        RECT 194.800 139.700 219.600 140.300 ;
        RECT 194.800 139.600 195.600 139.700 ;
        RECT 218.800 139.600 219.600 139.700 ;
        RECT 68.400 138.300 69.200 138.400 ;
        RECT 76.400 138.300 77.200 138.400 ;
        RECT 84.400 138.300 85.200 138.400 ;
        RECT 68.400 137.700 85.200 138.300 ;
        RECT 68.400 137.600 69.200 137.700 ;
        RECT 76.400 137.600 77.200 137.700 ;
        RECT 84.400 137.600 85.200 137.700 ;
        RECT 111.600 138.300 112.400 138.400 ;
        RECT 114.800 138.300 115.600 138.400 ;
        RECT 111.600 137.700 115.600 138.300 ;
        RECT 111.600 137.600 112.400 137.700 ;
        RECT 114.800 137.600 115.600 137.700 ;
        RECT 158.000 138.300 158.800 138.400 ;
        RECT 177.200 138.300 178.000 138.400 ;
        RECT 158.000 137.700 178.000 138.300 ;
        RECT 158.000 137.600 158.800 137.700 ;
        RECT 177.200 137.600 178.000 137.700 ;
        RECT 186.800 138.300 187.600 138.400 ;
        RECT 206.000 138.300 206.800 138.400 ;
        RECT 241.200 138.300 242.000 138.400 ;
        RECT 246.000 138.300 246.800 138.400 ;
        RECT 186.800 137.700 206.800 138.300 ;
        RECT 186.800 137.600 187.600 137.700 ;
        RECT 206.000 137.600 206.800 137.700 ;
        RECT 236.500 137.700 246.800 138.300 ;
        RECT 236.500 136.400 237.100 137.700 ;
        RECT 241.200 137.600 242.000 137.700 ;
        RECT 246.000 137.600 246.800 137.700 ;
        RECT 7.600 136.300 8.400 136.400 ;
        RECT 41.200 136.300 42.000 136.400 ;
        RECT 7.600 135.700 42.000 136.300 ;
        RECT 7.600 135.600 8.400 135.700 ;
        RECT 41.200 135.600 42.000 135.700 ;
        RECT 42.800 136.300 43.600 136.400 ;
        RECT 50.800 136.300 51.600 136.400 ;
        RECT 42.800 135.700 51.600 136.300 ;
        RECT 42.800 135.600 43.600 135.700 ;
        RECT 50.800 135.600 51.600 135.700 ;
        RECT 111.600 136.300 112.400 136.400 ;
        RECT 135.600 136.300 136.400 136.400 ;
        RECT 138.800 136.300 139.600 136.400 ;
        RECT 111.600 135.700 136.400 136.300 ;
        RECT 111.600 135.600 112.400 135.700 ;
        RECT 135.600 135.600 136.400 135.700 ;
        RECT 137.300 135.700 139.600 136.300 ;
        RECT 26.800 134.300 27.600 134.400 ;
        RECT 47.600 134.300 48.400 134.400 ;
        RECT 26.800 133.700 48.400 134.300 ;
        RECT 26.800 133.600 27.600 133.700 ;
        RECT 47.600 133.600 48.400 133.700 ;
        RECT 78.000 134.300 78.800 134.400 ;
        RECT 79.600 134.300 80.400 134.400 ;
        RECT 78.000 133.700 80.400 134.300 ;
        RECT 78.000 133.600 78.800 133.700 ;
        RECT 79.600 133.600 80.400 133.700 ;
        RECT 135.600 134.300 136.400 134.400 ;
        RECT 137.300 134.300 137.900 135.700 ;
        RECT 138.800 135.600 139.600 135.700 ;
        RECT 162.800 136.300 163.600 136.400 ;
        RECT 166.000 136.300 166.800 136.400 ;
        RECT 162.800 135.700 166.800 136.300 ;
        RECT 162.800 135.600 163.600 135.700 ;
        RECT 166.000 135.600 166.800 135.700 ;
        RECT 191.600 136.300 192.400 136.400 ;
        RECT 202.800 136.300 203.600 136.400 ;
        RECT 191.600 135.700 203.600 136.300 ;
        RECT 191.600 135.600 192.400 135.700 ;
        RECT 202.800 135.600 203.600 135.700 ;
        RECT 215.600 136.300 216.400 136.400 ;
        RECT 220.400 136.300 221.200 136.400 ;
        RECT 215.600 135.700 221.200 136.300 ;
        RECT 215.600 135.600 216.400 135.700 ;
        RECT 220.400 135.600 221.200 135.700 ;
        RECT 226.800 136.300 227.600 136.400 ;
        RECT 231.600 136.300 232.400 136.400 ;
        RECT 226.800 135.700 232.400 136.300 ;
        RECT 226.800 135.600 227.600 135.700 ;
        RECT 231.600 135.600 232.400 135.700 ;
        RECT 236.400 135.600 237.200 136.400 ;
        RECT 238.000 136.300 238.800 136.400 ;
        RECT 241.200 136.300 242.000 136.400 ;
        RECT 244.400 136.300 245.200 136.400 ;
        RECT 238.000 135.700 245.200 136.300 ;
        RECT 238.000 135.600 238.800 135.700 ;
        RECT 241.200 135.600 242.000 135.700 ;
        RECT 244.400 135.600 245.200 135.700 ;
        RECT 135.600 133.700 137.900 134.300 ;
        RECT 135.600 133.600 136.400 133.700 ;
        RECT 177.200 133.600 178.000 134.400 ;
        RECT 190.000 134.300 190.800 134.400 ;
        RECT 204.400 134.300 205.200 134.400 ;
        RECT 212.400 134.300 213.200 134.400 ;
        RECT 217.200 134.300 218.000 134.400 ;
        RECT 190.000 133.700 218.000 134.300 ;
        RECT 190.000 133.600 190.800 133.700 ;
        RECT 204.400 133.600 205.200 133.700 ;
        RECT 212.400 133.600 213.200 133.700 ;
        RECT 217.200 133.600 218.000 133.700 ;
        RECT 220.400 134.300 221.200 134.400 ;
        RECT 238.100 134.300 238.700 135.600 ;
        RECT 220.400 133.700 238.700 134.300 ;
        RECT 220.400 133.600 221.200 133.700 ;
        RECT 46.000 132.300 46.800 132.400 ;
        RECT 54.000 132.300 54.800 132.400 ;
        RECT 62.000 132.300 62.800 132.400 ;
        RECT 46.000 131.700 62.800 132.300 ;
        RECT 46.000 131.600 46.800 131.700 ;
        RECT 54.000 131.600 54.800 131.700 ;
        RECT 62.000 131.600 62.800 131.700 ;
        RECT 81.200 132.300 82.000 132.400 ;
        RECT 87.600 132.300 88.400 132.400 ;
        RECT 81.200 131.700 88.400 132.300 ;
        RECT 81.200 131.600 82.000 131.700 ;
        RECT 87.600 131.600 88.400 131.700 ;
        RECT 177.200 132.300 178.000 132.400 ;
        RECT 196.400 132.300 197.200 132.400 ;
        RECT 177.200 131.700 197.200 132.300 ;
        RECT 177.200 131.600 178.000 131.700 ;
        RECT 196.400 131.600 197.200 131.700 ;
        RECT 199.600 132.300 200.400 132.400 ;
        RECT 202.800 132.300 203.600 132.400 ;
        RECT 199.600 131.700 203.600 132.300 ;
        RECT 199.600 131.600 200.400 131.700 ;
        RECT 202.800 131.600 203.600 131.700 ;
        RECT 222.000 132.300 222.800 132.400 ;
        RECT 226.800 132.300 227.600 132.400 ;
        RECT 222.000 131.700 227.600 132.300 ;
        RECT 222.000 131.600 222.800 131.700 ;
        RECT 226.800 131.600 227.600 131.700 ;
        RECT 233.200 132.300 234.000 132.400 ;
        RECT 238.000 132.300 238.800 132.400 ;
        RECT 233.200 131.700 238.800 132.300 ;
        RECT 233.200 131.600 234.000 131.700 ;
        RECT 238.000 131.600 238.800 131.700 ;
        RECT 49.200 130.300 50.000 130.400 ;
        RECT 74.800 130.300 75.600 130.400 ;
        RECT 49.200 129.700 75.600 130.300 ;
        RECT 49.200 129.600 50.000 129.700 ;
        RECT 74.800 129.600 75.600 129.700 ;
        RECT 98.800 130.300 99.600 130.400 ;
        RECT 111.600 130.300 112.400 130.400 ;
        RECT 98.800 129.700 112.400 130.300 ;
        RECT 98.800 129.600 99.600 129.700 ;
        RECT 111.600 129.600 112.400 129.700 ;
        RECT 166.000 130.300 166.800 130.400 ;
        RECT 178.800 130.300 179.600 130.400 ;
        RECT 166.000 129.700 179.600 130.300 ;
        RECT 166.000 129.600 166.800 129.700 ;
        RECT 178.800 129.600 179.600 129.700 ;
        RECT 206.000 130.300 206.800 130.400 ;
        RECT 234.800 130.300 235.600 130.400 ;
        RECT 238.000 130.300 238.800 130.400 ;
        RECT 206.000 129.700 238.800 130.300 ;
        RECT 206.000 129.600 206.800 129.700 ;
        RECT 234.800 129.600 235.600 129.700 ;
        RECT 238.000 129.600 238.800 129.700 ;
        RECT 62.000 128.300 62.800 128.400 ;
        RECT 86.000 128.300 86.800 128.400 ;
        RECT 62.000 127.700 86.800 128.300 ;
        RECT 62.000 127.600 62.800 127.700 ;
        RECT 86.000 127.600 86.800 127.700 ;
        RECT 199.600 126.300 200.400 126.400 ;
        RECT 202.800 126.300 203.600 126.400 ;
        RECT 199.600 125.700 203.600 126.300 ;
        RECT 199.600 125.600 200.400 125.700 ;
        RECT 202.800 125.600 203.600 125.700 ;
        RECT 44.400 124.300 45.200 124.400 ;
        RECT 50.800 124.300 51.600 124.400 ;
        RECT 78.000 124.300 78.800 124.400 ;
        RECT 44.400 123.700 78.800 124.300 ;
        RECT 44.400 123.600 45.200 123.700 ;
        RECT 50.800 123.600 51.600 123.700 ;
        RECT 78.000 123.600 78.800 123.700 ;
        RECT 76.400 122.300 77.200 122.400 ;
        RECT 94.000 122.300 94.800 122.400 ;
        RECT 127.600 122.300 128.400 122.400 ;
        RECT 76.400 121.700 128.400 122.300 ;
        RECT 76.400 121.600 77.200 121.700 ;
        RECT 94.000 121.600 94.800 121.700 ;
        RECT 127.600 121.600 128.400 121.700 ;
        RECT 154.800 120.300 155.600 120.400 ;
        RECT 174.000 120.300 174.800 120.400 ;
        RECT 154.800 119.700 174.800 120.300 ;
        RECT 154.800 119.600 155.600 119.700 ;
        RECT 174.000 119.600 174.800 119.700 ;
        RECT 58.800 118.300 59.600 118.400 ;
        RECT 63.600 118.300 64.400 118.400 ;
        RECT 58.800 117.700 64.400 118.300 ;
        RECT 58.800 117.600 59.600 117.700 ;
        RECT 63.600 117.600 64.400 117.700 ;
        RECT 127.600 118.300 128.400 118.400 ;
        RECT 132.400 118.300 133.200 118.400 ;
        RECT 127.600 117.700 133.200 118.300 ;
        RECT 127.600 117.600 128.400 117.700 ;
        RECT 132.400 117.600 133.200 117.700 ;
        RECT 162.800 114.300 163.600 114.400 ;
        RECT 234.800 114.300 235.600 114.400 ;
        RECT 162.800 113.700 235.600 114.300 ;
        RECT 162.800 113.600 163.600 113.700 ;
        RECT 234.800 113.600 235.600 113.700 ;
        RECT 52.400 112.300 53.200 112.400 ;
        RECT 60.400 112.300 61.200 112.400 ;
        RECT 79.600 112.300 80.400 112.400 ;
        RECT 52.400 111.700 80.400 112.300 ;
        RECT 52.400 111.600 53.200 111.700 ;
        RECT 60.400 111.600 61.200 111.700 ;
        RECT 79.600 111.600 80.400 111.700 ;
        RECT 148.400 112.300 149.200 112.400 ;
        RECT 164.400 112.300 165.200 112.400 ;
        RECT 148.400 111.700 165.200 112.300 ;
        RECT 148.400 111.600 149.200 111.700 ;
        RECT 164.400 111.600 165.200 111.700 ;
        RECT 201.200 112.300 202.000 112.400 ;
        RECT 214.000 112.300 214.800 112.400 ;
        RECT 201.200 111.700 214.800 112.300 ;
        RECT 201.200 111.600 202.000 111.700 ;
        RECT 214.000 111.600 214.800 111.700 ;
        RECT 42.800 109.600 43.600 110.400 ;
        RECT 71.600 110.300 72.400 110.400 ;
        RECT 74.800 110.300 75.600 110.400 ;
        RECT 89.200 110.300 90.000 110.400 ;
        RECT 71.600 109.700 90.000 110.300 ;
        RECT 71.600 109.600 72.400 109.700 ;
        RECT 74.800 109.600 75.600 109.700 ;
        RECT 89.200 109.600 90.000 109.700 ;
        RECT 135.600 110.300 136.400 110.400 ;
        RECT 145.200 110.300 146.000 110.400 ;
        RECT 135.600 109.700 146.000 110.300 ;
        RECT 135.600 109.600 136.400 109.700 ;
        RECT 145.200 109.600 146.000 109.700 ;
        RECT 148.400 110.300 149.200 110.400 ;
        RECT 151.600 110.300 152.400 110.400 ;
        RECT 148.400 109.700 152.400 110.300 ;
        RECT 148.400 109.600 149.200 109.700 ;
        RECT 151.600 109.600 152.400 109.700 ;
        RECT 161.200 110.300 162.000 110.400 ;
        RECT 174.000 110.300 174.800 110.400 ;
        RECT 177.200 110.300 178.000 110.400 ;
        RECT 161.200 109.700 178.000 110.300 ;
        RECT 161.200 109.600 162.000 109.700 ;
        RECT 174.000 109.600 174.800 109.700 ;
        RECT 177.200 109.600 178.000 109.700 ;
        RECT 196.400 110.300 197.200 110.400 ;
        RECT 247.600 110.300 248.400 110.400 ;
        RECT 196.400 109.700 248.400 110.300 ;
        RECT 196.400 109.600 197.200 109.700 ;
        RECT 247.600 109.600 248.400 109.700 ;
        RECT 42.800 108.300 43.600 108.400 ;
        RECT 50.800 108.300 51.600 108.400 ;
        RECT 42.800 107.700 51.600 108.300 ;
        RECT 42.800 107.600 43.600 107.700 ;
        RECT 50.800 107.600 51.600 107.700 ;
        RECT 54.000 108.300 54.800 108.400 ;
        RECT 58.800 108.300 59.600 108.400 ;
        RECT 54.000 107.700 59.600 108.300 ;
        RECT 54.000 107.600 54.800 107.700 ;
        RECT 58.800 107.600 59.600 107.700 ;
        RECT 90.800 108.300 91.600 108.400 ;
        RECT 108.400 108.300 109.200 108.400 ;
        RECT 90.800 107.700 109.200 108.300 ;
        RECT 90.800 107.600 91.600 107.700 ;
        RECT 108.400 107.600 109.200 107.700 ;
        RECT 134.000 108.300 134.800 108.400 ;
        RECT 143.600 108.300 144.400 108.400 ;
        RECT 148.400 108.300 149.200 108.400 ;
        RECT 156.400 108.300 157.200 108.400 ;
        RECT 166.000 108.300 166.800 108.400 ;
        RECT 134.000 107.700 166.800 108.300 ;
        RECT 134.000 107.600 134.800 107.700 ;
        RECT 143.600 107.600 144.400 107.700 ;
        RECT 148.400 107.600 149.200 107.700 ;
        RECT 156.400 107.600 157.200 107.700 ;
        RECT 166.000 107.600 166.800 107.700 ;
        RECT 178.800 108.300 179.600 108.400 ;
        RECT 183.600 108.300 184.400 108.400 ;
        RECT 178.800 107.700 184.400 108.300 ;
        RECT 178.800 107.600 179.600 107.700 ;
        RECT 183.600 107.600 184.400 107.700 ;
        RECT 204.400 108.300 205.200 108.400 ;
        RECT 222.000 108.300 222.800 108.400 ;
        RECT 204.400 107.700 222.800 108.300 ;
        RECT 204.400 107.600 205.200 107.700 ;
        RECT 222.000 107.600 222.800 107.700 ;
        RECT 7.600 106.300 8.400 106.400 ;
        RECT 47.600 106.300 48.400 106.400 ;
        RECT 7.600 105.700 48.400 106.300 ;
        RECT 7.600 105.600 8.400 105.700 ;
        RECT 47.600 105.600 48.400 105.700 ;
        RECT 57.200 106.300 58.000 106.400 ;
        RECT 60.400 106.300 61.200 106.400 ;
        RECT 57.200 105.700 61.200 106.300 ;
        RECT 57.200 105.600 58.000 105.700 ;
        RECT 60.400 105.600 61.200 105.700 ;
        RECT 130.800 106.300 131.600 106.400 ;
        RECT 150.000 106.300 150.800 106.400 ;
        RECT 130.800 105.700 150.800 106.300 ;
        RECT 130.800 105.600 131.600 105.700 ;
        RECT 150.000 105.600 150.800 105.700 ;
        RECT 153.200 106.300 154.000 106.400 ;
        RECT 158.000 106.300 158.800 106.400 ;
        RECT 153.200 105.700 158.800 106.300 ;
        RECT 153.200 105.600 154.000 105.700 ;
        RECT 158.000 105.600 158.800 105.700 ;
        RECT 190.000 106.300 190.800 106.400 ;
        RECT 198.000 106.300 198.800 106.400 ;
        RECT 190.000 105.700 198.800 106.300 ;
        RECT 190.000 105.600 190.800 105.700 ;
        RECT 198.000 105.600 198.800 105.700 ;
        RECT 209.200 106.300 210.000 106.400 ;
        RECT 212.400 106.300 213.200 106.400 ;
        RECT 209.200 105.700 213.200 106.300 ;
        RECT 209.200 105.600 210.000 105.700 ;
        RECT 212.400 105.600 213.200 105.700 ;
        RECT 218.800 106.300 219.600 106.400 ;
        RECT 225.200 106.300 226.000 106.400 ;
        RECT 218.800 105.700 226.000 106.300 ;
        RECT 218.800 105.600 219.600 105.700 ;
        RECT 225.200 105.600 226.000 105.700 ;
        RECT 26.800 104.300 27.600 104.400 ;
        RECT 44.400 104.300 45.200 104.400 ;
        RECT 26.800 103.700 45.200 104.300 ;
        RECT 26.800 103.600 27.600 103.700 ;
        RECT 44.400 103.600 45.200 103.700 ;
        RECT 78.000 104.300 78.800 104.400 ;
        RECT 87.600 104.300 88.400 104.400 ;
        RECT 78.000 103.700 88.400 104.300 ;
        RECT 78.000 103.600 78.800 103.700 ;
        RECT 87.600 103.600 88.400 103.700 ;
        RECT 129.200 104.300 130.000 104.400 ;
        RECT 159.600 104.300 160.400 104.400 ;
        RECT 129.200 103.700 160.400 104.300 ;
        RECT 129.200 103.600 130.000 103.700 ;
        RECT 159.600 103.600 160.400 103.700 ;
        RECT 177.200 104.300 178.000 104.400 ;
        RECT 212.400 104.300 213.200 104.400 ;
        RECT 239.600 104.300 240.400 104.400 ;
        RECT 177.200 103.700 240.400 104.300 ;
        RECT 177.200 103.600 178.000 103.700 ;
        RECT 212.400 103.600 213.200 103.700 ;
        RECT 239.600 103.600 240.400 103.700 ;
        RECT 74.800 102.300 75.600 102.400 ;
        RECT 92.400 102.300 93.200 102.400 ;
        RECT 100.400 102.300 101.200 102.400 ;
        RECT 140.400 102.300 141.200 102.400 ;
        RECT 154.800 102.300 155.600 102.400 ;
        RECT 159.600 102.300 160.400 102.400 ;
        RECT 74.800 101.700 160.400 102.300 ;
        RECT 74.800 101.600 75.600 101.700 ;
        RECT 92.400 101.600 93.200 101.700 ;
        RECT 100.400 101.600 101.200 101.700 ;
        RECT 140.400 101.600 141.200 101.700 ;
        RECT 154.800 101.600 155.600 101.700 ;
        RECT 159.600 101.600 160.400 101.700 ;
        RECT 194.800 102.300 195.600 102.400 ;
        RECT 202.800 102.300 203.600 102.400 ;
        RECT 194.800 101.700 203.600 102.300 ;
        RECT 194.800 101.600 195.600 101.700 ;
        RECT 202.800 101.600 203.600 101.700 ;
        RECT 206.000 102.300 206.800 102.400 ;
        RECT 226.800 102.300 227.600 102.400 ;
        RECT 206.000 101.700 227.600 102.300 ;
        RECT 206.000 101.600 206.800 101.700 ;
        RECT 226.800 101.600 227.600 101.700 ;
        RECT 238.000 102.300 238.800 102.400 ;
        RECT 241.200 102.300 242.000 102.400 ;
        RECT 238.000 101.700 242.000 102.300 ;
        RECT 238.000 101.600 238.800 101.700 ;
        RECT 241.200 101.600 242.000 101.700 ;
        RECT 76.400 100.300 77.200 100.400 ;
        RECT 79.600 100.300 80.400 100.400 ;
        RECT 76.400 99.700 80.400 100.300 ;
        RECT 76.400 99.600 77.200 99.700 ;
        RECT 79.600 99.600 80.400 99.700 ;
        RECT 116.400 100.300 117.200 100.400 ;
        RECT 158.000 100.300 158.800 100.400 ;
        RECT 170.800 100.300 171.600 100.400 ;
        RECT 177.200 100.300 178.000 100.400 ;
        RECT 116.400 99.700 178.000 100.300 ;
        RECT 116.400 99.600 117.200 99.700 ;
        RECT 158.000 99.600 158.800 99.700 ;
        RECT 170.800 99.600 171.600 99.700 ;
        RECT 177.200 99.600 178.000 99.700 ;
        RECT 76.400 98.300 77.200 98.400 ;
        RECT 78.000 98.300 78.800 98.400 ;
        RECT 76.400 97.700 78.800 98.300 ;
        RECT 76.400 97.600 77.200 97.700 ;
        RECT 78.000 97.600 78.800 97.700 ;
        RECT 98.800 98.300 99.600 98.400 ;
        RECT 111.600 98.300 112.400 98.400 ;
        RECT 132.400 98.300 133.200 98.400 ;
        RECT 98.800 97.700 133.200 98.300 ;
        RECT 98.800 97.600 99.600 97.700 ;
        RECT 111.600 97.600 112.400 97.700 ;
        RECT 132.400 97.600 133.200 97.700 ;
        RECT 167.600 98.300 168.400 98.400 ;
        RECT 170.800 98.300 171.600 98.400 ;
        RECT 175.600 98.300 176.400 98.400 ;
        RECT 196.400 98.300 197.200 98.400 ;
        RECT 167.600 97.700 197.200 98.300 ;
        RECT 167.600 97.600 168.400 97.700 ;
        RECT 170.800 97.600 171.600 97.700 ;
        RECT 175.600 97.600 176.400 97.700 ;
        RECT 196.400 97.600 197.200 97.700 ;
        RECT 201.200 98.300 202.000 98.400 ;
        RECT 207.600 98.300 208.400 98.400 ;
        RECT 201.200 97.700 208.400 98.300 ;
        RECT 201.200 97.600 202.000 97.700 ;
        RECT 207.600 97.600 208.400 97.700 ;
        RECT 210.800 98.300 211.600 98.400 ;
        RECT 225.200 98.300 226.000 98.400 ;
        RECT 210.800 97.700 226.000 98.300 ;
        RECT 210.800 97.600 211.600 97.700 ;
        RECT 225.200 97.600 226.000 97.700 ;
        RECT 228.400 98.300 229.200 98.400 ;
        RECT 247.600 98.300 248.400 98.400 ;
        RECT 228.400 97.700 248.400 98.300 ;
        RECT 228.400 97.600 229.200 97.700 ;
        RECT 247.600 97.600 248.400 97.700 ;
        RECT 42.800 96.300 43.600 96.400 ;
        RECT 44.400 96.300 45.200 96.400 ;
        RECT 42.800 95.700 45.200 96.300 ;
        RECT 42.800 95.600 43.600 95.700 ;
        RECT 44.400 95.600 45.200 95.700 ;
        RECT 161.200 96.300 162.000 96.400 ;
        RECT 164.400 96.300 165.200 96.400 ;
        RECT 161.200 95.700 165.200 96.300 ;
        RECT 161.200 95.600 162.000 95.700 ;
        RECT 164.400 95.600 165.200 95.700 ;
        RECT 169.200 96.300 170.000 96.400 ;
        RECT 180.400 96.300 181.200 96.400 ;
        RECT 169.200 95.700 181.200 96.300 ;
        RECT 169.200 95.600 170.000 95.700 ;
        RECT 180.400 95.600 181.200 95.700 ;
        RECT 206.000 96.300 206.800 96.400 ;
        RECT 214.000 96.300 214.800 96.400 ;
        RECT 206.000 95.700 214.800 96.300 ;
        RECT 206.000 95.600 206.800 95.700 ;
        RECT 214.000 95.600 214.800 95.700 ;
        RECT 217.200 96.300 218.000 96.400 ;
        RECT 222.000 96.300 222.800 96.400 ;
        RECT 217.200 95.700 222.800 96.300 ;
        RECT 217.200 95.600 218.000 95.700 ;
        RECT 222.000 95.600 222.800 95.700 ;
        RECT 241.200 96.300 242.000 96.400 ;
        RECT 246.000 96.300 246.800 96.400 ;
        RECT 241.200 95.700 246.800 96.300 ;
        RECT 241.200 95.600 242.000 95.700 ;
        RECT 246.000 95.600 246.800 95.700 ;
        RECT 26.800 94.300 27.600 94.400 ;
        RECT 42.800 94.300 43.600 94.400 ;
        RECT 26.800 93.700 43.600 94.300 ;
        RECT 26.800 93.600 27.600 93.700 ;
        RECT 42.800 93.600 43.600 93.700 ;
        RECT 47.600 94.300 48.400 94.400 ;
        RECT 62.000 94.300 62.800 94.400 ;
        RECT 47.600 93.700 62.800 94.300 ;
        RECT 47.600 93.600 48.400 93.700 ;
        RECT 62.000 93.600 62.800 93.700 ;
        RECT 73.200 94.300 74.000 94.400 ;
        RECT 102.000 94.300 102.800 94.400 ;
        RECT 73.200 93.700 102.800 94.300 ;
        RECT 73.200 93.600 74.000 93.700 ;
        RECT 102.000 93.600 102.800 93.700 ;
        RECT 150.000 94.300 150.800 94.400 ;
        RECT 174.000 94.300 174.800 94.400 ;
        RECT 198.000 94.300 198.800 94.400 ;
        RECT 223.600 94.300 224.400 94.400 ;
        RECT 150.000 93.700 224.400 94.300 ;
        RECT 150.000 93.600 150.800 93.700 ;
        RECT 174.000 93.600 174.800 93.700 ;
        RECT 198.000 93.600 198.800 93.700 ;
        RECT 223.600 93.600 224.400 93.700 ;
        RECT 225.200 94.300 226.000 94.400 ;
        RECT 230.000 94.300 230.800 94.400 ;
        RECT 225.200 93.700 230.800 94.300 ;
        RECT 225.200 93.600 226.000 93.700 ;
        RECT 230.000 93.600 230.800 93.700 ;
        RECT 242.800 94.300 243.600 94.400 ;
        RECT 249.200 94.300 250.000 94.400 ;
        RECT 242.800 93.700 250.000 94.300 ;
        RECT 242.800 93.600 243.600 93.700 ;
        RECT 249.200 93.600 250.000 93.700 ;
        RECT 36.400 92.300 37.200 92.400 ;
        RECT 79.600 92.300 80.400 92.400 ;
        RECT 36.400 91.700 80.400 92.300 ;
        RECT 36.400 91.600 37.200 91.700 ;
        RECT 79.600 91.600 80.400 91.700 ;
        RECT 113.200 92.300 114.000 92.400 ;
        RECT 119.600 92.300 120.400 92.400 ;
        RECT 113.200 91.700 120.400 92.300 ;
        RECT 113.200 91.600 114.000 91.700 ;
        RECT 119.600 91.600 120.400 91.700 ;
        RECT 129.200 92.300 130.000 92.400 ;
        RECT 146.800 92.300 147.600 92.400 ;
        RECT 188.400 92.300 189.200 92.400 ;
        RECT 129.200 91.700 189.200 92.300 ;
        RECT 129.200 91.600 130.000 91.700 ;
        RECT 146.800 91.600 147.600 91.700 ;
        RECT 188.400 91.600 189.200 91.700 ;
        RECT 191.600 92.300 192.400 92.400 ;
        RECT 199.600 92.300 200.400 92.400 ;
        RECT 234.800 92.300 235.600 92.400 ;
        RECT 191.600 91.700 235.600 92.300 ;
        RECT 191.600 91.600 192.400 91.700 ;
        RECT 199.600 91.600 200.400 91.700 ;
        RECT 234.800 91.600 235.600 91.700 ;
        RECT 7.600 90.300 8.400 90.400 ;
        RECT 58.800 90.300 59.600 90.400 ;
        RECT 7.600 89.700 59.600 90.300 ;
        RECT 7.600 89.600 8.400 89.700 ;
        RECT 58.800 89.600 59.600 89.700 ;
        RECT 169.200 90.300 170.000 90.400 ;
        RECT 175.600 90.300 176.400 90.400 ;
        RECT 169.200 89.700 176.400 90.300 ;
        RECT 169.200 89.600 170.000 89.700 ;
        RECT 175.600 89.600 176.400 89.700 ;
        RECT 193.200 90.300 194.000 90.400 ;
        RECT 196.400 90.300 197.200 90.400 ;
        RECT 217.200 90.300 218.000 90.400 ;
        RECT 193.200 89.700 218.000 90.300 ;
        RECT 193.200 89.600 194.000 89.700 ;
        RECT 196.400 89.600 197.200 89.700 ;
        RECT 217.200 89.600 218.000 89.700 ;
        RECT 218.800 90.300 219.600 90.400 ;
        RECT 238.000 90.300 238.800 90.400 ;
        RECT 218.800 89.700 238.800 90.300 ;
        RECT 218.800 89.600 219.600 89.700 ;
        RECT 238.000 89.600 238.800 89.700 ;
        RECT 159.600 88.300 160.400 88.400 ;
        RECT 207.600 88.300 208.400 88.400 ;
        RECT 159.600 87.700 208.400 88.300 ;
        RECT 159.600 87.600 160.400 87.700 ;
        RECT 207.600 87.600 208.400 87.700 ;
        RECT 210.800 88.300 211.600 88.400 ;
        RECT 214.000 88.300 214.800 88.400 ;
        RECT 210.800 87.700 214.800 88.300 ;
        RECT 210.800 87.600 211.600 87.700 ;
        RECT 214.000 87.600 214.800 87.700 ;
        RECT 52.400 86.300 53.200 86.400 ;
        RECT 74.800 86.300 75.600 86.400 ;
        RECT 52.400 85.700 75.600 86.300 ;
        RECT 52.400 85.600 53.200 85.700 ;
        RECT 74.800 85.600 75.600 85.700 ;
        RECT 154.800 86.300 155.600 86.400 ;
        RECT 172.400 86.300 173.200 86.400 ;
        RECT 154.800 85.700 173.200 86.300 ;
        RECT 154.800 85.600 155.600 85.700 ;
        RECT 172.400 85.600 173.200 85.700 ;
        RECT 142.000 84.300 142.800 84.400 ;
        RECT 148.400 84.300 149.200 84.400 ;
        RECT 142.000 83.700 149.200 84.300 ;
        RECT 142.000 83.600 142.800 83.700 ;
        RECT 148.400 83.600 149.200 83.700 ;
        RECT 17.200 82.300 18.000 82.400 ;
        RECT 23.600 82.300 24.400 82.400 ;
        RECT 17.200 81.700 24.400 82.300 ;
        RECT 17.200 81.600 18.000 81.700 ;
        RECT 23.600 81.600 24.400 81.700 ;
        RECT 145.200 82.300 146.000 82.400 ;
        RECT 191.600 82.300 192.400 82.400 ;
        RECT 145.200 81.700 192.400 82.300 ;
        RECT 145.200 81.600 146.000 81.700 ;
        RECT 191.600 81.600 192.400 81.700 ;
        RECT 124.400 78.300 125.200 78.400 ;
        RECT 154.800 78.300 155.600 78.400 ;
        RECT 124.400 77.700 155.600 78.300 ;
        RECT 124.400 77.600 125.200 77.700 ;
        RECT 154.800 77.600 155.600 77.700 ;
        RECT 198.000 78.300 198.800 78.400 ;
        RECT 202.800 78.300 203.600 78.400 ;
        RECT 198.000 77.700 203.600 78.300 ;
        RECT 198.000 77.600 198.800 77.700 ;
        RECT 202.800 77.600 203.600 77.700 ;
        RECT 217.200 78.300 218.000 78.400 ;
        RECT 222.000 78.300 222.800 78.400 ;
        RECT 217.200 77.700 222.800 78.300 ;
        RECT 217.200 77.600 218.000 77.700 ;
        RECT 222.000 77.600 222.800 77.700 ;
        RECT 97.200 76.300 98.000 76.400 ;
        RECT 151.600 76.300 152.400 76.400 ;
        RECT 97.200 75.700 152.400 76.300 ;
        RECT 97.200 75.600 98.000 75.700 ;
        RECT 151.600 75.600 152.400 75.700 ;
        RECT 154.800 76.300 155.600 76.400 ;
        RECT 161.200 76.300 162.000 76.400 ;
        RECT 154.800 75.700 162.000 76.300 ;
        RECT 154.800 75.600 155.600 75.700 ;
        RECT 161.200 75.600 162.000 75.700 ;
        RECT 196.400 76.300 197.200 76.400 ;
        RECT 201.200 76.300 202.000 76.400 ;
        RECT 222.000 76.300 222.800 76.400 ;
        RECT 196.400 75.700 222.800 76.300 ;
        RECT 196.400 75.600 197.200 75.700 ;
        RECT 201.200 75.600 202.000 75.700 ;
        RECT 222.000 75.600 222.800 75.700 ;
        RECT 36.400 74.300 37.200 74.400 ;
        RECT 41.200 74.300 42.000 74.400 ;
        RECT 50.800 74.300 51.600 74.400 ;
        RECT 36.400 73.700 51.600 74.300 ;
        RECT 36.400 73.600 37.200 73.700 ;
        RECT 41.200 73.600 42.000 73.700 ;
        RECT 50.800 73.600 51.600 73.700 ;
        RECT 57.200 74.300 58.000 74.400 ;
        RECT 60.400 74.300 61.200 74.400 ;
        RECT 154.800 74.300 155.600 74.400 ;
        RECT 57.200 73.700 155.600 74.300 ;
        RECT 57.200 73.600 58.000 73.700 ;
        RECT 60.400 73.600 61.200 73.700 ;
        RECT 154.800 73.600 155.600 73.700 ;
        RECT 239.600 74.300 240.400 74.400 ;
        RECT 242.800 74.300 243.600 74.400 ;
        RECT 239.600 73.700 243.600 74.300 ;
        RECT 239.600 73.600 240.400 73.700 ;
        RECT 242.800 73.600 243.600 73.700 ;
        RECT 246.000 74.300 246.800 74.400 ;
        RECT 250.800 74.300 251.600 74.400 ;
        RECT 246.000 73.700 251.600 74.300 ;
        RECT 246.000 73.600 246.800 73.700 ;
        RECT 250.800 73.600 251.600 73.700 ;
        RECT 7.600 72.300 8.400 72.400 ;
        RECT 38.000 72.300 38.800 72.400 ;
        RECT 46.000 72.300 46.800 72.400 ;
        RECT 7.600 71.700 46.800 72.300 ;
        RECT 7.600 71.600 8.400 71.700 ;
        RECT 38.000 71.600 38.800 71.700 ;
        RECT 46.000 71.600 46.800 71.700 ;
        RECT 116.400 72.300 117.200 72.400 ;
        RECT 122.800 72.300 123.600 72.400 ;
        RECT 116.400 71.700 123.600 72.300 ;
        RECT 116.400 71.600 117.200 71.700 ;
        RECT 122.800 71.600 123.600 71.700 ;
        RECT 138.800 72.300 139.600 72.400 ;
        RECT 148.400 72.300 149.200 72.400 ;
        RECT 138.800 71.700 149.200 72.300 ;
        RECT 138.800 71.600 139.600 71.700 ;
        RECT 148.400 71.600 149.200 71.700 ;
        RECT 162.800 72.300 163.600 72.400 ;
        RECT 174.000 72.300 174.800 72.400 ;
        RECT 162.800 71.700 174.800 72.300 ;
        RECT 162.800 71.600 163.600 71.700 ;
        RECT 174.000 71.600 174.800 71.700 ;
        RECT 201.200 72.300 202.000 72.400 ;
        RECT 218.800 72.300 219.600 72.400 ;
        RECT 201.200 71.700 219.600 72.300 ;
        RECT 201.200 71.600 202.000 71.700 ;
        RECT 218.800 71.600 219.600 71.700 ;
        RECT 226.800 72.300 227.600 72.400 ;
        RECT 244.400 72.300 245.200 72.400 ;
        RECT 226.800 71.700 245.200 72.300 ;
        RECT 226.800 71.600 227.600 71.700 ;
        RECT 244.400 71.600 245.200 71.700 ;
        RECT 39.600 70.300 40.400 70.400 ;
        RECT 52.400 70.300 53.200 70.400 ;
        RECT 39.600 69.700 53.200 70.300 ;
        RECT 39.600 69.600 40.400 69.700 ;
        RECT 52.400 69.600 53.200 69.700 ;
        RECT 82.800 70.300 83.600 70.400 ;
        RECT 126.000 70.300 126.800 70.400 ;
        RECT 82.800 69.700 126.800 70.300 ;
        RECT 82.800 69.600 83.600 69.700 ;
        RECT 126.000 69.600 126.800 69.700 ;
        RECT 220.400 70.300 221.200 70.400 ;
        RECT 228.400 70.300 229.200 70.400 ;
        RECT 220.400 69.700 229.200 70.300 ;
        RECT 220.400 69.600 221.200 69.700 ;
        RECT 228.400 69.600 229.200 69.700 ;
        RECT 231.600 70.300 232.400 70.400 ;
        RECT 244.400 70.300 245.200 70.400 ;
        RECT 247.600 70.300 248.400 70.400 ;
        RECT 231.600 69.700 248.400 70.300 ;
        RECT 231.600 69.600 232.400 69.700 ;
        RECT 244.400 69.600 245.200 69.700 ;
        RECT 247.600 69.600 248.400 69.700 ;
        RECT 42.800 68.300 43.600 68.400 ;
        RECT 47.600 68.300 48.400 68.400 ;
        RECT 55.600 68.300 56.400 68.400 ;
        RECT 71.600 68.300 72.400 68.400 ;
        RECT 42.800 67.700 72.400 68.300 ;
        RECT 42.800 67.600 43.600 67.700 ;
        RECT 47.600 67.600 48.400 67.700 ;
        RECT 55.600 67.600 56.400 67.700 ;
        RECT 71.600 67.600 72.400 67.700 ;
        RECT 135.600 68.300 136.400 68.400 ;
        RECT 150.000 68.300 150.800 68.400 ;
        RECT 154.800 68.300 155.600 68.400 ;
        RECT 135.600 67.700 155.600 68.300 ;
        RECT 135.600 67.600 136.400 67.700 ;
        RECT 150.000 67.600 150.800 67.700 ;
        RECT 154.800 67.600 155.600 67.700 ;
        RECT 156.400 68.300 157.200 68.400 ;
        RECT 162.800 68.300 163.600 68.400 ;
        RECT 156.400 67.700 163.600 68.300 ;
        RECT 156.400 67.600 157.200 67.700 ;
        RECT 162.800 67.600 163.600 67.700 ;
        RECT 166.000 68.300 166.800 68.400 ;
        RECT 177.200 68.300 178.000 68.400 ;
        RECT 230.000 68.300 230.800 68.400 ;
        RECT 166.000 67.700 230.800 68.300 ;
        RECT 166.000 67.600 166.800 67.700 ;
        RECT 177.200 67.600 178.000 67.700 ;
        RECT 230.000 67.600 230.800 67.700 ;
        RECT 100.400 66.300 101.200 66.400 ;
        RECT 121.200 66.300 122.000 66.400 ;
        RECT 100.400 65.700 122.000 66.300 ;
        RECT 100.400 65.600 101.200 65.700 ;
        RECT 121.200 65.600 122.000 65.700 ;
        RECT 161.200 66.300 162.000 66.400 ;
        RECT 167.600 66.300 168.400 66.400 ;
        RECT 161.200 65.700 168.400 66.300 ;
        RECT 161.200 65.600 162.000 65.700 ;
        RECT 167.600 65.600 168.400 65.700 ;
        RECT 169.200 66.300 170.000 66.400 ;
        RECT 225.200 66.300 226.000 66.400 ;
        RECT 169.200 65.700 226.000 66.300 ;
        RECT 169.200 65.600 170.000 65.700 ;
        RECT 225.200 65.600 226.000 65.700 ;
        RECT 174.000 64.300 174.800 64.400 ;
        RECT 191.600 64.300 192.400 64.400 ;
        RECT 174.000 63.700 192.400 64.300 ;
        RECT 174.000 63.600 174.800 63.700 ;
        RECT 191.600 63.600 192.400 63.700 ;
        RECT 217.200 64.300 218.000 64.400 ;
        RECT 246.000 64.300 246.800 64.400 ;
        RECT 217.200 63.700 246.800 64.300 ;
        RECT 217.200 63.600 218.000 63.700 ;
        RECT 246.000 63.600 246.800 63.700 ;
        RECT 4.400 62.300 5.200 62.400 ;
        RECT 34.800 62.300 35.600 62.400 ;
        RECT 46.000 62.300 46.800 62.400 ;
        RECT 49.200 62.300 50.000 62.400 ;
        RECT 4.400 61.700 50.000 62.300 ;
        RECT 4.400 61.600 5.200 61.700 ;
        RECT 34.800 61.600 35.600 61.700 ;
        RECT 46.000 61.600 46.800 61.700 ;
        RECT 49.200 61.600 50.000 61.700 ;
        RECT 230.000 62.300 230.800 62.400 ;
        RECT 241.200 62.300 242.000 62.400 ;
        RECT 230.000 61.700 242.000 62.300 ;
        RECT 230.000 61.600 230.800 61.700 ;
        RECT 241.200 61.600 242.000 61.700 ;
        RECT 26.800 60.300 27.600 60.400 ;
        RECT 31.600 60.300 32.400 60.400 ;
        RECT 62.000 60.300 62.800 60.400 ;
        RECT 26.800 59.700 62.800 60.300 ;
        RECT 26.800 59.600 27.600 59.700 ;
        RECT 31.600 59.600 32.400 59.700 ;
        RECT 62.000 59.600 62.800 59.700 ;
        RECT 138.800 60.300 139.600 60.400 ;
        RECT 153.200 60.300 154.000 60.400 ;
        RECT 174.000 60.300 174.800 60.400 ;
        RECT 138.800 59.700 174.800 60.300 ;
        RECT 138.800 59.600 139.600 59.700 ;
        RECT 153.200 59.600 154.000 59.700 ;
        RECT 174.000 59.600 174.800 59.700 ;
        RECT 204.400 60.300 205.200 60.400 ;
        RECT 239.600 60.300 240.400 60.400 ;
        RECT 242.800 60.300 243.600 60.400 ;
        RECT 204.400 59.700 243.600 60.300 ;
        RECT 204.400 59.600 205.200 59.700 ;
        RECT 239.600 59.600 240.400 59.700 ;
        RECT 242.800 59.600 243.600 59.700 ;
        RECT 6.000 56.300 6.800 56.400 ;
        RECT 9.200 56.300 10.000 56.400 ;
        RECT 6.000 55.700 10.000 56.300 ;
        RECT 6.000 55.600 6.800 55.700 ;
        RECT 9.200 55.600 10.000 55.700 ;
        RECT 30.000 56.300 30.800 56.400 ;
        RECT 42.800 56.300 43.600 56.400 ;
        RECT 30.000 55.700 43.600 56.300 ;
        RECT 30.000 55.600 30.800 55.700 ;
        RECT 42.800 55.600 43.600 55.700 ;
        RECT 137.200 56.300 138.000 56.400 ;
        RECT 142.000 56.300 142.800 56.400 ;
        RECT 161.200 56.300 162.000 56.400 ;
        RECT 137.200 55.700 162.000 56.300 ;
        RECT 137.200 55.600 138.000 55.700 ;
        RECT 142.000 55.600 142.800 55.700 ;
        RECT 161.200 55.600 162.000 55.700 ;
        RECT 38.000 54.300 38.800 54.400 ;
        RECT 46.000 54.300 46.800 54.400 ;
        RECT 38.000 53.700 46.800 54.300 ;
        RECT 38.000 53.600 38.800 53.700 ;
        RECT 46.000 53.600 46.800 53.700 ;
        RECT 47.600 54.300 48.400 54.400 ;
        RECT 65.200 54.300 66.000 54.400 ;
        RECT 47.600 53.700 66.000 54.300 ;
        RECT 47.600 53.600 48.400 53.700 ;
        RECT 65.200 53.600 66.000 53.700 ;
        RECT 87.600 54.300 88.400 54.400 ;
        RECT 95.600 54.300 96.400 54.400 ;
        RECT 102.000 54.300 102.800 54.400 ;
        RECT 87.600 53.700 102.800 54.300 ;
        RECT 87.600 53.600 88.400 53.700 ;
        RECT 95.600 53.600 96.400 53.700 ;
        RECT 102.000 53.600 102.800 53.700 ;
        RECT 103.600 54.300 104.400 54.400 ;
        RECT 138.800 54.300 139.600 54.400 ;
        RECT 103.600 53.700 139.600 54.300 ;
        RECT 103.600 53.600 104.400 53.700 ;
        RECT 138.800 53.600 139.600 53.700 ;
        RECT 172.400 54.300 173.200 54.400 ;
        RECT 196.400 54.300 197.200 54.400 ;
        RECT 172.400 53.700 197.200 54.300 ;
        RECT 172.400 53.600 173.200 53.700 ;
        RECT 196.400 53.600 197.200 53.700 ;
        RECT 242.800 54.300 243.600 54.400 ;
        RECT 252.400 54.300 253.200 54.400 ;
        RECT 242.800 53.700 253.200 54.300 ;
        RECT 242.800 53.600 243.600 53.700 ;
        RECT 252.400 53.600 253.200 53.700 ;
        RECT 39.600 52.300 40.400 52.400 ;
        RECT 54.000 52.300 54.800 52.400 ;
        RECT 39.600 51.700 54.800 52.300 ;
        RECT 39.600 51.600 40.400 51.700 ;
        RECT 54.000 51.600 54.800 51.700 ;
        RECT 74.800 52.300 75.600 52.400 ;
        RECT 76.400 52.300 77.200 52.400 ;
        RECT 79.600 52.300 80.400 52.400 ;
        RECT 74.800 51.700 80.400 52.300 ;
        RECT 74.800 51.600 75.600 51.700 ;
        RECT 76.400 51.600 77.200 51.700 ;
        RECT 79.600 51.600 80.400 51.700 ;
        RECT 82.800 52.300 83.600 52.400 ;
        RECT 89.200 52.300 90.000 52.400 ;
        RECT 94.000 52.300 94.800 52.400 ;
        RECT 82.800 51.700 94.800 52.300 ;
        RECT 82.800 51.600 83.600 51.700 ;
        RECT 89.200 51.600 90.000 51.700 ;
        RECT 94.000 51.600 94.800 51.700 ;
        RECT 100.400 51.600 101.200 52.400 ;
        RECT 196.400 52.300 197.200 52.400 ;
        RECT 201.200 52.300 202.000 52.400 ;
        RECT 196.400 51.700 202.000 52.300 ;
        RECT 196.400 51.600 197.200 51.700 ;
        RECT 201.200 51.600 202.000 51.700 ;
        RECT 244.400 52.300 245.200 52.400 ;
        RECT 252.400 52.300 253.200 52.400 ;
        RECT 244.400 51.700 253.200 52.300 ;
        RECT 244.400 51.600 245.200 51.700 ;
        RECT 252.400 51.600 253.200 51.700 ;
        RECT 196.400 49.600 197.200 50.400 ;
        RECT 207.600 50.300 208.400 50.400 ;
        RECT 234.800 50.300 235.600 50.400 ;
        RECT 207.600 49.700 235.600 50.300 ;
        RECT 207.600 49.600 208.400 49.700 ;
        RECT 234.800 49.600 235.600 49.700 ;
        RECT 154.800 48.300 155.600 48.400 ;
        RECT 199.600 48.300 200.400 48.400 ;
        RECT 154.800 47.700 200.400 48.300 ;
        RECT 154.800 47.600 155.600 47.700 ;
        RECT 199.600 47.600 200.400 47.700 ;
        RECT 164.400 42.300 165.200 42.400 ;
        RECT 169.200 42.300 170.000 42.400 ;
        RECT 164.400 41.700 170.000 42.300 ;
        RECT 164.400 41.600 165.200 41.700 ;
        RECT 169.200 41.600 170.000 41.700 ;
        RECT 78.000 38.300 78.800 38.400 ;
        RECT 108.400 38.300 109.200 38.400 ;
        RECT 78.000 37.700 109.200 38.300 ;
        RECT 78.000 37.600 78.800 37.700 ;
        RECT 108.400 37.600 109.200 37.700 ;
        RECT 44.400 32.300 45.200 32.400 ;
        RECT 50.800 32.300 51.600 32.400 ;
        RECT 44.400 31.700 51.600 32.300 ;
        RECT 44.400 31.600 45.200 31.700 ;
        RECT 50.800 31.600 51.600 31.700 ;
        RECT 172.400 32.300 173.200 32.400 ;
        RECT 210.800 32.300 211.600 32.400 ;
        RECT 215.600 32.300 216.400 32.400 ;
        RECT 172.400 31.700 216.400 32.300 ;
        RECT 172.400 31.600 173.200 31.700 ;
        RECT 210.800 31.600 211.600 31.700 ;
        RECT 215.600 31.600 216.400 31.700 ;
        RECT 23.600 30.300 24.400 30.400 ;
        RECT 26.800 30.300 27.600 30.400 ;
        RECT 23.600 29.700 27.600 30.300 ;
        RECT 23.600 29.600 24.400 29.700 ;
        RECT 26.800 29.600 27.600 29.700 ;
        RECT 41.200 30.300 42.000 30.400 ;
        RECT 47.600 30.300 48.400 30.400 ;
        RECT 41.200 29.700 48.400 30.300 ;
        RECT 41.200 29.600 42.000 29.700 ;
        RECT 47.600 29.600 48.400 29.700 ;
        RECT 55.600 30.300 56.400 30.400 ;
        RECT 95.600 30.300 96.400 30.400 ;
        RECT 55.600 29.700 96.400 30.300 ;
        RECT 55.600 29.600 56.400 29.700 ;
        RECT 95.600 29.600 96.400 29.700 ;
        RECT 98.800 30.300 99.600 30.400 ;
        RECT 102.000 30.300 102.800 30.400 ;
        RECT 106.800 30.300 107.600 30.400 ;
        RECT 116.400 30.300 117.200 30.400 ;
        RECT 124.400 30.300 125.200 30.400 ;
        RECT 98.800 29.700 125.200 30.300 ;
        RECT 98.800 29.600 99.600 29.700 ;
        RECT 102.000 29.600 102.800 29.700 ;
        RECT 106.800 29.600 107.600 29.700 ;
        RECT 116.400 29.600 117.200 29.700 ;
        RECT 124.400 29.600 125.200 29.700 ;
        RECT 146.800 30.300 147.600 30.400 ;
        RECT 151.600 30.300 152.400 30.400 ;
        RECT 146.800 29.700 152.400 30.300 ;
        RECT 146.800 29.600 147.600 29.700 ;
        RECT 151.600 29.600 152.400 29.700 ;
        RECT 26.800 28.300 27.600 28.400 ;
        RECT 42.800 28.300 43.600 28.400 ;
        RECT 26.800 27.700 43.600 28.300 ;
        RECT 26.800 27.600 27.600 27.700 ;
        RECT 42.800 27.600 43.600 27.700 ;
        RECT 76.400 28.300 77.200 28.400 ;
        RECT 102.000 28.300 102.800 28.400 ;
        RECT 76.400 27.700 102.800 28.300 ;
        RECT 76.400 27.600 77.200 27.700 ;
        RECT 102.000 27.600 102.800 27.700 ;
        RECT 148.400 28.300 149.200 28.400 ;
        RECT 180.400 28.300 181.200 28.400 ;
        RECT 194.800 28.300 195.600 28.400 ;
        RECT 148.400 27.700 195.600 28.300 ;
        RECT 148.400 27.600 149.200 27.700 ;
        RECT 180.400 27.600 181.200 27.700 ;
        RECT 194.800 27.600 195.600 27.700 ;
        RECT 210.800 28.300 211.600 28.400 ;
        RECT 220.400 28.300 221.200 28.400 ;
        RECT 210.800 27.700 221.200 28.300 ;
        RECT 210.800 27.600 211.600 27.700 ;
        RECT 220.400 27.600 221.200 27.700 ;
        RECT 7.600 26.300 8.400 26.400 ;
        RECT 47.600 26.300 48.400 26.400 ;
        RECT 7.600 25.700 48.400 26.300 ;
        RECT 7.600 25.600 8.400 25.700 ;
        RECT 47.600 25.600 48.400 25.700 ;
        RECT 62.000 26.300 62.800 26.400 ;
        RECT 79.600 26.300 80.400 26.400 ;
        RECT 62.000 25.700 80.400 26.300 ;
        RECT 62.000 25.600 62.800 25.700 ;
        RECT 79.600 25.600 80.400 25.700 ;
        RECT 140.400 26.300 141.200 26.400 ;
        RECT 164.400 26.300 165.200 26.400 ;
        RECT 172.400 26.300 173.200 26.400 ;
        RECT 223.600 26.300 224.400 26.400 ;
        RECT 140.400 25.700 224.400 26.300 ;
        RECT 140.400 25.600 141.200 25.700 ;
        RECT 164.400 25.600 165.200 25.700 ;
        RECT 172.400 25.600 173.200 25.700 ;
        RECT 223.600 25.600 224.400 25.700 ;
        RECT 100.400 24.300 101.200 24.400 ;
        RECT 143.600 24.300 144.400 24.400 ;
        RECT 100.400 23.700 144.400 24.300 ;
        RECT 100.400 23.600 101.200 23.700 ;
        RECT 143.600 23.600 144.400 23.700 ;
        RECT 74.800 20.300 75.600 20.400 ;
        RECT 79.600 20.300 80.400 20.400 ;
        RECT 74.800 19.700 80.400 20.300 ;
        RECT 74.800 19.600 75.600 19.700 ;
        RECT 79.600 19.600 80.400 19.700 ;
        RECT 223.600 20.300 224.400 20.400 ;
        RECT 228.400 20.300 229.200 20.400 ;
        RECT 223.600 19.700 229.200 20.300 ;
        RECT 223.600 19.600 224.400 19.700 ;
        RECT 228.400 19.600 229.200 19.700 ;
        RECT 94.000 18.300 94.800 18.400 ;
        RECT 100.400 18.300 101.200 18.400 ;
        RECT 94.000 17.700 101.200 18.300 ;
        RECT 94.000 17.600 94.800 17.700 ;
        RECT 100.400 17.600 101.200 17.700 ;
        RECT 26.800 16.300 27.600 16.400 ;
        RECT 47.600 16.300 48.400 16.400 ;
        RECT 26.800 15.700 48.400 16.300 ;
        RECT 26.800 15.600 27.600 15.700 ;
        RECT 47.600 15.600 48.400 15.700 ;
        RECT 121.200 16.300 122.000 16.400 ;
        RECT 142.000 16.300 142.800 16.400 ;
        RECT 121.200 15.700 142.800 16.300 ;
        RECT 121.200 15.600 122.000 15.700 ;
        RECT 142.000 15.600 142.800 15.700 ;
        RECT 188.400 16.300 189.200 16.400 ;
        RECT 201.200 16.300 202.000 16.400 ;
        RECT 188.400 15.700 202.000 16.300 ;
        RECT 188.400 15.600 189.200 15.700 ;
        RECT 201.200 15.600 202.000 15.700 ;
        RECT 7.600 14.300 8.400 14.400 ;
        RECT 41.200 14.300 42.000 14.400 ;
        RECT 7.600 13.700 42.000 14.300 ;
        RECT 7.600 13.600 8.400 13.700 ;
        RECT 41.200 13.600 42.000 13.700 ;
        RECT 90.800 14.300 91.600 14.400 ;
        RECT 169.200 14.300 170.000 14.400 ;
        RECT 190.000 14.300 190.800 14.400 ;
        RECT 90.800 13.700 190.800 14.300 ;
        RECT 90.800 13.600 91.600 13.700 ;
        RECT 169.200 13.600 170.000 13.700 ;
        RECT 190.000 13.600 190.800 13.700 ;
        RECT 198.000 14.300 198.800 14.400 ;
        RECT 225.200 14.300 226.000 14.400 ;
        RECT 198.000 13.700 226.000 14.300 ;
        RECT 198.000 13.600 198.800 13.700 ;
        RECT 225.200 13.600 226.000 13.700 ;
        RECT 44.400 12.300 45.200 12.400 ;
        RECT 52.400 12.300 53.200 12.400 ;
        RECT 44.400 11.700 53.200 12.300 ;
        RECT 44.400 11.600 45.200 11.700 ;
        RECT 52.400 11.600 53.200 11.700 ;
        RECT 111.600 12.300 112.400 12.400 ;
        RECT 122.800 12.300 123.600 12.400 ;
        RECT 111.600 11.700 123.600 12.300 ;
        RECT 111.600 11.600 112.400 11.700 ;
        RECT 122.800 11.600 123.600 11.700 ;
        RECT 151.600 12.300 152.400 12.400 ;
        RECT 159.600 12.300 160.400 12.400 ;
        RECT 151.600 11.700 160.400 12.300 ;
        RECT 151.600 11.600 152.400 11.700 ;
        RECT 159.600 11.600 160.400 11.700 ;
        RECT 201.200 12.300 202.000 12.400 ;
        RECT 204.400 12.300 205.200 12.400 ;
        RECT 201.200 11.700 205.200 12.300 ;
        RECT 201.200 11.600 202.000 11.700 ;
        RECT 204.400 11.600 205.200 11.700 ;
        RECT 215.600 11.600 216.400 12.400 ;
        RECT 244.400 12.300 245.200 12.400 ;
        RECT 249.200 12.300 250.000 12.400 ;
        RECT 244.400 11.700 250.000 12.300 ;
        RECT 244.400 11.600 245.200 11.700 ;
        RECT 249.200 11.600 250.000 11.700 ;
        RECT 119.600 10.300 120.400 10.400 ;
        RECT 124.400 10.300 125.200 10.400 ;
        RECT 119.600 9.700 125.200 10.300 ;
        RECT 119.600 9.600 120.400 9.700 ;
        RECT 124.400 9.600 125.200 9.700 ;
        RECT 207.600 10.300 208.400 10.400 ;
        RECT 244.400 10.300 245.200 10.400 ;
        RECT 207.600 9.700 245.200 10.300 ;
        RECT 207.600 9.600 208.400 9.700 ;
        RECT 244.400 9.600 245.200 9.700 ;
      LAYER metal4 ;
        RECT 42.600 95.400 43.800 110.600 ;
        RECT 77.800 97.400 79.000 134.600 ;
        RECT 87.400 53.400 88.600 150.600 ;
        RECT 132.200 117.400 133.400 140.600 ;
        RECT 148.200 107.400 149.400 170.600 ;
        RECT 177.000 137.400 178.200 144.600 ;
        RECT 100.200 51.400 101.400 102.600 ;
        RECT 177.000 99.400 178.200 134.600 ;
        RECT 196.200 49.400 197.400 76.600 ;
        RECT 218.600 71.400 219.800 176.600 ;
        RECT 234.600 129.400 235.800 168.600 ;
        RECT 237.800 135.400 239.000 156.600 ;
        RECT 215.400 11.400 216.600 32.600 ;
        RECT 244.200 11.400 245.400 70.600 ;
  END
END map9v3
END LIBRARY

